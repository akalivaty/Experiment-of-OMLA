//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1227;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n464), .A2(new_n466), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n466), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n465), .A2(KEYINPUT66), .A3(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT66), .B1(new_n465), .B2(G136), .ZN(new_n480));
  OAI221_X1 g055(.A(new_n476), .B1(new_n477), .B2(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT67), .ZN(G162));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n466), .A2(G114), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n489), .B(new_n491), .C1(new_n463), .C2(new_n462), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n466), .A2(G138), .ZN(new_n493));
  OR2_X1    g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n487), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(KEYINPUT69), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT69), .B1(new_n503), .B2(G543), .ZN(new_n504));
  OR2_X1    g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n505), .A2(G88), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n505), .A2(G62), .A3(new_n509), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND4_X1  g095(.A1(new_n505), .A2(G89), .A3(new_n508), .A4(new_n509), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT73), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n509), .B1(new_n504), .B2(new_n502), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  OR3_X1    g102(.A1(new_n526), .A2(KEYINPUT71), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT71), .B1(new_n526), .B2(new_n527), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n506), .A2(new_n507), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(KEYINPUT72), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n525), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT72), .B1(new_n530), .B2(new_n534), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(G168));
  NOR2_X1   g113(.A1(new_n526), .A2(new_n531), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G90), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT74), .B(G52), .Z(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n512), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n505), .A2(G64), .A3(new_n509), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(G171));
  XNOR2_X1  g122(.A(KEYINPUT75), .B(G43), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n539), .A2(G81), .B1(new_n533), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n526), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n505), .A2(G91), .A3(new_n508), .A4(new_n509), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n526), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(new_n537), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n572), .A2(new_n525), .A3(new_n535), .ZN(G286));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n526), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n505), .A2(G87), .A3(new_n508), .A4(new_n509), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n533), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n576), .A2(KEYINPUT76), .A3(new_n577), .A4(new_n578), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G288));
  AOI22_X1  g159(.A1(new_n539), .A2(G86), .B1(G48), .B2(new_n533), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n526), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n539), .A2(G85), .B1(G47), .B2(new_n533), .ZN(new_n591));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n526), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(new_n539), .A2(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n526), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n512), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n533), .A2(KEYINPUT77), .ZN(new_n608));
  AOI22_X1  g183(.A1(G651), .A2(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G171), .ZN(G284));
  OAI21_X1  g188(.A(new_n612), .B1(new_n611), .B2(G171), .ZN(G321));
  NAND2_X1  g189(.A1(G299), .A2(new_n611), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G168), .B2(new_n611), .ZN(G280));
  XOR2_X1   g191(.A(G280), .B(KEYINPUT78), .Z(G297));
  AND2_X1   g192(.A1(new_n601), .A2(new_n609), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT79), .B(G559), .Z(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(G860), .B2(new_n619), .ZN(G148));
  NAND3_X1  g195(.A1(new_n601), .A2(new_n609), .A3(new_n619), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n601), .A2(new_n609), .A3(KEYINPUT80), .A4(new_n619), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  MUX2_X1   g200(.A(new_n554), .B(new_n625), .S(G868), .Z(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n494), .A2(new_n495), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n467), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2100), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n465), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n475), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n466), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT81), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n640), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n646), .A2(KEYINPUT83), .A3(KEYINPUT14), .ZN(new_n647));
  AOI21_X1  g222(.A(KEYINPUT83), .B1(new_n646), .B2(KEYINPUT14), .ZN(new_n648));
  OAI22_X1  g223(.A1(new_n647), .A2(new_n648), .B1(new_n644), .B2(new_n645), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT17), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n664), .B2(new_n662), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT84), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n664), .A3(new_n662), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n664), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n673), .B1(new_n663), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n688), .B(new_n687), .S(new_n680), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT85), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT86), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n692), .A2(new_n696), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT87), .B(G1986), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n700), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n697), .B2(new_n698), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(G229));
  MUX2_X1   g279(.A(G24), .B(G290), .S(G16), .Z(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(G1986), .Z(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G25), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n465), .A2(G131), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n475), .A2(G119), .ZN(new_n710));
  OR2_X1    g285(.A1(G95), .A2(G2105), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n711), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n708), .B1(new_n714), .B2(new_n707), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G22), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G6), .B(G305), .S(G16), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT32), .B(G1981), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G23), .B(new_n579), .S(G16), .Z(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT33), .B(G1976), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n722), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n706), .B(new_n717), .C1(new_n729), .C2(KEYINPUT34), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT88), .Z(new_n731));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n729), .B2(KEYINPUT34), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(KEYINPUT36), .A3(new_n733), .ZN(new_n737));
  NOR2_X1   g312(.A1(G29), .A2(G35), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G162), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT29), .Z(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT94), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n618), .A2(new_n718), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G4), .B2(new_n718), .ZN(new_n745));
  INV_X1    g320(.A(G1348), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n748), .A2(G28), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n707), .B1(new_n748), .B2(G28), .ZN(new_n750));
  AND2_X1   g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  NOR2_X1   g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n749), .A2(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n707), .A2(G33), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n628), .A2(new_n466), .ZN(new_n757));
  INV_X1    g332(.A(G139), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n628), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(new_n466), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n754), .B1(new_n763), .B2(new_n707), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n753), .B1(new_n764), .B2(G2072), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n707), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  OAI211_X1 g342(.A(G140), .B(new_n466), .C1(new_n462), .C2(new_n463), .ZN(new_n768));
  OAI211_X1 g343(.A(G128), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n769));
  INV_X1    g344(.A(G116), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G104), .C2(G2105), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n768), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n707), .ZN(new_n774));
  INV_X1    g349(.A(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n765), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  NAND2_X1  g353(.A1(G160), .A2(G29), .ZN(new_n779));
  INV_X1    g354(.A(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n780), .B2(KEYINPUT24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(KEYINPUT24), .B2(new_n780), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n764), .A2(G2072), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n778), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n639), .B2(new_n707), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n747), .A2(new_n777), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n740), .A2(new_n741), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n718), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT95), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT23), .ZN(new_n791));
  INV_X1    g366(.A(G299), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n718), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT96), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n707), .A2(G32), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n475), .A2(G129), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT26), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n467), .A2(G105), .ZN(new_n802));
  INV_X1    g377(.A(G141), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n757), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n797), .B1(new_n807), .B2(new_n707), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT27), .B(G1996), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n746), .B2(new_n745), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n787), .A2(new_n788), .A3(new_n796), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n718), .A2(G21), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G168), .B2(new_n718), .ZN(new_n814));
  INV_X1    g389(.A(G1966), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n718), .A2(G19), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT90), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n555), .B2(new_n718), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT91), .ZN(new_n820));
  INV_X1    g395(.A(G1341), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n707), .A2(G27), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G164), .B2(new_n707), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT93), .ZN(new_n825));
  INV_X1    g400(.A(G2078), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n718), .A2(G5), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G171), .B2(new_n718), .ZN(new_n829));
  INV_X1    g404(.A(G1961), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n822), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n816), .B(new_n832), .C1(new_n821), .C2(new_n820), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n743), .A2(new_n812), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n736), .A2(new_n737), .A3(new_n834), .ZN(G150));
  INV_X1    g410(.A(G150), .ZN(G311));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(G67), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n526), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G651), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n539), .A2(G93), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n533), .A2(G55), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT98), .B(G860), .Z(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT97), .B1(new_n841), .B2(new_n844), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n840), .A2(new_n842), .A3(new_n850), .A4(new_n843), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n554), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n845), .A2(new_n555), .A3(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT38), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n618), .A2(G559), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n855), .B(new_n856), .Z(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n846), .B1(new_n858), .B2(KEYINPUT39), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n848), .B1(new_n859), .B2(new_n861), .ZN(G145));
  NAND2_X1  g437(.A1(new_n465), .A2(G142), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n475), .A2(G130), .ZN(new_n864));
  OR2_X1    g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n805), .B(KEYINPUT92), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n492), .B(KEYINPUT99), .C1(new_n496), .C2(new_n497), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n489), .B1(new_n462), .B2(new_n463), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT4), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT68), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n491), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT99), .B1(new_n876), .B2(new_n492), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n487), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n773), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n498), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n870), .ZN(new_n882));
  INV_X1    g457(.A(new_n773), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n487), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n879), .A2(KEYINPUT100), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n879), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n869), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n883), .B1(new_n882), .B2(new_n487), .ZN(new_n889));
  AOI211_X1 g464(.A(new_n486), .B(new_n773), .C1(new_n881), .C2(new_n870), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n879), .A2(KEYINPUT100), .A3(new_n884), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n807), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n762), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n805), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n889), .B2(new_n890), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n879), .A2(new_n805), .A3(new_n884), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n762), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n868), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n630), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n891), .A2(new_n807), .A3(new_n892), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n807), .B1(new_n891), .B2(new_n892), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n763), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n867), .A3(new_n898), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n901), .B1(new_n900), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n713), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n638), .B(G160), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(G162), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n894), .A2(new_n868), .A3(new_n899), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n867), .B1(new_n904), .B2(new_n898), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n630), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n900), .A2(new_n905), .A3(new_n901), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n714), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n908), .A2(new_n910), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT101), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n908), .A2(new_n915), .A3(new_n918), .A4(new_n910), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n910), .B1(new_n908), .B2(new_n915), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(G37), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n920), .A2(KEYINPUT40), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT40), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(G395));
  OAI21_X1  g500(.A(KEYINPUT106), .B1(new_n845), .B2(G868), .ZN(new_n926));
  XNOR2_X1  g501(.A(G290), .B(new_n579), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT104), .ZN(new_n928));
  XNOR2_X1  g503(.A(G303), .B(G305), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n927), .B2(KEYINPUT104), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n931), .A2(new_n932), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n930), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(G299), .A2(KEYINPUT103), .ZN(new_n939));
  INV_X1    g514(.A(new_n569), .ZN(new_n940));
  OR3_X1    g515(.A1(new_n940), .A2(KEYINPUT103), .A3(new_n564), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n618), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n610), .A2(KEYINPUT103), .A3(G299), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n623), .A2(KEYINPUT102), .A3(new_n624), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT102), .B1(new_n623), .B2(new_n624), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n854), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n854), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n625), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n952), .B2(new_n946), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n945), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n942), .A2(KEYINPUT41), .A3(new_n943), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT41), .B1(new_n942), .B2(new_n943), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n854), .B1(new_n947), .B2(new_n948), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n952), .A2(new_n950), .A3(new_n946), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n938), .B1(new_n961), .B2(KEYINPUT105), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n954), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n611), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n938), .A2(new_n963), .A3(new_n954), .A4(new_n960), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n926), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n944), .B1(new_n958), .B2(new_n959), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT105), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n938), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n964), .ZN(new_n973));
  AND4_X1   g548(.A1(new_n968), .A2(new_n973), .A3(G868), .A4(new_n966), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(new_n967), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(G868), .A3(new_n966), .ZN(new_n976));
  INV_X1    g551(.A(new_n926), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n978), .B(new_n979), .C1(KEYINPUT106), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(G295));
  NOR2_X1   g556(.A1(new_n967), .A2(new_n974), .ZN(G331));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  NAND3_X1  g558(.A1(G168), .A2(new_n983), .A3(G171), .ZN(new_n984));
  NAND2_X1  g559(.A1(G301), .A2(KEYINPUT108), .ZN(new_n985));
  NAND2_X1  g560(.A1(G171), .A2(new_n983), .ZN(new_n986));
  NAND3_X1  g561(.A1(G286), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n854), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n984), .A2(new_n950), .A3(new_n987), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n957), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n945), .A3(new_n990), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n994), .B2(new_n933), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n992), .A2(new_n935), .A3(new_n930), .A4(new_n993), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n1000));
  OR3_X1    g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n998), .B2(new_n999), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n878), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n468), .A2(G40), .A3(new_n472), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n878), .A2(KEYINPUT109), .A3(new_n1004), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n883), .B(new_n775), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n895), .A2(G1996), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1013), .B(new_n1014), .C1(new_n869), .C2(G1996), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT110), .Z(new_n1017));
  XOR2_X1   g592(.A(new_n713), .B(new_n716), .Z(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1011), .A2(G1986), .A3(G290), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT48), .Z(new_n1021));
  AND2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1011), .A2(G1996), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT46), .Z(new_n1024));
  AND2_X1   g599(.A1(new_n1013), .A2(new_n805), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1024), .B1(new_n1011), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1027));
  XOR2_X1   g602(.A(new_n1026), .B(new_n1027), .Z(new_n1028));
  NAND2_X1  g603(.A1(new_n714), .A2(new_n716), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1017), .A2(new_n1029), .B1(G2067), .B2(new_n883), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1022), .B(new_n1028), .C1(new_n1012), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT126), .ZN(new_n1032));
  XNOR2_X1  g607(.A(G290), .B(G1986), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1012), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1019), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n878), .A2(new_n1009), .A3(new_n1004), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1036), .B(G8), .C1(new_n579), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n581), .A2(new_n582), .A3(new_n1037), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(KEYINPUT115), .A3(new_n1040), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1040), .B1(new_n1038), .B2(KEYINPUT114), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(KEYINPUT114), .B2(new_n1038), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G305), .A2(G1981), .ZN(new_n1048));
  INV_X1    g623(.A(G1981), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n585), .A2(new_n1049), .A3(new_n589), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1036), .A2(G8), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1045), .A2(new_n1047), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n468), .A2(G40), .A3(new_n472), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n499), .A2(new_n1004), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(KEYINPUT50), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n487), .B2(new_n498), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT50), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT111), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1059), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n878), .A2(new_n1064), .A3(new_n1004), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n778), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT45), .B1(new_n878), .B2(new_n1004), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1009), .B1(new_n1060), .B2(new_n1008), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n815), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1058), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(G303), .B2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(KEYINPUT55), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n543), .B1(new_n515), .B2(new_n516), .ZN(new_n1078));
  OAI211_X1 g653(.A(G8), .B(new_n1077), .C1(new_n513), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1066), .A2(new_n741), .A3(new_n1067), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n878), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1060), .A2(new_n1008), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1009), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n721), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1072), .A2(new_n1087), .A3(G168), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT63), .B1(new_n1057), .B2(new_n1088), .ZN(new_n1089));
  AOI211_X1 g664(.A(G1976), .B(G288), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1050), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1054), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G8), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1094), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1064), .B1(new_n878), .B2(new_n1004), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1009), .B1(new_n1060), .B2(KEYINPUT50), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1098), .A2(new_n741), .B1(new_n1085), .B2(new_n721), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1081), .B1(new_n1099), .B2(new_n1058), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1081), .A2(new_n1058), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1101), .A2(KEYINPUT113), .A3(new_n1102), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1095), .A2(new_n1100), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1089), .B(new_n1092), .C1(new_n1107), .C2(new_n1057), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n830), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G2078), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1069), .A2(new_n1070), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1110), .A2(KEYINPUT123), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1961), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1114), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1083), .A2(new_n1084), .A3(new_n826), .A4(new_n1009), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(G301), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  AND4_X1   g699(.A1(new_n1047), .A2(new_n1100), .A3(new_n1045), .A4(new_n1056), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1093), .A2(G286), .ZN(new_n1128));
  NAND3_X1  g703(.A1(G168), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(G8), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1094), .A2(KEYINPUT122), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(KEYINPUT51), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(G8), .A3(new_n1129), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1127), .B1(KEYINPUT62), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1132), .A2(new_n1138), .A3(new_n1135), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1108), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1110), .A2(KEYINPUT125), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1083), .A2(new_n1009), .A3(new_n1112), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1143), .A2(new_n1144), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1118), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1141), .B1(new_n1148), .B2(G171), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1120), .A2(G301), .A3(new_n1123), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1100), .A2(new_n1045), .A3(new_n1047), .A4(new_n1056), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1136), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1096), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1059), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1956), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(KEYINPUT56), .B(G2072), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1083), .A2(new_n1084), .A3(new_n1009), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT117), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n795), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(new_n1163), .A3(new_n1159), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT57), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1165), .A2(KEYINPUT116), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(KEYINPUT116), .ZN(new_n1167));
  NAND3_X1  g742(.A1(G299), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n565), .A2(KEYINPUT116), .A3(new_n1165), .A4(new_n569), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1161), .A2(new_n1164), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(G1348), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1036), .A2(G2067), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1171), .B1(new_n610), .B2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1157), .A2(new_n1160), .A3(new_n1170), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(G1341), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1036), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT119), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1036), .A2(KEYINPUT119), .A3(new_n1180), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1183), .B(new_n1184), .C1(G1996), .C2(new_n1085), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT120), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1185), .A2(new_n555), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1187), .B1(new_n1185), .B2(new_n555), .ZN(new_n1189));
  OAI22_X1  g764(.A1(new_n1188), .A2(new_n1189), .B1(KEYINPUT120), .B2(new_n1186), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n610), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1174), .A2(KEYINPUT60), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT60), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1193), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1192), .A2(new_n618), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1190), .A2(new_n1191), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1162), .A2(new_n1159), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1197), .B1(new_n1176), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1171), .A2(new_n1177), .A3(KEYINPUT61), .ZN(new_n1202));
  OAI211_X1 g777(.A(KEYINPUT121), .B(new_n1197), .C1(new_n1176), .C2(new_n1198), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1178), .B1(new_n1196), .B2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1148), .A2(G171), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1141), .B1(new_n1124), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1154), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  AOI211_X1 g783(.A(new_n1032), .B(new_n1035), .C1(new_n1140), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1136), .A2(KEYINPUT62), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1210), .A2(new_n1124), .A3(new_n1153), .A4(new_n1139), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1108), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1190), .A2(new_n1191), .A3(new_n1195), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1204), .ZN(new_n1214));
  AOI22_X1  g789(.A1(new_n1213), .A2(new_n1214), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1207), .A2(new_n1136), .A3(new_n1153), .A4(new_n1151), .ZN(new_n1216));
  OAI211_X1 g791(.A(new_n1211), .B(new_n1212), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1035), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT126), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1031), .B1(new_n1209), .B2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g795(.A1(G227), .A2(new_n460), .ZN(new_n1222));
  OAI21_X1  g796(.A(new_n1222), .B1(new_n658), .B2(new_n659), .ZN(new_n1223));
  AOI21_X1  g797(.A(new_n1223), .B1(new_n701), .B2(new_n703), .ZN(new_n1224));
  OAI21_X1  g798(.A(new_n1224), .B1(new_n998), .B2(new_n999), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n1225), .B1(new_n920), .B2(new_n922), .ZN(G308));
  NAND2_X1  g800(.A1(new_n920), .A2(new_n922), .ZN(new_n1227));
  OAI211_X1 g801(.A(new_n1227), .B(new_n1224), .C1(new_n999), .C2(new_n998), .ZN(G225));
endmodule


