//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n559,
    new_n561, new_n562, new_n563, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n622, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT67), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT70), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(new_n462), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n471), .A2(G137), .A3(new_n472), .A4(new_n461), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT71), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND3_X1  g052(.A1(new_n471), .A2(G2105), .A3(new_n461), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT72), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n471), .A2(KEYINPUT72), .A3(G2105), .A4(new_n461), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n471), .A2(new_n472), .A3(new_n461), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n460), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n485), .A2(G136), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n471), .A2(G138), .A3(new_n472), .A4(new_n461), .ZN(new_n492));
  INV_X1    g067(.A(new_n464), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n494), .A2(new_n495), .A3(new_n472), .A4(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n494), .B2(new_n495), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n471), .A2(G126), .A3(G2105), .A4(new_n461), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n498), .A2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(G543), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT75), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n511), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n512));
  AND4_X1   g087(.A1(new_n504), .A2(new_n508), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  XOR2_X1   g088(.A(KEYINPUT76), .B(G88), .Z(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n504), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n508), .A2(G62), .A3(new_n510), .A4(new_n512), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n519), .B1(new_n522), .B2(G651), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  AOI211_X1 g099(.A(KEYINPUT77), .B(new_n524), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n515), .B(new_n518), .C1(new_n523), .C2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  AND3_X1   g102(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT78), .B(G51), .Z(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(new_n529), .B1(new_n517), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n513), .A2(G89), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT79), .B(KEYINPUT7), .Z(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  XNOR2_X1  g112(.A(KEYINPUT81), .B(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n513), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n517), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n508), .A2(G64), .A3(new_n510), .A4(new_n512), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n541), .B1(new_n544), .B2(G651), .ZN(new_n545));
  AOI211_X1 g120(.A(KEYINPUT80), .B(new_n524), .C1(new_n542), .C2(new_n543), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n539), .B(new_n540), .C1(new_n545), .C2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n517), .A2(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n513), .A2(G81), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT82), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n517), .A2(G53), .ZN(new_n565));
  AND2_X1   g140(.A1(KEYINPUT83), .A2(KEYINPUT9), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n550), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n513), .A2(G91), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(G299));
  OAI21_X1  g148(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n513), .A2(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n517), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND4_X1  g152(.A1(new_n508), .A2(G61), .A3(new_n510), .A4(new_n512), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n517), .A2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n513), .A2(G86), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n528), .A2(G60), .ZN(new_n585));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n524), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n517), .A2(G47), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n508), .A2(new_n504), .A3(new_n510), .A4(new_n512), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G301), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT84), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n513), .B2(G92), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n589), .A2(KEYINPUT84), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n550), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n513), .A2(new_n597), .A3(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT84), .B1(new_n589), .B2(new_n599), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n601), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n601), .A2(KEYINPUT85), .A3(new_n605), .A4(new_n608), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n595), .B1(new_n614), .B2(new_n594), .ZN(G284));
  AOI21_X1  g190(.A(new_n595), .B1(new_n614), .B2(new_n594), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G868), .ZN(G297));
  XOR2_X1   g194(.A(G297), .B(KEYINPUT86), .Z(G280));
  NOR2_X1   g195(.A1(new_n613), .A2(G559), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G860), .B2(new_n614), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT87), .ZN(G148));
  NAND2_X1  g198(.A1(new_n556), .A2(new_n594), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n621), .B2(new_n594), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n482), .A2(G123), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n485), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n462), .A2(new_n460), .A3(G2105), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n633), .B(new_n634), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2100), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n632), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT89), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G14), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT90), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n657), .B2(new_n660), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT92), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n671), .A2(new_n672), .ZN(new_n678));
  AOI22_X1  g253(.A1(new_n676), .A2(new_n677), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n673), .A2(new_n678), .A3(new_n675), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n680), .C1(new_n677), .C2(new_n676), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT94), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G21), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G168), .B2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(G1966), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G35), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT29), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n694), .B1(new_n698), .B2(G2090), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n480), .A2(G129), .A3(new_n481), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n485), .A2(G141), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT26), .Z(new_n704));
  NAND4_X1  g279(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G29), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G29), .B2(G32), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G11), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT31), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT28), .ZN(new_n713));
  INV_X1    g288(.A(G26), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G29), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(G29), .ZN(new_n716));
  OR2_X1    g291(.A1(G104), .A2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G116), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n460), .B1(new_n718), .B2(G2105), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n485), .A2(G140), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n480), .A2(G128), .A3(new_n481), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(G29), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(new_n713), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(G2067), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(G2067), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n710), .A2(new_n712), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n695), .A2(G27), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n695), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT104), .B(G2078), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n711), .A2(KEYINPUT31), .ZN(new_n732));
  NOR4_X1   g307(.A1(new_n699), .A2(new_n727), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n698), .A2(G2090), .ZN(new_n734));
  OR2_X1    g309(.A1(G29), .A2(G33), .ZN(new_n735));
  NAND2_X1  g310(.A1(G115), .A2(G2104), .ZN(new_n736));
  INV_X1    g311(.A(G127), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n464), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2105), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT100), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT25), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G139), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n484), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT99), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n741), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n735), .B1(new_n750), .B2(new_n695), .ZN(new_n751));
  INV_X1    g326(.A(G2072), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT103), .Z(new_n754));
  XOR2_X1   g329(.A(KEYINPUT101), .B(G34), .Z(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT24), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT24), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n756), .A2(new_n695), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT102), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n760), .B(new_n761), .C1(new_n476), .C2(new_n695), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n751), .A2(new_n752), .B1(new_n695), .B2(new_n765), .ZN(new_n766));
  AND4_X1   g341(.A1(new_n734), .A2(new_n754), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n690), .A2(G5), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G171), .B2(new_n690), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n708), .A2(new_n709), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n690), .A2(KEYINPUT23), .A3(G20), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT23), .ZN(new_n774));
  INV_X1    g349(.A(G20), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G16), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n776), .C1(new_n618), .C2(new_n690), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n772), .B(new_n778), .C1(new_n763), .C2(new_n762), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n733), .A2(new_n767), .A3(new_n771), .A4(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n690), .A2(G4), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n614), .B2(new_n690), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT97), .B(G1348), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n690), .A2(G6), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G305), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n789), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(G303), .A2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n690), .A2(G22), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n574), .A2(new_n575), .A3(G16), .A4(new_n576), .ZN(new_n798));
  NOR2_X1   g373(.A1(G16), .A2(G23), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT33), .B(G1976), .Z(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n793), .A2(new_n797), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n787), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n793), .A2(new_n804), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n797), .A2(new_n805), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n811), .A2(KEYINPUT96), .A3(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n690), .A2(G24), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n592), .B2(new_n690), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G1986), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n809), .A2(new_n810), .A3(new_n807), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(G1986), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n695), .A2(G25), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n482), .A2(G119), .ZN(new_n821));
  OR2_X1    g396(.A1(G95), .A2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(G107), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n460), .B1(new_n823), .B2(G2105), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n485), .A2(G131), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n820), .B1(new_n827), .B2(new_n695), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G1991), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  AND4_X1   g406(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n831), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n813), .A2(new_n814), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n814), .B1(new_n813), .B2(new_n832), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n781), .B(new_n786), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n631), .A2(new_n695), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n557), .A2(G16), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G16), .B2(G19), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT98), .B(G1341), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n835), .A2(new_n836), .A3(new_n841), .ZN(G311));
  INV_X1    g417(.A(new_n834), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n813), .A2(new_n832), .A3(new_n814), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n780), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n836), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n845), .A2(new_n846), .A3(new_n840), .A4(new_n786), .ZN(G150));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n589), .A2(new_n848), .B1(new_n849), .B2(new_n516), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI221_X1 g427(.A(KEYINPUT105), .B1(new_n516), .B2(new_n849), .C1(new_n589), .C2(new_n848), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(G80), .A2(G543), .ZN(new_n855));
  INV_X1    g430(.A(G67), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n550), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G651), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT106), .B(G860), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n557), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n854), .A2(new_n556), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n614), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n862), .B1(new_n869), .B2(new_n860), .ZN(G145));
  INV_X1    g445(.A(G142), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n484), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT109), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n482), .A2(G130), .ZN(new_n875));
  OR2_X1    g450(.A1(G106), .A2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n827), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n826), .A2(new_n875), .A3(new_n877), .A4(new_n874), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n635), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n635), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n497), .A2(new_n493), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n499), .A2(KEYINPUT107), .A3(new_n501), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT107), .B1(new_n499), .B2(new_n501), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n706), .A2(new_n722), .ZN(new_n892));
  INV_X1    g467(.A(new_n722), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n705), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n741), .A2(new_n748), .A3(new_n749), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT108), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n750), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n706), .A2(new_n722), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n893), .A2(new_n705), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n890), .A3(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n895), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n895), .A2(new_n903), .B1(KEYINPUT108), .B2(new_n896), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n881), .B(new_n884), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n884), .A2(new_n881), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n895), .A2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n897), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n895), .A2(new_n900), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n490), .B(new_n476), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n631), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n906), .A2(new_n911), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT110), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n906), .A2(new_n911), .A3(new_n919), .A4(new_n916), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g497(.A1(new_n621), .A2(new_n865), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n609), .A2(G299), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n618), .A2(new_n605), .A3(new_n608), .A4(new_n601), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n924), .A2(KEYINPUT41), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT41), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n865), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n613), .B2(G559), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n923), .A2(new_n930), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n924), .A2(new_n925), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g510(.A1(G166), .A2(G288), .ZN(new_n936));
  INV_X1    g511(.A(G288), .ZN(new_n937));
  NAND2_X1  g512(.A1(G303), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(G290), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G290), .B1(new_n936), .B2(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(G305), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  INV_X1    g518(.A(G305), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(new_n931), .C1(new_n932), .C2(new_n933), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n935), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n935), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n859), .A2(new_n594), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(G295));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n952), .ZN(G331));
  AND2_X1   g529(.A1(G301), .A2(G168), .ZN(new_n955));
  NOR2_X1   g530(.A1(G301), .A2(G168), .ZN(new_n956));
  INV_X1    g531(.A(new_n864), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n556), .B1(new_n854), .B2(new_n858), .ZN(new_n958));
  OAI22_X1  g533(.A1(new_n955), .A2(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n545), .A2(new_n546), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(G286), .A3(new_n539), .A4(new_n540), .ZN(new_n962));
  NAND2_X1  g537(.A1(G301), .A2(G168), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n962), .A2(new_n863), .A3(new_n963), .A4(new_n864), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n959), .A2(new_n960), .A3(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n865), .B(KEYINPUT111), .C1(new_n955), .C2(new_n956), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n928), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n968), .A3(new_n964), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n929), .A2(KEYINPUT112), .A3(new_n963), .A4(new_n962), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n933), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G37), .B1(new_n972), .B2(new_n946), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n942), .A2(new_n945), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(new_n971), .B2(new_n967), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT43), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n928), .A2(new_n969), .A3(new_n970), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n933), .B1(new_n965), .B2(new_n966), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n928), .A2(new_n965), .A3(new_n966), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n969), .A2(new_n970), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n946), .B(new_n980), .C1(new_n981), .C2(new_n933), .ZN(new_n982));
  INV_X1    g557(.A(G37), .ZN(new_n983));
  AND4_X1   g558(.A1(KEYINPUT43), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n976), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n973), .B2(new_n975), .ZN(new_n988));
  AND4_X1   g563(.A1(new_n987), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n985), .A2(new_n990), .ZN(G397));
  NAND4_X1  g566(.A1(new_n467), .A2(G40), .A3(new_n473), .A4(new_n475), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n890), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT45), .B(new_n993), .C1(new_n498), .C2(new_n502), .ZN(new_n997));
  AOI21_X1  g572(.A(G1966), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n498), .B2(new_n502), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n992), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n890), .A2(new_n1001), .A3(new_n993), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1002), .A3(new_n763), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(G8), .B(G168), .C1(new_n998), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT118), .ZN(new_n1006));
  INV_X1    g581(.A(new_n992), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n502), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n499), .A2(KEYINPUT107), .A3(new_n501), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1011), .B2(new_n887), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1007), .B(new_n997), .C1(new_n1012), .C2(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n693), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n1003), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(G8), .A4(G168), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1006), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n581), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n580), .A2(G651), .B1(new_n513), .B2(G86), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(G1981), .A4(new_n582), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n524), .B1(new_n578), .B2(new_n579), .ZN(new_n1023));
  OAI21_X1  g598(.A(G1981), .B1(new_n1023), .B2(KEYINPUT114), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G305), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(KEYINPUT115), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT49), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n994), .A2(new_n992), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1022), .A2(new_n1025), .A3(KEYINPUT115), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1027), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT116), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1027), .A2(new_n1035), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1030), .B1(new_n1038), .B2(G288), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n937), .B2(G1976), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1030), .B(new_n1042), .C1(new_n1038), .C2(G288), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n1045));
  AND3_X1   g620(.A1(G303), .A2(new_n1045), .A3(G8), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(G303), .B2(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n992), .B1(new_n999), .B2(new_n995), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n890), .A2(KEYINPUT45), .A3(new_n993), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n795), .ZN(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1000), .A2(new_n1002), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1029), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1018), .A2(new_n1037), .A3(new_n1044), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT63), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1034), .A2(new_n1036), .B1(new_n1043), .B2(new_n1041), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1001), .B(new_n993), .C1(new_n498), .C2(new_n502), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(new_n1007), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(new_n1053), .C1(new_n1001), .C2(new_n1012), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1029), .B1(new_n1052), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(new_n1048), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1017), .B2(new_n1006), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT113), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT55), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n1070));
  NAND3_X1  g645(.A1(G303), .A2(new_n1045), .A3(G8), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1067), .A2(new_n1072), .A3(new_n1055), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1059), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(G288), .A2(G1976), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT117), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1077));
  NOR2_X1   g652(.A1(G305), .A2(G1981), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1030), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1058), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1029), .B1(new_n1014), .B2(new_n1003), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G286), .A2(G8), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT121), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1081), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(new_n1083), .B(KEYINPUT121), .Z(new_n1086));
  NAND2_X1  g661(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1088), .A2(new_n763), .B1(new_n1013), .B2(new_n693), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT122), .B(new_n1086), .C1(new_n1089), .C2(new_n1029), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(new_n1090), .A3(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1015), .A2(new_n1084), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT51), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1081), .B(new_n1093), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT62), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1051), .B2(G2078), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1087), .A2(new_n770), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G2078), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n996), .A2(KEYINPUT53), .A3(new_n1101), .A4(new_n997), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(G171), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT123), .B(G171), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1048), .A2(new_n1064), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1073), .A2(new_n1109), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1110), .A2(new_n1059), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1091), .A2(new_n1112), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1096), .A2(new_n1108), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1087), .A2(new_n785), .ZN(new_n1116));
  INV_X1    g691(.A(G2067), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1028), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n613), .B(new_n1115), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n784), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n994), .A2(G2067), .A3(new_n992), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1120), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n613), .B2(new_n1115), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT120), .B1(new_n611), .B2(new_n612), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1121), .B(new_n1122), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  INV_X1    g704(.A(G1956), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1012), .A2(new_n1001), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1061), .A2(new_n1007), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n1134));
  XNOR2_X1  g709(.A(G299), .B(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1049), .A2(new_n1050), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1129), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1135), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT61), .A3(new_n1138), .ZN(new_n1145));
  INV_X1    g720(.A(G1996), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1049), .A2(new_n1050), .A3(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n994), .B2(new_n992), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n556), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT59), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1150), .B(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1128), .A2(new_n1141), .A3(new_n1145), .A4(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1138), .A2(new_n1119), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1140), .B1(new_n1155), .B2(new_n614), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  AND4_X1   g732(.A1(KEYINPUT53), .A2(new_n996), .A3(new_n1101), .A4(new_n1050), .ZN(new_n1158));
  OAI21_X1  g733(.A(G171), .B1(new_n1100), .B2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1102), .A2(new_n1098), .A3(G301), .A4(new_n1099), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(KEYINPUT54), .A3(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1110), .A2(new_n1059), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1100), .A2(new_n1158), .A3(G171), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1108), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1157), .A2(new_n1162), .A3(new_n1165), .A4(new_n1095), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1080), .A2(new_n1114), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n706), .A2(new_n1146), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n893), .A2(new_n1117), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n722), .A2(G2067), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n705), .A2(G1996), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n829), .B2(new_n826), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n827), .A2(new_n830), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OR2_X1    g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  NAND2_X1  g751(.A1(G290), .A2(G1986), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1012), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1167), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n994), .A2(new_n995), .A3(new_n1007), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1175), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1176), .A2(new_n1182), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT48), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1179), .A2(KEYINPUT46), .A3(new_n1146), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1169), .A2(new_n706), .A3(new_n1170), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1179), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT46), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(new_n1182), .B2(G1996), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1187), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT125), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n1193), .B(KEYINPUT47), .Z(new_n1194));
  XOR2_X1   g769(.A(new_n1174), .B(KEYINPUT124), .Z(new_n1195));
  OAI21_X1  g770(.A(new_n1169), .B1(new_n1195), .B2(new_n1172), .ZN(new_n1196));
  AOI211_X1 g771(.A(new_n1186), .B(new_n1194), .C1(new_n1179), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1181), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g773(.A(G319), .ZN(new_n1200));
  OR2_X1    g774(.A1(G227), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1201), .A2(KEYINPUT126), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n652), .A2(new_n1202), .ZN(new_n1203));
  OR2_X1    g777(.A1(new_n1201), .A2(KEYINPUT126), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n921), .A2(new_n688), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n982), .A2(new_n983), .ZN(new_n1206));
  INV_X1    g780(.A(new_n975), .ZN(new_n1207));
  OAI21_X1  g781(.A(KEYINPUT43), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n973), .A2(new_n987), .A3(new_n979), .ZN(new_n1209));
  AOI211_X1 g783(.A(new_n1203), .B(new_n1205), .C1(new_n1208), .C2(new_n1209), .ZN(G308));
  AOI21_X1  g784(.A(new_n1205), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1211));
  INV_X1    g785(.A(new_n1203), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1211), .A2(new_n1212), .ZN(G225));
endmodule


