//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT65), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT24), .ZN(new_n212));
  OR2_X1    g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT24), .A3(new_n211), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n216), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n210), .A2(new_n212), .A3(new_n214), .A4(new_n221), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n221), .A2(new_n212), .A3(new_n214), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G169gat), .ZN(new_n226));
  AOI21_X1  g025(.A(G176gat), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT25), .B1(new_n227), .B2(KEYINPUT23), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n222), .A2(KEYINPUT25), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT27), .B(G183gat), .ZN(new_n232));
  INV_X1    g031(.A(G190gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n231), .B(new_n233), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n230), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT26), .B1(new_n206), .B2(new_n208), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n215), .B1(new_n205), .B2(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT66), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(KEYINPUT28), .A3(new_n237), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n239), .A2(new_n243), .A3(new_n211), .A4(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n249), .B2(new_n248), .ZN(new_n251));
  XOR2_X1   g050(.A(G127gat), .B(G134gat), .Z(new_n252));
  INV_X1    g051(.A(G120gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G113gat), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT68), .B(G113gat), .Z(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(new_n253), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n251), .A2(new_n252), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n229), .A2(new_n247), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n229), .B2(new_n247), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n204), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G15gat), .B(G43gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(G71gat), .B(G99gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT33), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n261), .A2(KEYINPUT32), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n258), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n245), .A2(KEYINPUT28), .A3(new_n237), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT28), .B1(new_n245), .B2(new_n237), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n211), .B1(new_n240), .B2(new_n242), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n223), .A2(new_n228), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n221), .A2(new_n212), .A3(new_n214), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n217), .B1(new_n206), .B2(new_n208), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT25), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n270), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n229), .A2(new_n247), .A3(new_n258), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT32), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n282), .A2(new_n204), .B1(new_n283), .B2(KEYINPUT33), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n269), .B1(new_n284), .B2(new_n264), .ZN(new_n285));
  INV_X1    g084(.A(new_n204), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n286), .A3(new_n281), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT34), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT34), .A4(new_n286), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n290), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n293), .B(new_n269), .C1(new_n264), .C2(new_n284), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT70), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT36), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n292), .A2(new_n294), .A3(new_n300), .ZN(new_n301));
  OR3_X1    g100(.A1(new_n285), .A2(new_n291), .A3(new_n300), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n299), .B1(KEYINPUT36), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n274), .B2(new_n279), .ZN(new_n306));
  NAND2_X1  g105(.A1(G226gat), .A2(G233gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n274), .B2(new_n279), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT73), .ZN(new_n311));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT72), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n314));
  INV_X1    g113(.A(G197gat), .ZN(new_n315));
  INV_X1    g114(.A(G204gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G197gat), .A2(G204gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n313), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n229), .A2(new_n247), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n309), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n308), .A2(new_n311), .A3(new_n320), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n320), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n309), .B1(new_n321), .B2(new_n305), .ZN(new_n326));
  INV_X1    g125(.A(new_n310), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G36gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT74), .B(G8gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(KEYINPUT75), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n324), .A2(new_n328), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339));
  AND4_X1   g138(.A1(new_n339), .A2(new_n329), .A3(KEYINPUT30), .A4(new_n333), .ZN(new_n340));
  INV_X1    g139(.A(new_n333), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n324), .B2(new_n328), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n339), .B1(new_n342), .B2(KEYINPUT30), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n345));
  INV_X1    g144(.A(G148gat), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT77), .B1(new_n346), .B2(G141gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348));
  INV_X1    g147(.A(G141gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(G148gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(G141gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G155gat), .B(G162gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n355));
  AND2_X1   g154(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT79), .B(G162gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n345), .B1(new_n354), .B2(new_n360), .ZN(new_n361));
  OR2_X1    g160(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n362));
  INV_X1    g161(.A(G162gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G162gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n362), .A2(new_n364), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT2), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n369), .A2(KEYINPUT80), .A3(new_n353), .A4(new_n352), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n361), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n349), .A2(G148gat), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT2), .B1(new_n351), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(new_n353), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT82), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n361), .B2(new_n370), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n372), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n383), .B1(new_n371), .B2(new_n376), .ZN(new_n384));
  AOI211_X1 g183(.A(KEYINPUT81), .B(new_n375), .C1(new_n361), .C2(new_n370), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n386), .A3(new_n270), .ZN(new_n387));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n379), .A2(new_n258), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT4), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n387), .A2(KEYINPUT5), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT5), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n270), .B1(new_n384), .B2(new_n385), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n389), .ZN(new_n395));
  INV_X1    g194(.A(new_n388), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n391), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G85gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT0), .B(G57gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n402), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(new_n391), .C1(new_n392), .C2(new_n397), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n405), .A2(new_n407), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n344), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n379), .B(new_n383), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n372), .B1(new_n320), .B2(KEYINPUT29), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n378), .B2(new_n381), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n413), .B(new_n414), .C1(new_n415), .C2(new_n325), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n382), .A2(new_n305), .ZN(new_n417));
  INV_X1    g216(.A(new_n379), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n417), .A2(new_n320), .B1(new_n418), .B2(new_n412), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n416), .B1(new_n419), .B2(new_n414), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n423), .A2(G22gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n416), .B(new_n429), .C1(new_n419), .C2(new_n414), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n304), .B1(new_n410), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT76), .B1(new_n334), .B2(new_n337), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n342), .A2(new_n339), .A3(KEYINPUT30), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT85), .B1(new_n436), .B2(new_n338), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n338), .B(KEYINPUT85), .C1(new_n340), .C2(new_n343), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n387), .A2(KEYINPUT39), .A3(new_n390), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT39), .B1(new_n387), .B2(new_n390), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n396), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n395), .A2(KEYINPUT39), .A3(new_n388), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n402), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n443), .A2(new_n402), .A3(new_n446), .A4(new_n444), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n405), .A2(KEYINPUT87), .ZN(new_n450));
  INV_X1    g249(.A(new_n389), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n411), .B2(new_n270), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT5), .B1(new_n452), .B2(new_n388), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n404), .A4(new_n391), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n448), .A2(new_n449), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n433), .B1(new_n440), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n450), .A2(new_n457), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n404), .B1(new_n455), .B2(new_n391), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n406), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n464));
  NAND2_X1  g263(.A1(new_n329), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n465), .B(new_n341), .C1(new_n466), .C2(new_n329), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n342), .B1(new_n467), .B2(KEYINPUT38), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n308), .A2(new_n310), .A3(new_n320), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n308), .A2(new_n311), .A3(new_n323), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT37), .B(new_n469), .C1(new_n470), .C2(new_n320), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n471), .A2(new_n465), .A3(new_n472), .A4(new_n335), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n463), .A2(new_n409), .A3(new_n468), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n432), .B1(new_n459), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT35), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n302), .A2(new_n301), .B1(new_n428), .B2(new_n430), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n437), .B2(new_n439), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n405), .A2(new_n407), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n460), .B2(new_n462), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n298), .A2(new_n431), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n410), .A2(KEYINPUT35), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT89), .B1(new_n475), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n448), .A2(new_n449), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n344), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n486), .A2(new_n460), .A3(new_n488), .A4(new_n438), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n474), .A3(new_n431), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n295), .B2(new_n297), .ZN(new_n492));
  INV_X1    g291(.A(new_n303), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n491), .ZN(new_n494));
  INV_X1    g293(.A(new_n410), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n433), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n479), .B1(new_n462), .B2(new_n405), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n298), .A2(new_n431), .A3(KEYINPUT35), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n499), .A2(new_n500), .A3(new_n344), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n488), .A2(new_n438), .ZN(new_n502));
  AOI211_X1 g301(.A(new_n406), .B(new_n461), .C1(new_n450), .C2(new_n457), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n502), .B(new_n477), .C1(new_n503), .C2(new_n479), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n504), .B2(new_n476), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n497), .A2(new_n498), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n485), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(new_n315), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT11), .B(G169gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  XOR2_X1   g310(.A(new_n511), .B(KEYINPUT12), .Z(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(KEYINPUT16), .A3(new_n515), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(G8gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(G8gat), .ZN(new_n521));
  INV_X1    g320(.A(G8gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n516), .A2(new_n517), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n526), .A2(G29gat), .A3(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(G29gat), .ZN(new_n528));
  INV_X1    g327(.A(G36gat), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT14), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT91), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT92), .B(G36gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G29gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(G50gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G43gat), .ZN(new_n537));
  INV_X1    g336(.A(G43gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G50gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(KEYINPUT15), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT15), .B1(new_n539), .B2(KEYINPUT93), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n540), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n537), .B(new_n539), .C1(KEYINPUT93), .C2(KEYINPUT15), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n544), .A2(new_n531), .A3(new_n534), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(KEYINPUT17), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n542), .B2(new_n548), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n525), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT96), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n525), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n556), .A2(new_n557), .A3(new_n549), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n556), .B2(new_n549), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n553), .B(new_n554), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n554), .B(KEYINPUT13), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n558), .A2(new_n559), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n556), .A2(new_n549), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n556), .A2(new_n549), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT97), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n556), .A2(new_n557), .A3(new_n549), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n571), .A2(KEYINPUT18), .A3(new_n554), .A4(new_n553), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n562), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n513), .B1(new_n573), .B2(KEYINPUT90), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(KEYINPUT90), .A3(new_n513), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n507), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT98), .Z(new_n581));
  INV_X1    g380(.A(G57gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(G64gat), .ZN(new_n583));
  INV_X1    g382(.A(G64gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G57gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  INV_X1    g386(.A(G71gat), .ZN(new_n588));
  INV_X1    g387(.A(G78gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n585), .B(KEYINPUT100), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n583), .B(KEYINPUT99), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n590), .B(new_n580), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT101), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n598), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G211gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n596), .A2(new_n597), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n556), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G183gat), .ZN(new_n610));
  OR3_X1    g409(.A1(new_n556), .A2(G183gat), .A3(new_n608), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n611), .A3(new_n607), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n605), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n616), .A2(new_n612), .A3(new_n604), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n602), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n604), .B1(new_n616), .B2(new_n612), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n613), .A2(new_n614), .A3(new_n605), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n601), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT7), .ZN(new_n624));
  INV_X1    g423(.A(G99gat), .ZN(new_n625));
  INV_X1    g424(.A(G106gat), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT8), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n624), .B(new_n627), .C1(G85gat), .C2(G92gat), .ZN(new_n628));
  XOR2_X1   g427(.A(G99gat), .B(G106gat), .Z(new_n629));
  OR2_X1    g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n592), .A3(new_n631), .A4(new_n595), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT103), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n592), .A2(new_n595), .ZN(new_n635));
  INV_X1    g434(.A(new_n631), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n628), .A2(new_n629), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n635), .A2(new_n638), .A3(new_n639), .A4(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n630), .A2(new_n631), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n596), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT102), .B(KEYINPUT10), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n632), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G230gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n203), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT105), .B(G204gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT104), .B(G176gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n643), .A2(new_n632), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n650), .B(new_n656), .C1(new_n649), .C2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n648), .B1(new_n641), .B2(new_n645), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n649), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n642), .B1(new_n550), .B2(new_n552), .ZN(new_n663));
  NAND3_X1  g462(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n549), .A2(new_n638), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G190gat), .B(G218gat), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  XNOR2_X1  g468(.A(G134gat), .B(G162gat), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n666), .A2(new_n667), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n666), .A2(new_n667), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n662), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n622), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n579), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n499), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n515), .ZN(G1324gat));
  INV_X1    g482(.A(new_n680), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT16), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n522), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n522), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n684), .A2(new_n440), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G8gat), .B1(new_n680), .B2(new_n502), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(G1325gat));
  AND3_X1   g493(.A1(new_n684), .A2(G15gat), .A3(new_n494), .ZN(new_n695));
  AOI21_X1  g494(.A(G15gat), .B1(new_n684), .B2(new_n303), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(G1326gat));
  OR3_X1    g496(.A1(new_n680), .A2(G22gat), .A3(new_n431), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n699));
  OAI21_X1  g498(.A(G22gat), .B1(new_n680), .B2(new_n431), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(G1327gat));
  OAI21_X1  g502(.A(new_n673), .B1(new_n668), .B2(new_n669), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n675), .A2(new_n672), .A3(new_n676), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n577), .A2(new_n622), .A3(new_n662), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n507), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n528), .A3(new_n499), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT107), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n708), .A2(new_n712), .A3(new_n528), .A4(new_n499), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n711), .B1(new_n710), .B2(new_n713), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n485), .A2(new_n506), .ZN(new_n717));
  INV_X1    g516(.A(new_n706), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n475), .B2(new_n484), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n497), .A2(KEYINPUT108), .A3(new_n505), .ZN(new_n723));
  AOI211_X1 g522(.A(new_n706), .B(new_n720), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n707), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n725), .A2(new_n499), .A3(new_n726), .ZN(new_n727));
  OAI22_X1  g526(.A1(new_n714), .A2(new_n715), .B1(new_n528), .B2(new_n727), .ZN(G1328gat));
  INV_X1    g527(.A(new_n533), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n708), .A2(new_n729), .A3(new_n440), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT46), .Z(new_n731));
  AND3_X1   g530(.A1(new_n725), .A2(new_n440), .A3(new_n726), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n729), .B2(new_n732), .ZN(G1329gat));
  OAI211_X1 g532(.A(new_n494), .B(new_n726), .C1(new_n719), .C2(new_n724), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G43gat), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n708), .A2(new_n538), .A3(new_n303), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1330gat));
  OAI211_X1 g538(.A(new_n433), .B(new_n726), .C1(new_n719), .C2(new_n724), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n708), .A2(new_n536), .A3(new_n433), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1331gat));
  AOI21_X1  g544(.A(new_n622), .B1(new_n722), .B2(new_n723), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n577), .A2(new_n718), .A3(new_n662), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n681), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT110), .B(G57gat), .Z(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1332gat));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n746), .A2(KEYINPUT111), .A3(new_n747), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n502), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  AOI21_X1  g558(.A(new_n304), .B1(new_n753), .B2(new_n754), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n303), .A2(new_n588), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n760), .A2(new_n588), .B1(new_n748), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n762), .B(new_n764), .ZN(G1334gat));
  AOI21_X1  g564(.A(new_n431), .B1(new_n753), .B2(new_n754), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(new_n589), .ZN(G1335gat));
  AND2_X1   g566(.A1(new_n618), .A2(new_n621), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n577), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n662), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n725), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(G85gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n772), .A2(new_n773), .A3(new_n681), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n770), .B1(new_n497), .B2(new_n505), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n776), .A3(new_n718), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n769), .B(new_n718), .C1(new_n475), .C2(new_n484), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n662), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n499), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n774), .B1(new_n773), .B2(new_n783), .ZN(G1336gat));
  OAI211_X1 g583(.A(new_n440), .B(new_n771), .C1(new_n719), .C2(new_n724), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n502), .A2(G92gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n781), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n662), .B1(new_n778), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n775), .A2(KEYINPUT113), .A3(new_n776), .A4(new_n718), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n779), .A4(new_n788), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT114), .B1(new_n795), .B2(KEYINPUT52), .ZN(new_n796));
  INV_X1    g595(.A(new_n794), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n785), .B2(G92gat), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n798), .A2(new_n799), .A3(new_n787), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n790), .B1(new_n796), .B2(new_n800), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n772), .B2(new_n304), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n625), .A3(new_n303), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT115), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n780), .B2(new_n804), .ZN(G1338gat));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n433), .B(new_n771), .C1(new_n719), .C2(new_n724), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n431), .A2(G106gat), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n792), .A2(new_n793), .A3(new_n779), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n777), .A2(new_n779), .A3(new_n782), .A4(new_n810), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n807), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n808), .B2(G106gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n806), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n811), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n808), .B2(G106gat), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n818), .B(KEYINPUT116), .C1(new_n807), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n816), .A2(new_n821), .ZN(G1339gat));
  NAND3_X1  g621(.A1(new_n641), .A2(new_n648), .A3(new_n645), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n656), .B1(new_n659), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n658), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n705), .A3(new_n704), .ZN(new_n832));
  INV_X1    g631(.A(new_n511), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n565), .A2(new_n566), .A3(new_n564), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n554), .B1(new_n571), .B2(new_n553), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT117), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n573), .A2(new_n513), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n832), .A2(new_n678), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n831), .ZN(new_n843));
  INV_X1    g642(.A(new_n576), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n843), .B(new_n706), .C1(new_n844), .C2(new_n574), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n768), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n577), .A2(new_n622), .A3(new_n678), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n499), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n502), .A3(new_n477), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n578), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n502), .A3(new_n482), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n578), .A2(new_n255), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n850), .B2(new_n662), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n782), .A2(new_n253), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n852), .B2(new_n856), .ZN(G1341gat));
  INV_X1    g656(.A(G127gat), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n850), .A2(new_n858), .A3(new_n622), .ZN(new_n859));
  INV_X1    g658(.A(new_n852), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n768), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n859), .B1(new_n861), .B2(new_n858), .ZN(G1342gat));
  NOR3_X1   g661(.A1(new_n852), .A2(G134gat), .A3(new_n706), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n850), .B2(new_n706), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1343gat));
  OAI21_X1  g665(.A(new_n433), .B1(new_n846), .B2(new_n847), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n681), .A2(new_n440), .A3(new_n494), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n349), .A3(new_n577), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n869), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n867), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(KEYINPUT57), .B(new_n433), .C1(new_n846), .C2(new_n847), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n879), .A2(KEYINPUT118), .A3(new_n577), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT118), .B1(new_n879), .B2(new_n577), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n874), .B1(new_n882), .B2(G141gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n577), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G141gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n873), .B1(new_n885), .B2(new_n872), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT119), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n886), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n880), .A2(new_n881), .A3(new_n349), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n874), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n891), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n878), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n782), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n875), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n346), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT120), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(KEYINPUT59), .C1(new_n895), .C2(new_n346), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n871), .A2(new_n346), .A3(new_n782), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1345gat));
  AOI21_X1  g703(.A(new_n358), .B1(new_n871), .B2(new_n768), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n622), .A2(new_n357), .A3(new_n356), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n879), .B2(new_n906), .ZN(G1346gat));
  NAND2_X1  g706(.A1(new_n879), .A2(new_n718), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n359), .A3(new_n910), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n870), .A2(new_n359), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n706), .B2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n502), .A2(new_n499), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n848), .A2(new_n477), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n578), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n848), .A2(new_n482), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n224), .A2(new_n226), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n577), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n916), .B1(new_n918), .B2(new_n920), .ZN(G1348gat));
  INV_X1    g720(.A(new_n915), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(G176gat), .A3(new_n782), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT122), .ZN(new_n924));
  INV_X1    g723(.A(new_n918), .ZN(new_n925));
  AOI21_X1  g724(.A(G176gat), .B1(new_n925), .B2(new_n782), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n924), .A2(new_n926), .ZN(G1349gat));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n768), .A3(new_n232), .ZN(new_n928));
  OAI21_X1  g727(.A(G183gat), .B1(new_n915), .B2(new_n622), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n928), .A2(new_n929), .B1(KEYINPUT123), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT123), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(G1350gat));
  AOI21_X1  g732(.A(new_n233), .B1(new_n922), .B2(new_n718), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n233), .A3(new_n718), .ZN(new_n942));
  NAND2_X1  g741(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n939), .A2(new_n940), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n936), .A2(new_n937), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n914), .A2(new_n304), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n867), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT126), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n315), .A3(new_n577), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n877), .B2(new_n878), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n577), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n951), .B1(new_n953), .B2(new_n315), .ZN(G1352gat));
  NOR3_X1   g753(.A1(new_n867), .A2(G204gat), .A3(new_n947), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n955), .A2(new_n782), .B1(KEYINPUT127), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(KEYINPUT127), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(G204gat), .B1(new_n894), .B2(new_n947), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n957), .A2(new_n958), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G1353gat));
  NAND2_X1  g761(.A1(new_n952), .A2(new_n768), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n622), .A2(G211gat), .ZN(new_n966));
  OAI22_X1  g765(.A1(new_n964), .A2(new_n965), .B1(new_n949), .B2(new_n966), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n950), .B2(new_n718), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n718), .A2(G218gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n952), .B2(new_n969), .ZN(G1355gat));
endmodule


