//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n218), .B1(new_n202), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT64), .B(G77), .Z(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT65), .B(G244), .Z(new_n222));
  AOI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n217), .B1(new_n212), .B2(new_n211), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  OR2_X1    g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1698), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g0053(.A1(G222), .A2(new_n250), .B1(new_n221), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n248), .A2(new_n249), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G1698), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n260), .A2(new_n263), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G226), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT73), .B1(new_n270), .B2(G190), .ZN(new_n271));
  INV_X1    g0071(.A(G200), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n262), .A2(KEYINPUT73), .A3(G190), .A4(new_n268), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n208), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n213), .ZN(new_n276));
  INV_X1    g0076(.A(G13), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G50), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n206), .B2(G20), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n281), .A2(new_n283), .B1(new_n282), .B2(new_n280), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n207), .A2(new_n285), .A3(KEYINPUT68), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(G20), .B2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G150), .ZN(new_n290));
  OAI21_X1  g0090(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n207), .A2(G33), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n290), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n276), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n274), .B1(new_n297), .B2(KEYINPUT9), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n284), .A2(new_n295), .A3(KEYINPUT9), .ZN(new_n299));
  NOR4_X1   g0099(.A1(new_n271), .A2(new_n273), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n273), .A2(KEYINPUT72), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT72), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n270), .B2(new_n272), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n271), .A2(new_n298), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n300), .A2(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n309), .A2(KEYINPUT69), .A3(new_n293), .ZN(new_n310));
  INV_X1    g0110(.A(new_n292), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n289), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n221), .A2(G20), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT69), .B1(new_n309), .B2(new_n293), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n310), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n221), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n315), .A2(new_n276), .B1(new_n316), .B2(new_n280), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n208), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n279), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n206), .A2(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G77), .ZN(new_n321));
  OR3_X1    g0121(.A1(new_n319), .A2(KEYINPUT70), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT70), .B1(new_n319), .B2(new_n321), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n250), .A2(G232), .B1(new_n253), .B2(G107), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n219), .B2(new_n257), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n261), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n266), .B1(new_n267), .B2(new_n222), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n325), .B1(G200), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT71), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n328), .A2(new_n329), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n331), .A2(new_n332), .B1(G190), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n332), .B2(new_n331), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n269), .A2(G169), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(new_n269), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n296), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(G179), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n330), .A2(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n325), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n308), .A2(new_n335), .A3(new_n339), .A4(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT75), .A2(G169), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n346));
  INV_X1    g0146(.A(G1698), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n256), .A2(G226), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n261), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT13), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n266), .B1(new_n267), .B2(G238), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n351), .B2(new_n353), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n345), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT14), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n355), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n351), .A2(new_n353), .A3(KEYINPUT74), .A4(new_n352), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(G179), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n345), .C1(new_n354), .C2(new_n355), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n357), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT76), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n357), .A2(KEYINPUT76), .A3(new_n363), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n289), .A2(G50), .ZN(new_n371));
  INV_X1    g0171(.A(new_n293), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n318), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT11), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n278), .A2(G20), .A3(new_n202), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT12), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n320), .A2(G68), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n375), .B(new_n377), .C1(new_n319), .C2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n374), .A2(KEYINPUT11), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n370), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n360), .A2(new_n361), .A3(G190), .A4(new_n362), .ZN(new_n384));
  OAI21_X1  g0184(.A(G200), .B1(new_n354), .B2(new_n355), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n344), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n248), .A2(new_n207), .A3(new_n249), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT7), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n202), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n289), .A2(G159), .ZN(new_n394));
  XNOR2_X1  g0194(.A(G58), .B(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G20), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n393), .A2(new_n397), .A3(KEYINPUT16), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n253), .B2(new_n207), .ZN(new_n400));
  NOR4_X1   g0200(.A1(new_n251), .A2(new_n252), .A3(new_n390), .A4(G20), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n289), .A2(G159), .B1(new_n395), .B2(G20), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n276), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n292), .B1(new_n206), .B2(G20), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n281), .A2(new_n406), .B1(new_n280), .B2(new_n292), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT77), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT16), .B1(new_n393), .B2(new_n397), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n399), .A3(new_n403), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n318), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  INV_X1    g0212(.A(new_n407), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(G226), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n416));
  OAI211_X1 g0216(.A(G223), .B(new_n347), .C1(new_n251), .C2(new_n252), .ZN(new_n417));
  INV_X1    g0217(.A(G87), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n285), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n261), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n260), .A2(G232), .A3(new_n263), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT78), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT78), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n260), .A2(new_n263), .A3(new_n425), .A4(G232), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(new_n265), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G169), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n424), .A2(new_n426), .A3(new_n265), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G179), .A3(new_n422), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n429), .A2(KEYINPUT79), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT79), .B1(new_n429), .B2(new_n431), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT80), .B1(new_n415), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n405), .A2(KEYINPUT77), .A3(new_n407), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT80), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT79), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n428), .A2(new_n337), .ZN(new_n441));
  INV_X1    g0241(.A(G169), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n430), .B2(new_n422), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n429), .A2(KEYINPUT79), .A3(new_n431), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n438), .A2(new_n439), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT18), .B1(new_n435), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n439), .B1(new_n438), .B2(new_n446), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n434), .A2(KEYINPUT80), .A3(new_n437), .A4(new_n436), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  INV_X1    g0253(.A(G190), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n430), .A2(KEYINPUT81), .A3(new_n454), .A4(new_n422), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n428), .B2(new_n272), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n428), .A2(G190), .ZN(new_n458));
  OAI211_X1 g0258(.A(KEYINPUT82), .B(new_n455), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n411), .A2(new_n413), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n430), .A2(new_n454), .A3(new_n422), .ZN(new_n462));
  AOI21_X1  g0262(.A(G200), .B1(new_n430), .B2(new_n422), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n456), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT82), .B1(new_n464), .B2(new_n455), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n453), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT83), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT82), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(KEYINPUT17), .A3(new_n460), .A4(new_n459), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n467), .B1(new_n466), .B2(new_n471), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n448), .B(new_n452), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n388), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n256), .A2(new_n207), .A3(G68), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT19), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n207), .B1(new_n349), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n418), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(G107), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n478), .B1(new_n349), .B2(G20), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n477), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n276), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n280), .A2(new_n309), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n206), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n318), .A2(new_n279), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT84), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT84), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n318), .A2(new_n490), .A3(new_n279), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n485), .B(new_n486), .C1(new_n492), .C2(new_n309), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n256), .A2(G244), .A3(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G116), .ZN(new_n495));
  INV_X1    g0295(.A(new_n250), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n494), .B(new_n495), .C1(new_n496), .C2(new_n219), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n261), .ZN(new_n498));
  INV_X1    g0298(.A(G45), .ZN(new_n499));
  OAI21_X1  g0299(.A(G250), .B1(new_n499), .B2(G1), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n502), .A2(new_n260), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n337), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n503), .B1(new_n497), .B2(new_n261), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n442), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n493), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n489), .A2(G87), .A3(new_n491), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n510), .A2(new_n485), .A3(new_n486), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n505), .A2(G190), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n507), .A2(G200), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n289), .A2(G77), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  INV_X1    g0318(.A(G107), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n480), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n517), .B1(new_n524), .B2(new_n207), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n519), .B1(new_n391), .B2(new_n392), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n276), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n280), .A2(new_n480), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n528), .C1(new_n480), .C2(new_n492), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n347), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n256), .A2(G244), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n256), .A2(G250), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n347), .B1(new_n534), .B2(KEYINPUT4), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n261), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G41), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n206), .B(G45), .C1(new_n537), .C2(KEYINPUT5), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT85), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT86), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT5), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(G41), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(KEYINPUT86), .A3(KEYINPUT5), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n260), .A2(new_n543), .A3(G274), .A4(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n543), .A2(new_n544), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n260), .B1(new_n547), .B2(new_n538), .ZN(new_n548));
  INV_X1    g0348(.A(G257), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n536), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n442), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n538), .B(KEYINPUT85), .ZN(new_n554));
  INV_X1    g0354(.A(new_n545), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT87), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(new_n557), .C1(new_n549), .C2(new_n548), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT87), .B1(new_n546), .B2(new_n550), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(new_n536), .A4(new_n337), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n529), .A2(new_n553), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n558), .A3(new_n536), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT88), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT88), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n558), .A2(new_n559), .A3(new_n536), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n272), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n552), .A2(new_n454), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(new_n529), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n516), .B(new_n561), .C1(new_n566), .C2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n285), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(G20), .B1(new_n572), .B2(new_n531), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n207), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n571), .B1(new_n576), .B2(new_n318), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n276), .B(KEYINPUT20), .C1(new_n573), .C2(new_n575), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n488), .A2(G116), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G116), .B2(new_n280), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n253), .A2(G303), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n496), .C2(new_n549), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n261), .ZN(new_n585));
  INV_X1    g0385(.A(new_n548), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT89), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(G270), .ZN(new_n588));
  INV_X1    g0388(.A(G270), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT89), .B1(new_n548), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n585), .A2(new_n588), .A3(new_n556), .A4(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n591), .A2(new_n272), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(G190), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n579), .B(new_n581), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n581), .A2(new_n579), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n595), .A3(G169), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n591), .A2(new_n595), .A3(KEYINPUT21), .A4(G169), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n591), .A2(new_n337), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n595), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n594), .A2(new_n598), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n256), .A2(new_n207), .A3(G87), .ZN(new_n603));
  XNOR2_X1  g0403(.A(KEYINPUT90), .B(KEYINPUT22), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n604), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(new_n207), .A3(G87), .A4(new_n256), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT23), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(G20), .B2(new_n519), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n495), .A2(G20), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT24), .A4(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n276), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(new_n607), .A3(new_n612), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT24), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n489), .A2(G107), .A3(new_n491), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n278), .A2(G20), .A3(new_n519), .ZN(new_n620));
  XOR2_X1   g0420(.A(new_n620), .B(KEYINPUT25), .Z(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n256), .A2(G250), .A3(new_n347), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT91), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n256), .A2(KEYINPUT91), .A3(G250), .A4(new_n347), .ZN(new_n626));
  NAND2_X1  g0426(.A1(G33), .A2(G294), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n256), .A2(G257), .A3(G1698), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n261), .B1(G264), .B2(new_n586), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n630), .A2(G179), .A3(new_n556), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n442), .B1(new_n630), .B2(new_n556), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n622), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n619), .A2(new_n621), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n630), .A2(new_n454), .A3(new_n556), .ZN(new_n635));
  AOI21_X1  g0435(.A(G200), .B1(new_n630), .B2(new_n556), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n618), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NOR4_X1   g0438(.A1(new_n476), .A2(new_n570), .A3(new_n602), .A4(new_n638), .ZN(G372));
  AOI22_X1  g0439(.A1(new_n340), .A2(new_n341), .B1(new_n324), .B2(new_n317), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n386), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n383), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n466), .A2(new_n471), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT83), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n460), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n445), .A3(new_n444), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT18), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n434), .A2(new_n450), .A3(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n308), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(new_n339), .ZN(new_n654));
  INV_X1    g0454(.A(new_n509), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n515), .A2(new_n561), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n515), .B2(new_n561), .ZN(new_n659));
  INV_X1    g0459(.A(new_n633), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n598), .A2(new_n601), .A3(new_n599), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n637), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n658), .B(new_n659), .C1(new_n570), .C2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n654), .B1(new_n476), .B2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(G330), .ZN(new_n666));
  INV_X1    g0466(.A(new_n602), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT92), .ZN(new_n668));
  INV_X1    g0468(.A(new_n278), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .A3(G20), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT27), .B1(new_n669), .B2(G20), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n667), .A2(new_n668), .B1(new_n595), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n668), .B2(new_n667), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n661), .A2(new_n595), .A3(new_n674), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n666), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n633), .A2(new_n674), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n622), .A2(new_n674), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n637), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n660), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n674), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n661), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n680), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0492(.A(new_n210), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n481), .A2(G107), .A3(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n215), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  NAND2_X1  g0499(.A1(new_n663), .A2(new_n687), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT29), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n602), .A2(new_n638), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n561), .A2(new_n509), .A3(new_n514), .ZN(new_n703));
  INV_X1    g0503(.A(new_n566), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(new_n568), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n705), .A3(new_n687), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT94), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n630), .A2(new_n551), .A3(new_n536), .A4(new_n507), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n546), .B1(new_n261), .B2(new_n584), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(G179), .A3(new_n590), .A4(new_n588), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n707), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n707), .B(KEYINPUT30), .C1(new_n708), .C2(new_n710), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n630), .A2(new_n556), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n507), .A2(G179), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n562), .A3(new_n591), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  INV_X1    g0521(.A(new_n718), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n713), .B2(new_n714), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n721), .B1(new_n723), .B2(new_n687), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n706), .A2(new_n720), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n701), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n699), .B1(new_n729), .B2(new_n206), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT95), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n277), .A2(G20), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G45), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n695), .A2(G1), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n676), .A2(new_n666), .A3(new_n677), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n679), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n676), .A2(new_n677), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n207), .A2(G190), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n272), .A2(G179), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G283), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G329), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G303), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n207), .A2(new_n454), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n742), .ZN(new_n753));
  INV_X1    g0553(.A(G326), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n337), .A2(new_n272), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n750), .B1(new_n751), .B2(new_n753), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n337), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n741), .A2(new_n758), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G322), .A2(new_n760), .B1(new_n762), .B2(G311), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n755), .A2(new_n741), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT33), .B(G317), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n256), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G294), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n746), .A2(G190), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n763), .B(new_n767), .C1(new_n768), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n757), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT99), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n756), .A2(new_n282), .B1(new_n759), .B2(new_n201), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n221), .B2(new_n762), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  NOR2_X1   g0577(.A1(new_n743), .A2(new_n519), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n256), .B1(new_n753), .B2(new_n418), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n778), .B(new_n779), .C1(G68), .C2(new_n765), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n771), .A2(new_n480), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT98), .B(G159), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n747), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n777), .A2(new_n780), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n773), .A2(KEYINPUT99), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n774), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n213), .B1(G20), .B2(new_n442), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n734), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n693), .A2(new_n253), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G355), .B1(new_n574), .B2(new_n693), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n216), .A2(G45), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n243), .B2(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n693), .A2(new_n256), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n792), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(KEYINPUT96), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT96), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n739), .A2(new_n789), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n740), .B(new_n790), .C1(new_n798), .C2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n736), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  INV_X1    g0604(.A(new_n734), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT101), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n343), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n640), .A2(KEYINPUT101), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n325), .A2(new_n674), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n335), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n663), .A2(new_n687), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n812), .A2(KEYINPUT102), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n809), .A2(new_n335), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n640), .A2(new_n674), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n663), .B2(new_n687), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n813), .B(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n805), .B1(new_n819), .B2(new_n727), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n727), .B2(new_n819), .ZN(new_n821));
  INV_X1    g0621(.A(new_n789), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G143), .A2(new_n760), .B1(new_n765), .B2(G150), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n756), .C1(new_n761), .C2(new_n783), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n256), .B1(new_n747), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n753), .A2(new_n282), .B1(new_n743), .B2(new_n202), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(G58), .C2(new_n770), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n827), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n753), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n256), .B(new_n781), .C1(G107), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n764), .A2(new_n836), .B1(new_n761), .B2(new_n574), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT100), .Z(new_n838));
  NOR2_X1   g0638(.A1(new_n743), .A2(new_n418), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n759), .A2(new_n768), .B1(new_n747), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n756), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n839), .B(new_n841), .C1(G303), .C2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n835), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n822), .B1(new_n833), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G77), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n789), .A2(new_n737), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n734), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n816), .B2(new_n738), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n821), .A2(new_n849), .ZN(G384));
  INV_X1    g0650(.A(new_n524), .ZN(new_n851));
  OAI211_X1 g0651(.A(G116), .B(new_n214), .C1(new_n851), .C2(KEYINPUT35), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(KEYINPUT35), .B2(new_n851), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT36), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n216), .B(new_n221), .C1(new_n201), .C2(new_n202), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n282), .A2(G68), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n206), .B(G13), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n809), .A2(new_n674), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n812), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n381), .A2(new_n687), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n387), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n381), .B1(new_n368), .B2(new_n369), .ZN(new_n863));
  INV_X1    g0663(.A(new_n386), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n863), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  INV_X1    g0670(.A(new_n672), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n648), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n875), .B2(new_n646), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n434), .A2(new_n437), .A3(new_n436), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n436), .A2(new_n437), .A3(new_n871), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n470), .A2(new_n460), .A3(new_n459), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n649), .A3(new_n872), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n880), .A2(new_n881), .B1(KEYINPUT37), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n870), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n872), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n474), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n883), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n869), .A2(new_n889), .B1(new_n652), .B2(new_n672), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n881), .A2(new_n649), .A3(new_n879), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n880), .A2(new_n881), .B1(KEYINPUT37), .B2(new_n891), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n892), .A2(KEYINPUT104), .ZN(new_n893));
  INV_X1    g0693(.A(new_n879), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n650), .A2(new_n466), .A3(new_n471), .A4(new_n651), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n892), .A2(KEYINPUT104), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n870), .B(new_n883), .C1(new_n474), .C2(new_n885), .ZN(new_n898));
  XNOR2_X1  g0698(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n886), .B2(new_n887), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT39), .B1(new_n901), .B2(new_n898), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT103), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT103), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n889), .A2(new_n904), .A3(KEYINPUT39), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n900), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n863), .A2(new_n687), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n890), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT29), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n663), .B2(new_n687), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n339), .B(new_n653), .C1(new_n912), .C2(new_n476), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n908), .B(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT106), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n915), .A2(KEYINPUT31), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n719), .A2(new_n674), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n916), .B1(new_n723), .B2(new_n687), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n706), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n861), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n383), .B2(new_n386), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n920), .B(new_n816), .C1(new_n922), .C2(new_n865), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n889), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n924), .B(KEYINPUT40), .C1(new_n897), .C2(new_n898), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n388), .A2(new_n475), .A3(new_n920), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(G330), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n914), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n206), .B2(new_n732), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n914), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n858), .B1(new_n935), .B2(new_n936), .ZN(G367));
  NOR2_X1   g0737(.A1(new_n796), .A2(new_n239), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n800), .B1(new_n210), .B2(new_n309), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n805), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n834), .A2(KEYINPUT46), .A3(G116), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n941), .B(new_n253), .C1(new_n768), .C2(new_n764), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n744), .A2(G97), .ZN(new_n943));
  INV_X1    g0743(.A(G317), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n747), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n756), .A2(new_n840), .B1(new_n759), .B2(new_n751), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT46), .B1(new_n834), .B2(G116), .ZN(new_n947));
  NOR4_X1   g0747(.A1(new_n942), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n771), .A2(new_n519), .B1(new_n836), .B2(new_n761), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT107), .ZN(new_n950));
  XNOR2_X1  g0750(.A(KEYINPUT108), .B(G137), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n256), .B1(new_n747), .B2(new_n951), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n316), .A2(new_n743), .B1(new_n282), .B2(new_n761), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(G68), .C2(new_n770), .ZN(new_n954));
  INV_X1    g0754(.A(G150), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n955), .A2(new_n759), .B1(new_n764), .B2(new_n783), .ZN(new_n956));
  INV_X1    g0756(.A(G143), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n756), .A2(new_n957), .B1(new_n753), .B2(new_n201), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n948), .A2(new_n950), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n960), .A2(KEYINPUT47), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n822), .B1(new_n960), .B2(KEYINPUT47), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n940), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n511), .A2(new_n687), .ZN(new_n964));
  MUX2_X1   g0764(.A(new_n516), .B(new_n655), .S(new_n964), .Z(new_n965));
  INV_X1    g0765(.A(new_n739), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n733), .A2(G1), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n569), .A2(new_n566), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n529), .A2(new_n674), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n561), .A2(new_n970), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n969), .A2(new_n971), .B1(new_n561), .B2(new_n687), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n690), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT45), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n690), .A2(new_n972), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT44), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n686), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n976), .B(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n685), .B1(new_n980), .B2(new_n974), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n684), .B(new_n688), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n678), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n728), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n728), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n694), .B(KEYINPUT41), .Z(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n968), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n689), .A2(new_n972), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n561), .B1(new_n969), .B2(new_n633), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n687), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n991), .B2(KEYINPUT42), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n990), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n685), .A2(new_n972), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n967), .B1(new_n989), .B2(new_n1000), .ZN(G387));
  INV_X1    g0801(.A(new_n985), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1002), .A2(new_n695), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n728), .B2(new_n984), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n696), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n791), .A2(new_n1005), .B1(new_n519), .B2(new_n693), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n696), .B(new_n499), .C1(new_n202), .C2(new_n846), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT109), .Z(new_n1008));
  NAND2_X1  g0808(.A1(new_n311), .A2(new_n282), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT50), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n795), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n236), .A2(new_n499), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1006), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n734), .B1(new_n1013), .B2(new_n800), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n842), .A2(G159), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT110), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G50), .A2(new_n760), .B1(new_n765), .B2(new_n311), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(new_n256), .A3(new_n943), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G68), .A2(new_n762), .B1(new_n748), .B2(G150), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n316), .B2(new_n753), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n771), .A2(new_n309), .ZN(new_n1021));
  NOR4_X1   g0821(.A1(new_n1016), .A2(new_n1018), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n834), .A2(G294), .B1(new_n770), .B2(G283), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G317), .A2(new_n760), .B1(new_n762), .B2(G303), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(KEYINPUT111), .B(G322), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n840), .B2(new_n764), .C1(new_n756), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n253), .B1(new_n747), .B2(new_n754), .C1(new_n574), .C2(new_n743), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n1029), .B2(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1022), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1014), .B1(new_n1033), .B2(new_n822), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n684), .B2(new_n739), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n984), .B2(new_n968), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1004), .A2(new_n1036), .ZN(G393));
  INV_X1    g0837(.A(new_n982), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n968), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n771), .A2(new_n846), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n764), .A2(new_n282), .B1(new_n761), .B2(new_n292), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n253), .A4(new_n839), .ZN(new_n1042));
  INV_X1    g0842(.A(G159), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n756), .A2(new_n955), .B1(new_n759), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT51), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n753), .A2(new_n202), .B1(new_n747), .B2(new_n957), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT112), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1042), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n756), .A2(new_n944), .B1(new_n759), .B2(new_n840), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n753), .A2(new_n836), .B1(new_n761), .B2(new_n768), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n764), .A2(new_n751), .B1(new_n747), .B2(new_n1025), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n256), .B(new_n778), .C1(G116), .C2(new_n770), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1050), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n822), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n800), .B1(new_n480), .B2(new_n210), .C1(new_n796), .C2(new_n246), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n805), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n972), .B2(new_n966), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1038), .A2(new_n1002), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n694), .B1(new_n982), .B2(new_n985), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1039), .B(new_n1060), .C1(new_n1061), .C2(new_n1062), .ZN(G390));
  INV_X1    g0863(.A(KEYINPUT114), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n930), .A2(new_n666), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n913), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n811), .A2(new_n809), .B1(new_n640), .B2(new_n674), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n862), .B2(new_n866), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n860), .B1(new_n1068), .B2(new_n727), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n666), .B1(new_n814), .B2(new_n815), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n920), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n922), .A2(new_n865), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n1072), .A3(KEYINPUT115), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1069), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1072), .B1(new_n726), .B2(new_n1067), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n867), .A2(new_n920), .A3(new_n1070), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n860), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n701), .A2(new_n475), .A3(new_n388), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n931), .A2(G330), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(new_n654), .A4(KEYINPUT114), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1066), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n900), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n868), .A2(new_n907), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n904), .B1(new_n889), .B2(KEYINPUT39), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT39), .ZN(new_n1090));
  AOI211_X1 g0890(.A(KEYINPUT103), .B(new_n1090), .C1(new_n884), .C2(new_n888), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1087), .B(new_n1088), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n726), .A2(new_n1072), .A3(new_n1067), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n897), .A2(new_n898), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n907), .B(KEYINPUT113), .Z(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n868), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1092), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1095), .A2(new_n868), .A3(new_n1096), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n906), .B2(new_n1088), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1086), .B(new_n1098), .C1(new_n1100), .C2(new_n1079), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n694), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(KEYINPUT116), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT116), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1104), .A3(new_n694), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1086), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1098), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1079), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1103), .A2(new_n1105), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n968), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n734), .B1(new_n292), .B2(new_n847), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT117), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n256), .B1(new_n743), .B2(new_n282), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  INV_X1    g0916(.A(G125), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n756), .A2(new_n1116), .B1(new_n747), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1115), .B(new_n1118), .C1(G159), .C2(new_n770), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n753), .A2(new_n955), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT53), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n764), .A2(new_n951), .B1(new_n761), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G132), .B2(new_n760), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1119), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n256), .B(new_n1040), .C1(G87), .C2(new_n834), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G107), .A2(new_n765), .B1(new_n762), .B2(G97), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G283), .A2(new_n842), .B1(new_n760), .B2(G116), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n743), .A2(new_n202), .B1(new_n747), .B2(new_n768), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT118), .Z(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n822), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1114), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n906), .B2(new_n737), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1112), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1110), .A2(new_n1140), .ZN(G378));
  AOI21_X1  g0941(.A(new_n734), .B1(new_n282), .B2(new_n847), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(G33), .A2(G41), .ZN(new_n1143));
  INV_X1    g0943(.A(G124), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1143), .B1(new_n747), .B2(new_n1144), .C1(new_n743), .C2(new_n783), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n756), .A2(new_n1117), .B1(new_n764), .B2(new_n829), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n762), .A2(G137), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n1116), .B2(new_n759), .C1(new_n753), .C2(new_n1122), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(G150), .C2(new_n770), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1145), .B1(new_n1150), .B2(KEYINPUT59), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(KEYINPUT59), .B2(new_n1150), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G41), .B(new_n256), .C1(new_n834), .C2(new_n221), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n201), .B2(new_n743), .C1(new_n836), .C2(new_n747), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT120), .Z(new_n1155));
  OAI22_X1  g0955(.A1(new_n764), .A2(new_n480), .B1(new_n761), .B2(new_n309), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n756), .A2(new_n574), .B1(new_n759), .B2(new_n519), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(G68), .C2(new_n770), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(KEYINPUT58), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1152), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT58), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G50), .B(new_n1143), .C1(new_n253), .C2(new_n537), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n306), .A2(new_n307), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n271), .A2(new_n298), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n273), .A2(new_n299), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n301), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n339), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT121), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT121), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n308), .A2(new_n1171), .A3(new_n339), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n297), .A2(new_n672), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT55), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1170), .A2(new_n1175), .A3(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT123), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1177), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1142), .B1(new_n822), .B2(new_n1163), .C1(new_n1185), .C2(new_n738), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT124), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n923), .B1(new_n884), .B2(new_n888), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n928), .B(G330), .C1(KEYINPUT40), .C2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1185), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n927), .A2(new_n1185), .A3(G330), .A4(new_n928), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n908), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1087), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n907), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1197), .A2(new_n890), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1187), .B1(new_n1199), .B2(new_n968), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1066), .A2(new_n1085), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1101), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n694), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1199), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1200), .B1(new_n1207), .B2(new_n1208), .ZN(G375));
  INV_X1    g1009(.A(new_n1082), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1201), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1106), .A2(new_n988), .A3(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n867), .A2(new_n738), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT125), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n951), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G132), .A2(new_n842), .B1(new_n760), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n253), .B1(new_n744), .B2(G58), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n282), .C2(new_n771), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n747), .A2(new_n1116), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1043), .A2(new_n753), .B1(new_n764), .B2(new_n1122), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G150), .C2(new_n762), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n764), .A2(new_n574), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n480), .A2(new_n753), .B1(new_n759), .B2(new_n836), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G294), .C2(new_n842), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n846), .A2(new_n743), .B1(new_n761), .B2(new_n519), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n253), .B1(new_n747), .B2(new_n751), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1021), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1219), .A2(new_n1222), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(new_n822), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n734), .B(new_n1230), .C1(new_n202), .C2(new_n847), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1082), .A2(new_n968), .B1(new_n1214), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1212), .A2(new_n1232), .ZN(G381));
  OR2_X1    g1033(.A1(new_n1112), .A2(new_n1139), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n1103), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1101), .A2(new_n1202), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1206), .B(new_n694), .C1(KEYINPUT57), .C2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1200), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(G390), .ZN(new_n1240));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1004), .A2(new_n803), .A3(new_n1036), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1244));
  OR4_X1    g1044(.A1(G387), .A2(new_n1239), .A3(G381), .A4(new_n1244), .ZN(G407));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G343), .C2(new_n1239), .ZN(G409));
  NAND2_X1  g1046(.A1(G387), .A2(new_n1240), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT126), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n803), .B1(new_n1004), .B2(new_n1036), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1248), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G390), .B(new_n967), .C1(new_n989), .C2(new_n1000), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1247), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n989), .A2(new_n1000), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1254), .A2(new_n1250), .A3(new_n967), .A4(G390), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1243), .A2(new_n1249), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G387), .A2(new_n1240), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1253), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1203), .A2(new_n988), .A3(new_n1199), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1200), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1110), .A3(new_n1140), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(G375), .B2(new_n1236), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  INV_X1    g1064(.A(G213), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(G343), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1211), .A2(KEYINPUT60), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1211), .A2(KEYINPUT60), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n694), .B(new_n1106), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(G384), .A3(new_n1232), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(G384), .B1(new_n1271), .B2(new_n1232), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1263), .A2(new_n1264), .A3(new_n1267), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G378), .A2(new_n1200), .A3(new_n1238), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1266), .B1(new_n1278), .B2(new_n1262), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G2897), .B(new_n1266), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1274), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1266), .A2(G2897), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1272), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1276), .B(new_n1277), .C1(new_n1279), .C2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1264), .B1(new_n1279), .B2(new_n1275), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1259), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT63), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1279), .A2(new_n1275), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1258), .A2(new_n1277), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1263), .A2(new_n1267), .A3(new_n1275), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(KEYINPUT63), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1287), .A2(new_n1294), .ZN(G405));
  XNOR2_X1  g1095(.A(new_n1258), .B(new_n1275), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G375), .A2(G378), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1239), .A2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1296), .B(new_n1298), .ZN(G402));
endmodule


