

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723;

  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n433) );
  INV_X1 U376 ( .A(G953), .ZN(n711) );
  XNOR2_X2 U377 ( .A(n462), .B(n461), .ZN(n522) );
  NOR2_X1 U378 ( .A1(n651), .A2(n707), .ZN(n652) );
  NOR2_X1 U379 ( .A1(n663), .A2(n707), .ZN(n665) );
  NOR2_X1 U380 ( .A1(n657), .A2(n707), .ZN(n658) );
  OR2_X1 U381 ( .A1(n579), .A2(n472), .ZN(n509) );
  XNOR2_X1 U382 ( .A(G143), .B(G128), .ZN(n406) );
  BUF_X1 U383 ( .A(n644), .Z(n623) );
  XNOR2_X1 U384 ( .A(n514), .B(KEYINPUT39), .ZN(n568) );
  NOR2_X1 U385 ( .A1(n611), .A2(n478), .ZN(n479) );
  AND2_X1 U386 ( .A1(n650), .A2(G953), .ZN(n707) );
  NOR2_X1 U387 ( .A1(n623), .A2(n710), .ZN(n578) );
  AND2_X1 U388 ( .A1(n614), .A2(n354), .ZN(n615) );
  NOR2_X1 U389 ( .A1(n569), .A2(n572), .ZN(n535) );
  XOR2_X1 U390 ( .A(n451), .B(n450), .Z(n353) );
  XOR2_X1 U391 ( .A(n613), .B(KEYINPUT122), .Z(n354) );
  AND2_X1 U392 ( .A1(n547), .A2(n546), .ZN(n355) );
  NOR2_X1 U393 ( .A1(n666), .A2(n622), .ZN(n471) );
  AND2_X1 U394 ( .A1(n355), .A2(n562), .ZN(n563) );
  AND2_X1 U395 ( .A1(n564), .A2(n563), .ZN(n567) );
  XNOR2_X1 U396 ( .A(n406), .B(n366), .ZN(n367) );
  NOR2_X1 U397 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U398 ( .A(n368), .B(n367), .ZN(n371) );
  OR2_X1 U399 ( .A1(n474), .A2(n473), .ZN(n477) );
  OR2_X1 U400 ( .A1(n512), .A2(n517), .ZN(n380) );
  XNOR2_X1 U401 ( .A(n503), .B(KEYINPUT45), .ZN(n644) );
  OR2_X1 U402 ( .A1(n696), .A2(G902), .ZN(n432) );
  XNOR2_X1 U403 ( .A(n477), .B(n476), .ZN(n611) );
  XNOR2_X1 U404 ( .A(n460), .B(KEYINPUT25), .ZN(n461) );
  BUF_X1 U405 ( .A(n642), .Z(n710) );
  AND2_X1 U406 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U407 ( .A(n466), .B(n465), .ZN(n666) );
  XNOR2_X1 U408 ( .A(n619), .B(n618), .ZN(G75) );
  XNOR2_X1 U409 ( .A(G116), .B(G113), .ZN(n357) );
  XNOR2_X1 U410 ( .A(KEYINPUT3), .B(G119), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n438) );
  XNOR2_X1 U412 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n358), .B(G122), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n438), .B(n359), .ZN(n363) );
  XNOR2_X1 U415 ( .A(G107), .B(G104), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n360), .B(G110), .ZN(n362) );
  XNOR2_X1 U417 ( .A(G101), .B(KEYINPUT73), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n429) );
  XNOR2_X1 U419 ( .A(n363), .B(n429), .ZN(n629) );
  XOR2_X1 U420 ( .A(KEYINPUT18), .B(KEYINPUT90), .Z(n365) );
  XNOR2_X1 U421 ( .A(KEYINPUT75), .B(KEYINPUT17), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n368) );
  NAND2_X1 U423 ( .A1(n711), .A2(G224), .ZN(n366) );
  INV_X1 U424 ( .A(G146), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n369), .B(G125), .ZN(n390) );
  XNOR2_X1 U426 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n423) );
  XNOR2_X1 U427 ( .A(n390), .B(n423), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n629), .B(n372), .ZN(n654) );
  XNOR2_X1 U430 ( .A(G902), .B(KEYINPUT15), .ZN(n637) );
  NAND2_X1 U431 ( .A1(n654), .A2(n637), .ZN(n377) );
  INV_X1 U432 ( .A(G902), .ZN(n443) );
  INV_X1 U433 ( .A(G237), .ZN(n373) );
  NAND2_X1 U434 ( .A1(n443), .A2(n373), .ZN(n378) );
  NAND2_X1 U435 ( .A1(n378), .A2(G210), .ZN(n375) );
  INV_X1 U436 ( .A(KEYINPUT77), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n512) );
  NAND2_X1 U439 ( .A1(n378), .A2(G214), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n379), .B(KEYINPUT91), .ZN(n517) );
  XNOR2_X1 U441 ( .A(n380), .B(KEYINPUT19), .ZN(n539) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n381), .B(KEYINPUT14), .ZN(n384) );
  AND2_X1 U444 ( .A1(G953), .A2(n384), .ZN(n382) );
  NAND2_X1 U445 ( .A1(G902), .A2(n382), .ZN(n505) );
  NOR2_X1 U446 ( .A1(G898), .A2(n505), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n383), .B(KEYINPUT92), .ZN(n385) );
  NAND2_X1 U448 ( .A1(G952), .A2(n384), .ZN(n609) );
  NOR2_X1 U449 ( .A1(G953), .A2(n609), .ZN(n508) );
  NOR2_X1 U450 ( .A1(n385), .A2(n508), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n386), .B(KEYINPUT93), .ZN(n387) );
  NAND2_X1 U452 ( .A1(n539), .A2(n387), .ZN(n389) );
  XNOR2_X1 U453 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n388) );
  XNOR2_X2 U454 ( .A(n389), .B(n388), .ZN(n490) );
  XNOR2_X1 U455 ( .A(n390), .B(KEYINPUT10), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n391), .B(KEYINPUT67), .ZN(n709) );
  XNOR2_X1 U457 ( .A(G113), .B(G143), .ZN(n392) );
  INV_X1 U458 ( .A(G140), .ZN(n620) );
  XNOR2_X1 U459 ( .A(n620), .B(G131), .ZN(n426) );
  XNOR2_X1 U460 ( .A(n392), .B(n426), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n709), .B(n393), .ZN(n401) );
  XOR2_X1 U462 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n395) );
  NAND2_X1 U463 ( .A1(G214), .A2(n433), .ZN(n394) );
  XNOR2_X1 U464 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U465 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n397) );
  XNOR2_X1 U466 ( .A(G104), .B(G122), .ZN(n396) );
  XNOR2_X1 U467 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n647) );
  NAND2_X1 U470 ( .A1(n647), .A2(n443), .ZN(n405) );
  XOR2_X1 U471 ( .A(KEYINPUT13), .B(KEYINPUT99), .Z(n403) );
  XNOR2_X1 U472 ( .A(KEYINPUT100), .B(G475), .ZN(n402) );
  XOR2_X1 U473 ( .A(n403), .B(n402), .Z(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n493) );
  INV_X1 U475 ( .A(n493), .ZN(n555) );
  XNOR2_X1 U476 ( .A(n406), .B(G134), .ZN(n425) );
  XOR2_X1 U477 ( .A(KEYINPUT9), .B(G122), .Z(n408) );
  XNOR2_X1 U478 ( .A(G116), .B(G107), .ZN(n407) );
  XNOR2_X1 U479 ( .A(n408), .B(n407), .ZN(n413) );
  XOR2_X1 U480 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n411) );
  NAND2_X1 U481 ( .A1(G234), .A2(n711), .ZN(n409) );
  XOR2_X1 U482 ( .A(KEYINPUT8), .B(n409), .Z(n455) );
  NAND2_X1 U483 ( .A1(G217), .A2(n455), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U485 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U486 ( .A(n425), .B(n414), .ZN(n702) );
  NAND2_X1 U487 ( .A1(n702), .A2(n443), .ZN(n417) );
  INV_X1 U488 ( .A(KEYINPUT102), .ZN(n415) );
  XNOR2_X1 U489 ( .A(n415), .B(G478), .ZN(n416) );
  XNOR2_X1 U490 ( .A(n417), .B(n416), .ZN(n548) );
  NAND2_X1 U491 ( .A1(n555), .A2(n548), .ZN(n598) );
  NAND2_X1 U492 ( .A1(n637), .A2(G234), .ZN(n418) );
  XNOR2_X1 U493 ( .A(n418), .B(KEYINPUT20), .ZN(n459) );
  AND2_X1 U494 ( .A1(n459), .A2(G221), .ZN(n420) );
  INV_X1 U495 ( .A(KEYINPUT21), .ZN(n419) );
  XNOR2_X1 U496 ( .A(n420), .B(n419), .ZN(n579) );
  NOR2_X1 U497 ( .A1(n598), .A2(n579), .ZN(n421) );
  NAND2_X1 U498 ( .A1(n490), .A2(n421), .ZN(n422) );
  XOR2_X1 U499 ( .A(KEYINPUT22), .B(n422), .Z(n499) );
  XNOR2_X1 U500 ( .A(n423), .B(G137), .ZN(n424) );
  XNOR2_X1 U501 ( .A(n425), .B(n424), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n442), .B(n426), .ZN(n708) );
  NAND2_X1 U503 ( .A1(n711), .A2(G227), .ZN(n427) );
  XNOR2_X1 U504 ( .A(n427), .B(G146), .ZN(n428) );
  XNOR2_X1 U505 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U506 ( .A(n708), .B(n430), .ZN(n696) );
  XNOR2_X1 U507 ( .A(KEYINPUT70), .B(G469), .ZN(n431) );
  XNOR2_X2 U508 ( .A(n432), .B(n431), .ZN(n551) );
  XNOR2_X2 U509 ( .A(n551), .B(KEYINPUT1), .ZN(n586) );
  XNOR2_X1 U510 ( .A(n586), .B(KEYINPUT88), .ZN(n537) );
  NAND2_X1 U511 ( .A1(n433), .A2(G210), .ZN(n435) );
  XOR2_X1 U512 ( .A(KEYINPUT94), .B(G131), .Z(n434) );
  XNOR2_X1 U513 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U514 ( .A(n436), .B(G146), .Z(n440) );
  XNOR2_X1 U515 ( .A(G101), .B(KEYINPUT5), .ZN(n437) );
  XNOR2_X1 U516 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U517 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U518 ( .A(n442), .B(n441), .ZN(n660) );
  NAND2_X1 U519 ( .A1(n660), .A2(n443), .ZN(n444) );
  XNOR2_X2 U520 ( .A(n444), .B(G472), .ZN(n523) );
  INV_X1 U521 ( .A(KEYINPUT6), .ZN(n445) );
  XNOR2_X1 U522 ( .A(n523), .B(n445), .ZN(n530) );
  INV_X1 U523 ( .A(KEYINPUT23), .ZN(n446) );
  NAND2_X1 U524 ( .A1(KEYINPUT79), .A2(n446), .ZN(n449) );
  INV_X1 U525 ( .A(KEYINPUT79), .ZN(n447) );
  NAND2_X1 U526 ( .A1(n447), .A2(KEYINPUT23), .ZN(n448) );
  NAND2_X1 U527 ( .A1(n449), .A2(n448), .ZN(n451) );
  XNOR2_X1 U528 ( .A(G110), .B(KEYINPUT24), .ZN(n450) );
  XOR2_X1 U529 ( .A(G140), .B(G137), .Z(n453) );
  XNOR2_X1 U530 ( .A(G119), .B(G128), .ZN(n452) );
  XNOR2_X1 U531 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U532 ( .A(n353), .B(n454), .ZN(n457) );
  NAND2_X1 U533 ( .A1(G221), .A2(n455), .ZN(n456) );
  XNOR2_X1 U534 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U535 ( .A(n709), .B(n458), .ZN(n704) );
  NOR2_X1 U536 ( .A1(n704), .A2(G902), .ZN(n462) );
  NAND2_X1 U537 ( .A1(n459), .A2(G217), .ZN(n460) );
  XNOR2_X1 U538 ( .A(n522), .B(KEYINPUT104), .ZN(n581) );
  NOR2_X1 U539 ( .A1(n530), .A2(n581), .ZN(n463) );
  AND2_X1 U540 ( .A1(n537), .A2(n463), .ZN(n464) );
  AND2_X1 U541 ( .A1(n499), .A2(n464), .ZN(n466) );
  XNOR2_X1 U542 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n465) );
  INV_X1 U543 ( .A(n499), .ZN(n469) );
  INV_X1 U544 ( .A(n586), .ZN(n473) );
  NOR2_X1 U545 ( .A1(n523), .A2(n522), .ZN(n467) );
  NAND2_X1 U546 ( .A1(n473), .A2(n467), .ZN(n468) );
  NOR2_X1 U547 ( .A1(n469), .A2(n468), .ZN(n622) );
  INV_X1 U548 ( .A(KEYINPUT83), .ZN(n470) );
  XNOR2_X1 U549 ( .A(n471), .B(n470), .ZN(n483) );
  INV_X1 U550 ( .A(n522), .ZN(n472) );
  INV_X1 U551 ( .A(n509), .ZN(n585) );
  NAND2_X1 U552 ( .A1(n530), .A2(n585), .ZN(n474) );
  XNOR2_X1 U553 ( .A(KEYINPUT86), .B(KEYINPUT33), .ZN(n475) );
  XNOR2_X1 U554 ( .A(n475), .B(KEYINPUT71), .ZN(n476) );
  INV_X1 U555 ( .A(n490), .ZN(n478) );
  XNOR2_X1 U556 ( .A(n479), .B(KEYINPUT34), .ZN(n481) );
  NOR2_X1 U557 ( .A1(n555), .A2(n548), .ZN(n480) );
  NAND2_X1 U558 ( .A1(n481), .A2(n480), .ZN(n482) );
  XOR2_X1 U559 ( .A(KEYINPUT35), .B(n482), .Z(n667) );
  NAND2_X1 U560 ( .A1(n483), .A2(n667), .ZN(n484) );
  XNOR2_X1 U561 ( .A(n484), .B(KEYINPUT44), .ZN(n502) );
  AND2_X1 U562 ( .A1(n523), .A2(n585), .ZN(n485) );
  AND2_X1 U563 ( .A1(n586), .A2(n485), .ZN(n591) );
  NAND2_X1 U564 ( .A1(n490), .A2(n591), .ZN(n486) );
  XNOR2_X1 U565 ( .A(n486), .B(KEYINPUT31), .ZN(n687) );
  INV_X1 U566 ( .A(n551), .ZN(n488) );
  INV_X1 U567 ( .A(n523), .ZN(n584) );
  NAND2_X1 U568 ( .A1(n584), .A2(n585), .ZN(n487) );
  NOR2_X1 U569 ( .A1(n488), .A2(n487), .ZN(n489) );
  NAND2_X1 U570 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U571 ( .A(KEYINPUT95), .B(n491), .ZN(n673) );
  NOR2_X1 U572 ( .A1(n687), .A2(n673), .ZN(n492) );
  XNOR2_X1 U573 ( .A(n492), .B(KEYINPUT96), .ZN(n494) );
  NAND2_X1 U574 ( .A1(n493), .A2(n548), .ZN(n533) );
  INV_X1 U575 ( .A(n533), .ZN(n683) );
  NOR2_X1 U576 ( .A1(n548), .A2(n493), .ZN(n686) );
  NOR2_X1 U577 ( .A1(n683), .A2(n686), .ZN(n600) );
  NOR2_X1 U578 ( .A1(n494), .A2(n600), .ZN(n495) );
  XNOR2_X1 U579 ( .A(n495), .B(KEYINPUT103), .ZN(n500) );
  INV_X1 U580 ( .A(n530), .ZN(n496) );
  NAND2_X1 U581 ( .A1(n496), .A2(n581), .ZN(n497) );
  NOR2_X1 U582 ( .A1(n497), .A2(n586), .ZN(n498) );
  NAND2_X1 U583 ( .A1(n499), .A2(n498), .ZN(n668) );
  NAND2_X1 U584 ( .A1(n500), .A2(n668), .ZN(n501) );
  INV_X1 U585 ( .A(KEYINPUT40), .ZN(n516) );
  NOR2_X1 U586 ( .A1(n517), .A2(n584), .ZN(n504) );
  XOR2_X1 U587 ( .A(KEYINPUT30), .B(n504), .Z(n554) );
  XOR2_X1 U588 ( .A(n505), .B(KEYINPUT105), .Z(n506) );
  NOR2_X1 U589 ( .A1(G900), .A2(n506), .ZN(n507) );
  NOR2_X1 U590 ( .A1(n508), .A2(n507), .ZN(n556) );
  NOR2_X1 U591 ( .A1(n556), .A2(n509), .ZN(n510) );
  NAND2_X1 U592 ( .A1(n551), .A2(n510), .ZN(n511) );
  NOR2_X1 U593 ( .A1(n554), .A2(n511), .ZN(n513) );
  BUF_X1 U594 ( .A(n512), .Z(n572) );
  XNOR2_X1 U595 ( .A(n572), .B(KEYINPUT38), .ZN(n596) );
  NAND2_X1 U596 ( .A1(n513), .A2(n596), .ZN(n514) );
  NAND2_X1 U597 ( .A1(n568), .A2(n683), .ZN(n515) );
  XNOR2_X1 U598 ( .A(n516), .B(n515), .ZN(n721) );
  INV_X1 U599 ( .A(n517), .ZN(n595) );
  NAND2_X1 U600 ( .A1(n596), .A2(n595), .ZN(n601) );
  NOR2_X1 U601 ( .A1(n601), .A2(n598), .ZN(n519) );
  XNOR2_X1 U602 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n518) );
  XNOR2_X1 U603 ( .A(n519), .B(n518), .ZN(n612) );
  NOR2_X1 U604 ( .A1(n579), .A2(n556), .ZN(n520) );
  XNOR2_X1 U605 ( .A(n520), .B(KEYINPUT69), .ZN(n521) );
  NOR2_X1 U606 ( .A1(n522), .A2(n521), .ZN(n531) );
  AND2_X1 U607 ( .A1(n523), .A2(n531), .ZN(n524) );
  XNOR2_X1 U608 ( .A(n524), .B(KEYINPUT28), .ZN(n525) );
  NAND2_X1 U609 ( .A1(n525), .A2(n551), .ZN(n541) );
  NOR2_X1 U610 ( .A1(n612), .A2(n541), .ZN(n526) );
  XNOR2_X1 U611 ( .A(KEYINPUT42), .B(n526), .ZN(n720) );
  NOR2_X1 U612 ( .A1(n721), .A2(n720), .ZN(n528) );
  XNOR2_X1 U613 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n527) );
  XNOR2_X1 U614 ( .A(n528), .B(n527), .ZN(n564) );
  XNOR2_X1 U615 ( .A(KEYINPUT84), .B(KEYINPUT109), .ZN(n529) );
  XNOR2_X1 U616 ( .A(n529), .B(KEYINPUT36), .ZN(n536) );
  NAND2_X1 U617 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U618 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U619 ( .A1(n534), .A2(n595), .ZN(n569) );
  XOR2_X1 U620 ( .A(n536), .B(n535), .Z(n538) );
  NAND2_X1 U621 ( .A1(n538), .A2(n537), .ZN(n691) );
  XNOR2_X1 U622 ( .A(KEYINPUT82), .B(n691), .ZN(n547) );
  INV_X1 U623 ( .A(KEYINPUT47), .ZN(n543) );
  INV_X1 U624 ( .A(n539), .ZN(n540) );
  NOR2_X1 U625 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U626 ( .A(n542), .B(KEYINPUT76), .ZN(n680) );
  XNOR2_X1 U627 ( .A(n543), .B(n680), .ZN(n545) );
  NAND2_X1 U628 ( .A1(n543), .A2(n600), .ZN(n544) );
  NAND2_X1 U629 ( .A1(n545), .A2(n544), .ZN(n546) );
  INV_X1 U630 ( .A(n548), .ZN(n549) );
  NAND2_X1 U631 ( .A1(n549), .A2(n585), .ZN(n550) );
  NOR2_X1 U632 ( .A1(n550), .A2(n572), .ZN(n552) );
  NAND2_X1 U633 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U634 ( .A1(n554), .A2(n553), .ZN(n558) );
  NOR2_X1 U635 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U636 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U637 ( .A(KEYINPUT107), .B(n559), .ZN(n722) );
  NAND2_X1 U638 ( .A1(n600), .A2(KEYINPUT47), .ZN(n560) );
  XOR2_X1 U639 ( .A(KEYINPUT78), .B(n560), .Z(n561) );
  NOR2_X1 U640 ( .A1(n722), .A2(n561), .ZN(n562) );
  XOR2_X1 U641 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n565) );
  XNOR2_X1 U642 ( .A(KEYINPUT81), .B(n565), .ZN(n566) );
  XNOR2_X1 U643 ( .A(n567), .B(n566), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n568), .A2(n686), .ZN(n693) );
  INV_X1 U645 ( .A(n693), .ZN(n575) );
  NOR2_X1 U646 ( .A1(n569), .A2(n586), .ZN(n571) );
  XNOR2_X1 U647 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n570) );
  XNOR2_X1 U648 ( .A(n571), .B(n570), .ZN(n574) );
  INV_X1 U649 ( .A(n572), .ZN(n573) );
  NOR2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n621) );
  NOR2_X1 U651 ( .A1(n575), .A2(n621), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n642) );
  XNOR2_X1 U653 ( .A(n578), .B(KEYINPUT2), .ZN(n616) );
  INV_X1 U654 ( .A(n579), .ZN(n580) );
  NOR2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U656 ( .A(n582), .B(KEYINPUT49), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n587), .B(KEYINPUT50), .ZN(n588) );
  NOR2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U661 ( .A(KEYINPUT119), .B(n590), .Z(n592) );
  NOR2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U663 ( .A(KEYINPUT51), .B(n593), .Z(n594) );
  NOR2_X1 U664 ( .A1(n612), .A2(n594), .ZN(n606) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U667 ( .A(n599), .B(KEYINPUT120), .ZN(n603) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U670 ( .A1(n604), .A2(n611), .ZN(n605) );
  NOR2_X1 U671 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U672 ( .A(n607), .B(KEYINPUT52), .ZN(n608) );
  NOR2_X1 U673 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U674 ( .A(KEYINPUT121), .B(n610), .ZN(n614) );
  NOR2_X1 U675 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U676 ( .A1(n711), .A2(n617), .ZN(n619) );
  XNOR2_X1 U677 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n618) );
  XNOR2_X1 U678 ( .A(n621), .B(n620), .ZN(G42) );
  XOR2_X1 U679 ( .A(G110), .B(n622), .Z(G12) );
  NOR2_X1 U680 ( .A1(n623), .A2(G953), .ZN(n624) );
  XNOR2_X1 U681 ( .A(n624), .B(KEYINPUT125), .ZN(n628) );
  NAND2_X1 U682 ( .A1(G953), .A2(G224), .ZN(n625) );
  XNOR2_X1 U683 ( .A(KEYINPUT61), .B(n625), .ZN(n626) );
  NAND2_X1 U684 ( .A1(n626), .A2(G898), .ZN(n627) );
  NAND2_X1 U685 ( .A1(n628), .A2(n627), .ZN(n633) );
  INV_X1 U686 ( .A(n629), .ZN(n631) );
  NOR2_X1 U687 ( .A1(G898), .A2(n711), .ZN(n630) );
  NOR2_X1 U688 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U689 ( .A(n633), .B(n632), .ZN(G69) );
  INV_X1 U690 ( .A(n644), .ZN(n636) );
  XNOR2_X1 U691 ( .A(n642), .B(KEYINPUT74), .ZN(n634) );
  NOR2_X1 U692 ( .A1(n634), .A2(n637), .ZN(n635) );
  NAND2_X1 U693 ( .A1(n636), .A2(n635), .ZN(n640) );
  XOR2_X1 U694 ( .A(KEYINPUT80), .B(n637), .Z(n638) );
  NAND2_X1 U695 ( .A1(n638), .A2(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U696 ( .A1(n640), .A2(n639), .ZN(n646) );
  INV_X1 U697 ( .A(KEYINPUT2), .ZN(n641) );
  OR2_X1 U698 ( .A1(n642), .A2(n641), .ZN(n643) );
  OR2_X1 U699 ( .A1(n644), .A2(n643), .ZN(n645) );
  AND2_X2 U700 ( .A1(n646), .A2(n645), .ZN(n700) );
  NAND2_X1 U701 ( .A1(n700), .A2(G475), .ZN(n649) );
  XNOR2_X1 U702 ( .A(n647), .B(KEYINPUT59), .ZN(n648) );
  XNOR2_X1 U703 ( .A(n649), .B(n648), .ZN(n651) );
  INV_X1 U704 ( .A(G952), .ZN(n650) );
  XNOR2_X1 U705 ( .A(n652), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U706 ( .A1(n700), .A2(G210), .ZN(n656) );
  XNOR2_X1 U707 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n653) );
  XNOR2_X1 U708 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U709 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U710 ( .A(n658), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U711 ( .A1(n700), .A2(G472), .ZN(n662) );
  XNOR2_X1 U712 ( .A(KEYINPUT87), .B(KEYINPUT62), .ZN(n659) );
  XNOR2_X1 U713 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U714 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U715 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n664) );
  XNOR2_X1 U716 ( .A(n665), .B(n664), .ZN(G57) );
  XOR2_X1 U717 ( .A(G119), .B(n666), .Z(G21) );
  XNOR2_X1 U718 ( .A(n667), .B(G122), .ZN(G24) );
  XNOR2_X1 U719 ( .A(n668), .B(G101), .ZN(n669) );
  XNOR2_X1 U720 ( .A(KEYINPUT110), .B(n669), .ZN(G3) );
  NAND2_X1 U721 ( .A1(n673), .A2(n683), .ZN(n670) );
  XNOR2_X1 U722 ( .A(n670), .B(G104), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n672) );
  XNOR2_X1 U724 ( .A(KEYINPUT111), .B(KEYINPUT27), .ZN(n671) );
  XNOR2_X1 U725 ( .A(n672), .B(n671), .ZN(n677) );
  XNOR2_X1 U726 ( .A(G107), .B(KEYINPUT26), .ZN(n675) );
  NAND2_X1 U727 ( .A1(n686), .A2(n673), .ZN(n674) );
  XNOR2_X1 U728 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U729 ( .A(n677), .B(n676), .ZN(G9) );
  XOR2_X1 U730 ( .A(G128), .B(KEYINPUT29), .Z(n679) );
  NAND2_X1 U731 ( .A1(n686), .A2(n680), .ZN(n678) );
  XNOR2_X1 U732 ( .A(n679), .B(n678), .ZN(G30) );
  XOR2_X1 U733 ( .A(G146), .B(KEYINPUT115), .Z(n682) );
  NAND2_X1 U734 ( .A1(n683), .A2(n680), .ZN(n681) );
  XNOR2_X1 U735 ( .A(n682), .B(n681), .ZN(G48) );
  NAND2_X1 U736 ( .A1(n687), .A2(n683), .ZN(n684) );
  XNOR2_X1 U737 ( .A(n684), .B(KEYINPUT116), .ZN(n685) );
  XNOR2_X1 U738 ( .A(G113), .B(n685), .ZN(G15) );
  XOR2_X1 U739 ( .A(G116), .B(KEYINPUT117), .Z(n689) );
  NAND2_X1 U740 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U741 ( .A(n689), .B(n688), .ZN(G18) );
  XOR2_X1 U742 ( .A(KEYINPUT118), .B(KEYINPUT37), .Z(n690) );
  XNOR2_X1 U743 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U744 ( .A(G125), .B(n692), .ZN(G27) );
  XNOR2_X1 U745 ( .A(G134), .B(n693), .ZN(G36) );
  NAND2_X1 U746 ( .A1(n700), .A2(G469), .ZN(n698) );
  XOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XNOR2_X1 U748 ( .A(n694), .B(KEYINPUT124), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U750 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U751 ( .A1(n707), .A2(n699), .ZN(G54) );
  NAND2_X1 U752 ( .A1(n700), .A2(G478), .ZN(n701) );
  XOR2_X1 U753 ( .A(n702), .B(n701), .Z(n703) );
  NOR2_X1 U754 ( .A1(n707), .A2(n703), .ZN(G63) );
  NAND2_X1 U755 ( .A1(n700), .A2(G217), .ZN(n705) );
  XNOR2_X1 U756 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U757 ( .A1(n707), .A2(n706), .ZN(G66) );
  XOR2_X1 U758 ( .A(n709), .B(n708), .Z(n713) );
  XNOR2_X1 U759 ( .A(n710), .B(n713), .ZN(n712) );
  NAND2_X1 U760 ( .A1(n712), .A2(n711), .ZN(n718) );
  XNOR2_X1 U761 ( .A(n713), .B(G227), .ZN(n714) );
  XNOR2_X1 U762 ( .A(n714), .B(KEYINPUT126), .ZN(n715) );
  NAND2_X1 U763 ( .A1(n715), .A2(G900), .ZN(n716) );
  NAND2_X1 U764 ( .A1(n716), .A2(G953), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U766 ( .A(KEYINPUT127), .B(n719), .Z(G72) );
  XOR2_X1 U767 ( .A(G137), .B(n720), .Z(G39) );
  XOR2_X1 U768 ( .A(n721), .B(G131), .Z(G33) );
  XOR2_X1 U769 ( .A(G143), .B(n722), .Z(n723) );
  XNOR2_X1 U770 ( .A(KEYINPUT114), .B(n723), .ZN(G45) );
endmodule

