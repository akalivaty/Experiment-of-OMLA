//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT77), .Z(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n193), .A2(new_n194), .A3(G107), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(G104), .A2(G107), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT79), .B(G107), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G104), .ZN(new_n199));
  OAI211_X1 g013(.A(G101), .B(new_n196), .C1(new_n199), .C2(KEYINPUT3), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT80), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT79), .A2(G107), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT79), .A2(G107), .ZN(new_n203));
  OAI21_X1  g017(.A(G104), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n197), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n193), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G101), .A4(new_n196), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT3), .B1(new_n204), .B2(new_n205), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(new_n195), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n209), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G143), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  OR2_X1    g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n218), .B1(new_n221), .B2(new_n219), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n200), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n213), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G137), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(G137), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  INV_X1    g049(.A(G131), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n233), .A3(new_n236), .A4(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(KEYINPUT82), .B(new_n194), .C1(new_n202), .C2(new_n203), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n194), .B2(G107), .ZN(new_n242));
  INV_X1    g056(.A(G107), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT81), .A3(G104), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT82), .B1(new_n198), .B2(new_n194), .ZN(new_n247));
  OAI21_X1  g061(.A(G101), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n212), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n215), .A2(new_n217), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(KEYINPUT65), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n215), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g070(.A1(KEYINPUT66), .A2(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT66), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n251), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(KEYINPUT65), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n252), .A2(KEYINPUT1), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n218), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n250), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n251), .A2(G128), .A3(new_n261), .A4(new_n262), .ZN(new_n267));
  AND2_X1   g081(.A1(KEYINPUT66), .A2(G128), .ZN(new_n268));
  NOR2_X1   g082(.A1(KEYINPUT66), .A2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n215), .B2(new_n263), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n267), .B(KEYINPUT68), .C1(new_n271), .C2(new_n251), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n249), .A2(KEYINPUT10), .A3(new_n266), .A4(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n217), .A2(new_n254), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(new_n264), .B2(new_n218), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n212), .A2(new_n248), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n227), .A2(new_n239), .A3(new_n273), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT84), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n266), .A2(new_n272), .A3(KEYINPUT10), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n282), .A2(new_n249), .B1(new_n277), .B2(new_n278), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT84), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n239), .A4(new_n227), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT86), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n227), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(new_n238), .ZN(new_n289));
  AOI211_X1 g103(.A(KEYINPUT86), .B(new_n239), .C1(new_n283), .C2(new_n227), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(G110), .B(G140), .Z(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT78), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G227), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n293), .B(new_n295), .Z(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n267), .B1(new_n271), .B2(new_n251), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n277), .B1(new_n249), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n238), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT12), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n286), .A2(new_n303), .A3(new_n296), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n192), .B1(new_n305), .B2(new_n190), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n286), .A2(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n297), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT85), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n286), .A2(new_n309), .A3(new_n296), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n213), .A2(new_n226), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n212), .A2(new_n248), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n266), .A2(new_n272), .A3(KEYINPUT10), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n279), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n238), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT86), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n288), .A2(new_n287), .A3(new_n238), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n297), .B1(new_n281), .B2(new_n285), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(new_n309), .ZN(new_n321));
  OAI211_X1 g135(.A(G469), .B(new_n308), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n189), .B1(new_n306), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT67), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G119), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(G128), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n257), .A2(KEYINPUT23), .A3(G119), .A4(new_n258), .ZN(new_n329));
  AOI21_X1  g143(.A(G128), .B1(new_n325), .B2(new_n327), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G110), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT71), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT16), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(G125), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(G146), .B(new_n336), .C1(new_n340), .C2(new_n334), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT72), .ZN(new_n342));
  XNOR2_X1  g156(.A(G125), .B(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G146), .A4(new_n336), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n336), .B1(new_n340), .B2(new_n334), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n214), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n325), .A2(new_n327), .A3(G128), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n268), .A2(new_n269), .A3(new_n324), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT24), .B(G110), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT71), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n331), .A2(new_n356), .A3(G110), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n333), .A2(new_n349), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT73), .B(G110), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n331), .A2(new_n359), .B1(new_n352), .B2(new_n354), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n343), .A2(new_n214), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n341), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n360), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n360), .B2(new_n362), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n358), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT75), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G137), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n358), .B(KEYINPUT76), .C1(new_n364), .C2(new_n365), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n368), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n366), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT76), .A3(new_n372), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G217), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(G234), .B2(new_n191), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT25), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n383), .A3(new_n191), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n380), .ZN(new_n385));
  AOI21_X1  g199(.A(G902), .B1(new_n375), .B2(new_n377), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n383), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n382), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n231), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n229), .A2(G137), .ZN(new_n390));
  OAI21_X1  g204(.A(G131), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n391), .A2(new_n237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n266), .A2(new_n272), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n325), .A2(new_n327), .A3(G116), .ZN(new_n394));
  INV_X1    g208(.A(G116), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G119), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT2), .B(G113), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n399), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n220), .A2(new_n222), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n238), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n393), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT28), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n393), .A2(new_n406), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n403), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n407), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n412), .B2(KEYINPUT28), .ZN(new_n413));
  NOR2_X1   g227(.A1(G237), .A2(G953), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G210), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT27), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT26), .B(G101), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n299), .A2(new_n392), .ZN(new_n423));
  INV_X1    g237(.A(new_n406), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n403), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n408), .B1(new_n425), .B2(new_n407), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n418), .B(KEYINPUT69), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n426), .A2(new_n409), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n423), .B2(new_n424), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n393), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n403), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n407), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n419), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n420), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n422), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G472), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n433), .A2(new_n407), .A3(new_n418), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT31), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT31), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n433), .A2(new_n441), .A3(new_n407), .A4(new_n418), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n428), .B1(new_n426), .B2(new_n409), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G472), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n191), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT70), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT32), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT32), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n388), .B1(new_n438), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G214), .B1(G237), .B2(G902), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G122), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n403), .B1(KEYINPUT4), .B2(new_n200), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n195), .B1(new_n206), .B2(new_n193), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n208), .B1(new_n460), .B2(G101), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n462), .B2(new_n209), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT5), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n325), .A2(new_n327), .A3(new_n464), .A4(G116), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n465), .A2(G113), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n394), .A2(KEYINPUT5), .A3(new_n396), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n401), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT87), .B1(new_n312), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n466), .A2(new_n467), .B1(new_n398), .B2(new_n400), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n212), .A4(new_n248), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n457), .B1(new_n463), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n224), .A2(new_n225), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n213), .A2(new_n403), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n477), .A2(new_n470), .A3(new_n473), .A4(new_n456), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n475), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT88), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n475), .A2(new_n481), .A3(new_n478), .A4(KEYINPUT6), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n475), .A2(KEYINPUT6), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n299), .A2(new_n338), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n405), .A2(G125), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n294), .A2(G224), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n486), .B(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n480), .A2(new_n482), .A3(new_n483), .A4(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n312), .B(new_n469), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n456), .B(KEYINPUT8), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT89), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n488), .A2(KEYINPUT7), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT90), .B1(new_n486), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n484), .A2(new_n498), .A3(new_n485), .A4(new_n495), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n497), .A2(new_n499), .B1(new_n486), .B2(new_n496), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n500), .A2(new_n478), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n490), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G210), .B1(G237), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n490), .A2(new_n504), .A3(new_n502), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n455), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT101), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(G104), .ZN(new_n511));
  INV_X1    g325(.A(G237), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n294), .A3(G214), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n216), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n414), .A2(G143), .A3(G214), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT18), .A2(G131), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT91), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n516), .A2(new_n520), .A3(KEYINPUT18), .A4(G131), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n340), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n343), .A2(KEYINPUT92), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(G146), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n526), .A2(new_n361), .B1(new_n517), .B2(new_n518), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT19), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n343), .A2(KEYINPUT19), .ZN(new_n531));
  AOI21_X1  g345(.A(G146), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n516), .A2(G131), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n514), .A2(new_n236), .A3(new_n515), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n341), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n511), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n349), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n533), .A2(new_n540), .A3(new_n534), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n516), .A2(KEYINPUT17), .A3(G131), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n533), .A2(KEYINPUT94), .A3(new_n540), .A4(new_n534), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n539), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n522), .A2(new_n527), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n511), .B(KEYINPUT93), .Z(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(G475), .A2(G902), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT20), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT20), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n554), .A3(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n546), .A2(new_n547), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n511), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n549), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n191), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G475), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n264), .A2(G143), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n259), .B2(new_n216), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G134), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n270), .B2(G143), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(new_n229), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT97), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G122), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G116), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n395), .A2(G122), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT95), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n198), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n395), .A2(G122), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n571), .B1(new_n577), .B2(KEYINPUT14), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(KEYINPUT14), .B2(new_n571), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(G107), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n564), .A2(G134), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n566), .A2(new_n229), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n568), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n198), .ZN(new_n586));
  INV_X1    g400(.A(new_n575), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n574), .B1(new_n570), .B2(new_n571), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n573), .A2(new_n198), .A3(new_n575), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT13), .B(new_n563), .C1(new_n259), .C2(new_n216), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n229), .B1(new_n562), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n592), .A2(new_n594), .B1(new_n566), .B2(new_n229), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n591), .B2(new_n595), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n585), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n187), .A2(new_n379), .A3(G953), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT98), .Z(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n601), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n585), .B(new_n603), .C1(new_n597), .C2(new_n598), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(KEYINPUT100), .A3(new_n191), .ZN(new_n606));
  INV_X1    g420(.A(G478), .ZN(new_n607));
  NOR2_X1   g421(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n611), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n605), .A2(KEYINPUT100), .A3(new_n191), .A4(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n556), .A2(new_n561), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(G234), .A2(G237), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(G952), .A3(new_n294), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT21), .B(G898), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(G902), .A3(G953), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n509), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n612), .A2(new_n614), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n553), .A2(new_n555), .B1(new_n560), .B2(G475), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(KEYINPUT101), .A3(new_n621), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n323), .A2(new_n453), .A3(new_n508), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  AOI21_X1  g444(.A(new_n296), .B1(new_n318), .B2(new_n286), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n286), .A2(new_n296), .A3(new_n303), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n190), .B(new_n191), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n192), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n322), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n189), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n444), .A2(new_n191), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G472), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n448), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n637), .A2(new_n388), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n490), .A2(new_n504), .A3(new_n502), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n504), .B1(new_n490), .B2(new_n502), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n454), .B(new_n621), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n645), .B1(new_n605), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n602), .A2(KEYINPUT103), .A3(KEYINPUT33), .A4(new_n604), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT102), .B1(new_n605), .B2(new_n646), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n650));
  AOI211_X1 g464(.A(new_n650), .B(KEYINPUT33), .C1(new_n602), .C2(new_n604), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(G478), .B1(new_n652), .B2(G902), .ZN(new_n653));
  INV_X1    g467(.A(new_n626), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n605), .A2(new_n607), .A3(new_n191), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n644), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n641), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT104), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  NAND3_X1  g475(.A1(new_n624), .A2(new_n626), .A3(new_n621), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT105), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n641), .A2(new_n508), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  INV_X1    g480(.A(new_n381), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n372), .A2(KEYINPUT36), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n366), .B(new_n668), .Z(new_n669));
  OAI22_X1  g483(.A1(new_n385), .A2(new_n387), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT106), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n667), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n386), .A2(new_n383), .ZN(new_n673));
  INV_X1    g487(.A(new_n380), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n386), .B2(new_n383), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n672), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n640), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n628), .A2(new_n636), .A3(new_n635), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n508), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  NAND2_X1  g498(.A1(new_n506), .A2(new_n507), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n671), .A3(new_n678), .A4(new_n454), .ZN(new_n686));
  INV_X1    g500(.A(new_n451), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n450), .B1(new_n444), .B2(new_n447), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n438), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n624), .A2(new_n626), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n617), .B(KEYINPUT107), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(G900), .B2(new_n620), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n635), .A2(new_n689), .A3(new_n636), .A4(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n686), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n264), .ZN(G30));
  XNOR2_X1  g511(.A(new_n692), .B(KEYINPUT39), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n635), .A2(new_n636), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n635), .A2(KEYINPUT108), .A3(new_n636), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT40), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT40), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n701), .A2(new_n705), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n412), .A2(new_n428), .ZN(new_n707));
  AOI21_X1  g521(.A(G902), .B1(new_n707), .B2(new_n439), .ZN(new_n708));
  OAI22_X1  g522(.A1(new_n687), .A2(new_n688), .B1(new_n445), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n625), .A2(new_n626), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n454), .A3(new_n676), .A4(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n685), .A2(KEYINPUT38), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n685), .A2(KEYINPUT38), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n704), .A2(new_n706), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  NAND4_X1  g530(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n692), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n689), .A3(new_n636), .A4(new_n635), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n686), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n214), .ZN(G48));
  AOI22_X1  g535(.A1(new_n291), .A2(new_n297), .B1(new_n303), .B2(new_n320), .ZN(new_n722));
  OAI21_X1  g536(.A(G469), .B1(new_n722), .B2(G902), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n636), .A3(new_n633), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n657), .A2(new_n453), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n725), .A2(new_n663), .A3(new_n453), .A4(new_n508), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NAND4_X1  g544(.A1(new_n628), .A2(new_n671), .A3(new_n678), .A4(new_n689), .ZN(new_n731));
  INV_X1    g545(.A(new_n633), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n316), .A2(new_n317), .B1(new_n281), .B2(new_n285), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n304), .B1(new_n733), .B2(new_n296), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n190), .B1(new_n734), .B2(new_n191), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n508), .A3(KEYINPUT109), .A4(new_n636), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n454), .B1(new_n642), .B2(new_n643), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n738), .B1(new_n724), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n731), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n324), .ZN(G21));
  AND4_X1   g556(.A1(new_n636), .A2(new_n723), .A3(new_n633), .A4(new_n621), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n454), .B(new_n710), .C1(new_n642), .C2(new_n643), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n440), .B(new_n442), .C1(new_n427), .C2(new_n413), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n447), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n639), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n388), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n743), .A2(new_n745), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n676), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n718), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n737), .B2(new_n740), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n338), .ZN(G27));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n642), .A2(new_n643), .A3(new_n455), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n453), .A2(new_n757), .A3(new_n636), .A4(new_n635), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n758), .B2(new_n717), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n506), .A2(new_n454), .A3(new_n507), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n637), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .A3(new_n453), .A4(new_n718), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NOR3_X1   g578(.A1(new_n758), .A2(new_n690), .A3(new_n693), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n229), .ZN(G36));
  OAI21_X1  g580(.A(new_n308), .B1(new_n319), .B2(new_n321), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT45), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n769), .B(new_n308), .C1(new_n319), .C2(new_n321), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(G469), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n634), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(G469), .C1(new_n771), .C2(G902), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n633), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n636), .A3(new_n698), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT110), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n776), .A2(new_n779), .A3(new_n636), .A4(new_n698), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n653), .A2(new_n626), .A3(new_n655), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT43), .B1(new_n781), .B2(KEYINPUT111), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n670), .A2(new_n640), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT44), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n784), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(KEYINPUT44), .A3(new_n782), .A4(new_n786), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n757), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n778), .A2(new_n780), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  INV_X1    g607(.A(new_n388), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n760), .A2(new_n717), .A3(new_n794), .A4(new_n689), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n776), .A2(KEYINPUT47), .A3(new_n636), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT47), .B1(new_n776), .B2(new_n636), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NOR2_X1   g613(.A1(G952), .A2(G953), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT117), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n783), .A2(new_n784), .A3(new_n691), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n724), .A2(new_n760), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n453), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT48), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n709), .A2(new_n388), .A3(new_n617), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(G952), .B(new_n294), .C1(new_n807), .C2(new_n656), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n802), .A2(new_n749), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n737), .A2(new_n740), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n712), .A2(new_n713), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n455), .A3(new_n725), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n809), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT50), .B1(new_n817), .B2(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n817), .A2(KEYINPUT50), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n817), .B2(KEYINPUT50), .ZN(new_n822));
  OAI22_X1  g636(.A1(new_n815), .A2(new_n809), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n802), .A2(new_n752), .A3(new_n803), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n803), .A2(new_n806), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n819), .A2(new_n823), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n810), .A2(new_n757), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT114), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n796), .A2(new_n797), .ZN(new_n830));
  INV_X1    g644(.A(new_n736), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n636), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n827), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n813), .B1(new_n833), .B2(KEYINPUT51), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(KEYINPUT51), .B2(new_n833), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n765), .B1(new_n762), .B2(new_n759), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n629), .A2(new_n729), .A3(new_n750), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n741), .ZN(new_n839));
  INV_X1    g653(.A(new_n644), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n388), .A2(new_n640), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n656), .A2(new_n690), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n323), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n682), .A2(new_n726), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n615), .A2(new_n693), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n671), .A2(new_n678), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n635), .A2(new_n689), .A3(new_n636), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n846), .A2(new_n847), .A3(new_n760), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n757), .A2(new_n636), .A3(new_n635), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n753), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n717), .A2(new_n676), .A3(new_n748), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n761), .A2(KEYINPUT112), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n848), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n837), .A2(new_n839), .A3(new_n844), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n696), .B1(new_n811), .B2(new_n852), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n693), .B(new_n672), .C1(new_n673), .C2(new_n675), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n635), .A2(new_n857), .A3(new_n709), .A4(new_n636), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n744), .ZN(new_n859));
  INV_X1    g673(.A(new_n686), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n847), .A2(new_n717), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n862), .A3(KEYINPUT52), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT52), .B1(new_n856), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n863), .B1(new_n864), .B2(KEYINPUT113), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n866), .B(KEYINPUT52), .C1(new_n856), .C2(new_n862), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n836), .B(new_n855), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n719), .A2(new_n686), .B1(new_n744), .B2(new_n858), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n869), .A2(new_n754), .A3(new_n870), .A4(new_n696), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n864), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n837), .A2(new_n839), .A3(new_n844), .A4(new_n854), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT53), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(KEYINPUT54), .A3(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(KEYINPUT53), .B(new_n855), .C1(new_n865), .C2(new_n867), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n836), .B1(new_n872), .B2(new_n873), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n801), .B1(new_n835), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n736), .B(KEYINPUT49), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n794), .A2(new_n454), .A3(new_n636), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n883), .A2(new_n781), .A3(new_n709), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n814), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n881), .A2(new_n885), .ZN(G75));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n876), .A2(new_n878), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(G902), .ZN(new_n889));
  INV_X1    g703(.A(G210), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT118), .Z(new_n893));
  XOR2_X1   g707(.A(new_n489), .B(KEYINPUT55), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n887), .B(new_n895), .C1(new_n889), .C2(new_n890), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n294), .A2(G952), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT119), .Z(new_n900));
  AND3_X1   g714(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(G51));
  INV_X1    g715(.A(new_n900), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n192), .B(KEYINPUT57), .ZN(new_n903));
  INV_X1    g717(.A(new_n879), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n734), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n889), .A2(new_n772), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n902), .B1(new_n907), .B2(new_n908), .ZN(G54));
  NAND2_X1  g723(.A1(KEYINPUT58), .A2(G475), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n889), .A2(new_n550), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n550), .B1(new_n889), .B2(new_n910), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n902), .B1(new_n911), .B2(new_n912), .ZN(G60));
  XNOR2_X1  g727(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n607), .A2(new_n191), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n914), .B(new_n915), .Z(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n880), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n652), .B(KEYINPUT120), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(KEYINPUT122), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n879), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n920), .A2(new_n916), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n902), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n916), .B1(new_n875), .B2(new_n879), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n919), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n921), .A2(new_n925), .A3(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n876), .B2(new_n878), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n900), .B1(new_n933), .B2(new_n378), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n669), .B(new_n932), .C1(new_n876), .C2(new_n878), .ZN(new_n936));
  OR3_X1    g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(G66));
  NAND2_X1  g753(.A1(new_n839), .A2(new_n844), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n294), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n619), .A2(G224), .A3(G953), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT123), .ZN(new_n945));
  INV_X1    g759(.A(G898), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n893), .B1(new_n946), .B2(G953), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G69));
  NAND2_X1  g762(.A1(new_n431), .A2(new_n432), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n530), .A2(new_n531), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(G900), .B2(G953), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n754), .A2(new_n720), .A3(new_n696), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n837), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n798), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n778), .A2(new_n453), .A3(new_n745), .A4(new_n780), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n955), .A2(new_n792), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n957), .B2(G953), .ZN(new_n958));
  INV_X1    g772(.A(new_n951), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n704), .A2(new_n706), .A3(new_n714), .ZN(new_n961));
  INV_X1    g775(.A(new_n720), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n856), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n715), .A2(new_n953), .A3(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n703), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n967), .A2(new_n453), .A3(new_n757), .A4(new_n842), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n966), .A2(new_n792), .A3(new_n798), .A4(new_n968), .ZN(new_n969));
  AOI211_X1 g783(.A(KEYINPUT124), .B(new_n959), .C1(new_n969), .C2(new_n294), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n964), .A2(new_n965), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n792), .A2(new_n798), .A3(new_n968), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n294), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n971), .B1(new_n974), .B2(new_n951), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n958), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n977), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n979), .B(new_n958), .C1(new_n970), .C2(new_n975), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(G72));
  XNOR2_X1  g795(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n445), .A2(new_n191), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT126), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n969), .B2(new_n940), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n418), .A3(new_n434), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n984), .B1(new_n435), .B2(new_n439), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n868), .A2(new_n874), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n434), .A2(new_n418), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n955), .A2(new_n792), .A3(new_n941), .A4(new_n956), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n985), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n995));
  OR3_X1    g809(.A1(new_n994), .A2(new_n995), .A3(new_n902), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n994), .B2(new_n902), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(new_n996), .B2(new_n997), .ZN(G57));
endmodule


