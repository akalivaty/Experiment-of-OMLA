//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G221), .A4(G218), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n451), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n460), .A2(new_n461), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n462), .A2(G136), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n468), .B1(new_n460), .B2(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  MUX2_X1   g051(.A(G100), .B(G112), .S(G2105), .Z(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n462), .A2(new_n481), .A3(G138), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n468), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G102), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT69), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n487), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n503), .B1(new_n500), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G62), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n505), .B1(new_n504), .B2(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(G88), .B1(G50), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND2_X1  g093(.A1(new_n515), .A2(G51), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT72), .B(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n504), .A2(new_n511), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n515), .A2(G51), .B1(new_n525), .B2(new_n524), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n530), .A2(KEYINPUT73), .A3(new_n521), .A4(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n512), .A2(new_n536), .B1(new_n537), .B2(new_n514), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(G43), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n513), .A2(G81), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n534), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(G78), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT77), .B1(new_n553), .B2(new_n502), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n553), .A2(new_n502), .A3(KEYINPUT77), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n500), .A2(G543), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n502), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT70), .B1(new_n502), .B2(KEYINPUT5), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n554), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n514), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n511), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n561), .A2(G651), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n512), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n504), .A2(KEYINPUT76), .A3(new_n511), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(G91), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  NAND3_X1  g148(.A1(new_n568), .A2(G87), .A3(new_n569), .ZN(new_n574));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n559), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n511), .A2(G49), .A3(G543), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n511), .A2(KEYINPUT78), .A3(G49), .A4(G543), .ZN(new_n580));
  AOI22_X1  g155(.A1(G651), .A2(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n574), .A2(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n568), .A2(G86), .A3(new_n569), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n559), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n515), .A2(G48), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n534), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n512), .A2(new_n592), .B1(new_n593), .B2(new_n514), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NOR2_X1   g172(.A1(G301), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n515), .A2(G54), .ZN(new_n599));
  OAI211_X1 g174(.A(G66), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n600), .A2(KEYINPUT80), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT80), .B1(new_n600), .B2(new_n601), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n600), .A2(new_n601), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n609), .A2(G651), .A3(new_n602), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n610), .A2(new_n611), .A3(new_n599), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n568), .A2(G92), .A3(new_n569), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n568), .A2(G92), .A3(new_n569), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n613), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n606), .A2(new_n612), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n598), .B1(new_n618), .B2(new_n597), .ZN(G284));
  XNOR2_X1  g194(.A(G284), .B(KEYINPUT82), .ZN(G321));
  NOR2_X1   g195(.A1(G168), .A2(new_n597), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT83), .B1(G299), .B2(new_n597), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n621), .B2(new_n624), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(new_n621), .B2(new_n624), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n618), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n617), .A2(new_n615), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n605), .A2(KEYINPUT81), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n611), .B1(new_n610), .B2(new_n599), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n627), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(KEYINPUT84), .B1(new_n618), .B2(new_n627), .ZN(new_n635));
  OAI21_X1  g210(.A(G868), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n462), .A2(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  MUX2_X1   g219(.A(G99), .B(G111), .S(G2105), .Z(new_n645));
  AOI22_X1  g220(.A1(G123), .A2(new_n475), .B1(new_n645), .B2(G2104), .ZN(new_n646));
  INV_X1    g221(.A(G135), .ZN(new_n647));
  INV_X1    g222(.A(new_n462), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n643), .A2(new_n644), .A3(new_n651), .ZN(G156));
  XOR2_X1   g227(.A(KEYINPUT15), .B(G2435), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT87), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT86), .B(G2438), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1341), .B(G1348), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G14), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n661), .B2(new_n667), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2072), .B(G2078), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n675), .B(KEYINPUT17), .Z(new_n678));
  INV_X1    g253(.A(new_n673), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(new_n674), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n675), .B(KEYINPUT88), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n679), .B1(new_n682), .B2(new_n674), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(KEYINPUT89), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n686));
  INV_X1    g261(.A(new_n674), .ZN(new_n687));
  OAI22_X1  g262(.A1(new_n683), .A2(new_n686), .B1(new_n687), .B2(new_n678), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n681), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(new_n650), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G2100), .ZN(G227));
  XOR2_X1   g266(.A(G1971), .B(G1976), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1956), .B(G2474), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1961), .B(G1966), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(new_n696), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT20), .Z(new_n700));
  AOI211_X1 g275(.A(new_n698), .B(new_n700), .C1(new_n693), .C2(new_n697), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n704), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  NOR2_X1   g284(.A1(G16), .A2(G21), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G168), .B2(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G1966), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT102), .ZN(new_n713));
  NAND2_X1  g288(.A1(G160), .A2(G29), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  AND2_X1   g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  NOR2_X1   g291(.A1(KEYINPUT24), .A2(G34), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT101), .ZN(new_n720));
  INV_X1    g295(.A(G2084), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G27), .A2(G29), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G164), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G2078), .Z(new_n725));
  INV_X1    g300(.A(G1961), .ZN(new_n726));
  NOR2_X1   g301(.A1(G5), .A2(G16), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G171), .B2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT104), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n722), .B(new_n725), .C1(new_n726), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G19), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n545), .B2(G16), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1341), .Z(new_n733));
  NOR2_X1   g308(.A1(G29), .A2(G33), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT100), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n465), .A2(G103), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n462), .A2(G139), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n737), .B(new_n738), .C1(new_n468), .C2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n735), .B1(new_n740), .B2(new_n715), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2072), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT26), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G105), .B2(new_n465), .ZN(new_n745));
  AOI22_X1  g320(.A1(G129), .A2(new_n475), .B1(new_n462), .B2(G141), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n715), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n715), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT103), .B(G28), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT30), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(new_n715), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n755), .B(new_n756), .C1(new_n649), .C2(new_n715), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n750), .B2(new_n751), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n733), .A2(new_n742), .A3(new_n752), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT29), .ZN(new_n762));
  INV_X1    g337(.A(G2090), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G1966), .B2(new_n711), .ZN(new_n765));
  OR4_X1    g340(.A1(new_n713), .A2(new_n730), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n475), .A2(G128), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT96), .Z(new_n768));
  NOR2_X1   g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT97), .Z(new_n770));
  INV_X1    g345(.A(G116), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n464), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n770), .A2(new_n772), .B1(G140), .B2(new_n462), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G29), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT98), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n715), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT99), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G2067), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G16), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G20), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT23), .Z(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G299), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1956), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n729), .A2(new_n726), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n782), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G4), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n618), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1348), .Z(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n766), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G95), .B(G107), .S(G2105), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G2104), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT91), .ZN(new_n798));
  AOI22_X1  g373(.A1(G119), .A2(new_n475), .B1(new_n462), .B2(G131), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G29), .ZN(new_n801));
  INV_X1    g376(.A(G25), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT90), .B1(new_n802), .B2(G29), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n802), .A2(KEYINPUT90), .A3(G29), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n805), .B(new_n806), .Z(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G24), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n595), .B2(G16), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(G1986), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(G1986), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n807), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n813));
  OR2_X1    g388(.A1(G305), .A2(new_n783), .ZN(new_n814));
  OR2_X1    g389(.A1(G6), .A2(G16), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT92), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n814), .A2(KEYINPUT92), .A3(new_n815), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT32), .B(G1981), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n821), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n818), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G16), .A2(G22), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G166), .B2(G16), .ZN(new_n828));
  INV_X1    g403(.A(G1971), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n574), .A2(new_n581), .A3(KEYINPUT93), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT93), .B1(new_n574), .B2(new_n581), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G16), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G16), .B2(G23), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT33), .B(G1976), .Z(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n830), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n813), .B1(new_n826), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(new_n838), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n841), .A2(KEYINPUT94), .A3(new_n825), .A4(new_n830), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT34), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n812), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(new_n842), .A3(KEYINPUT34), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(KEYINPUT95), .A2(KEYINPUT36), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n795), .B1(new_n850), .B2(new_n851), .ZN(G311));
  INV_X1    g427(.A(new_n851), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n848), .B1(new_n845), .B2(new_n846), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n794), .B1(new_n853), .B2(new_n854), .ZN(G150));
  NAND2_X1  g430(.A1(new_n618), .A2(G559), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  INV_X1    g434(.A(G55), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n512), .A2(new_n859), .B1(new_n860), .B2(new_n514), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n504), .A2(G67), .ZN(new_n862));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n534), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT106), .ZN(new_n865));
  OR3_X1    g440(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n861), .B2(new_n864), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n544), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n543), .B(new_n541), .C1(new_n864), .C2(new_n861), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n858), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT107), .ZN(new_n874));
  AOI21_X1  g449(.A(G860), .B1(new_n871), .B2(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n866), .A2(new_n867), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(G145));
  INV_X1    g455(.A(new_n493), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n487), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n747), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n774), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n740), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n884), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n740), .A2(new_n886), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  MUX2_X1   g466(.A(G106), .B(G118), .S(G2105), .Z(new_n892));
  AOI22_X1  g467(.A1(G130), .A2(new_n475), .B1(new_n892), .B2(G2104), .ZN(new_n893));
  INV_X1    g468(.A(G142), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n648), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n640), .B(new_n895), .Z(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(new_n800), .Z(new_n897));
  AND3_X1   g472(.A1(new_n891), .A2(KEYINPUT110), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n891), .B1(KEYINPUT110), .B2(new_n897), .ZN(new_n899));
  XNOR2_X1  g474(.A(G160), .B(new_n479), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(new_n649), .Z(new_n901));
  NOR3_X1   g476(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(KEYINPUT109), .B(G37), .ZN(new_n903));
  INV_X1    g478(.A(new_n891), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n904), .B2(new_n897), .ZN(new_n905));
  INV_X1    g480(.A(new_n897), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n891), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT40), .Z(G395));
  AOI221_X4 g485(.A(G299), .B1(new_n617), .B2(new_n615), .C1(new_n606), .C2(new_n612), .ZN(new_n911));
  INV_X1    g486(.A(G299), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n606), .A2(new_n612), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(new_n629), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT41), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G299), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(new_n912), .A3(new_n629), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n632), .A2(new_n633), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n618), .A2(KEYINPUT84), .A3(new_n627), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n870), .ZN(new_n924));
  INV_X1    g499(.A(new_n870), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n634), .B2(new_n635), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n911), .A2(new_n914), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n922), .A2(new_n923), .A3(new_n870), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n870), .B1(new_n922), .B2(new_n923), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n833), .A2(new_n595), .ZN(new_n932));
  OAI21_X1  g507(.A(G290), .B1(new_n831), .B2(new_n832), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(G303), .A2(G305), .ZN(new_n935));
  NAND2_X1  g510(.A1(G303), .A2(G305), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n932), .A2(new_n933), .A3(new_n936), .A4(new_n935), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n938), .A2(new_n939), .B1(KEYINPUT111), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n927), .A2(new_n931), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n927), .B2(new_n931), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n940), .A2(KEYINPUT111), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n927), .A2(new_n931), .ZN(new_n947));
  INV_X1    g522(.A(new_n941), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n927), .A2(new_n931), .A3(new_n941), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(G868), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n877), .A2(G868), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT112), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n945), .B1(new_n942), .B2(new_n943), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n949), .A2(new_n944), .A3(new_n950), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n597), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n958), .A2(new_n959), .A3(new_n953), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n955), .A2(new_n960), .ZN(G295));
  NOR2_X1   g536(.A1(new_n958), .A2(new_n953), .ZN(G331));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n963));
  XNOR2_X1  g538(.A(G168), .B(G301), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n870), .ZN(new_n965));
  AOI21_X1  g540(.A(G301), .B1(new_n531), .B2(new_n529), .ZN(new_n966));
  NOR2_X1   g541(.A1(G168), .A2(G171), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n869), .B(new_n868), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(KEYINPUT113), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n925), .B(new_n970), .C1(new_n967), .C2(new_n966), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n965), .A2(new_n968), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n972), .A2(new_n928), .B1(new_n921), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n938), .A2(new_n939), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n903), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n915), .A2(new_n978), .A3(new_n920), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n928), .A2(KEYINPUT114), .A3(new_n918), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n971), .A3(new_n980), .A4(new_n969), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n928), .A2(new_n968), .A3(new_n965), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n963), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n974), .A2(new_n975), .ZN(new_n986));
  INV_X1    g561(.A(G37), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(KEYINPUT43), .A3(new_n987), .A4(new_n976), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n984), .A2(new_n988), .A3(KEYINPUT115), .A4(new_n985), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n977), .B2(new_n983), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n986), .A2(new_n963), .A3(new_n987), .A4(new_n976), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(KEYINPUT44), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n992), .A3(new_n995), .ZN(G397));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n882), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  INV_X1    g574(.A(G40), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n467), .A2(new_n472), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n774), .B(new_n781), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n748), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1002), .ZN(new_n1005));
  INV_X1    g580(.A(G1996), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT117), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1008), .B2(KEYINPUT46), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(KEYINPUT46), .B2(new_n1008), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT47), .Z(new_n1011));
  NOR2_X1   g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT116), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n1005), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT48), .Z(new_n1015));
  OAI21_X1  g590(.A(new_n1003), .B1(new_n1006), .B2(new_n748), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1008), .A2(new_n748), .B1(new_n1005), .B2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n800), .A2(new_n806), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n800), .A2(new_n806), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1005), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1017), .A2(new_n1019), .B1(new_n781), .B2(new_n884), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1015), .A2(new_n1021), .B1(new_n1022), .B2(new_n1002), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1011), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n1001), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT45), .B1(new_n497), .B2(new_n997), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(G2078), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1025), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n998), .A2(new_n999), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(G2078), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1001), .A3(new_n1032), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1028), .A2(KEYINPUT53), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n470), .A2(new_n471), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G2105), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1036), .A2(G40), .A3(new_n466), .A4(new_n463), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n497), .A2(KEYINPUT50), .A3(new_n997), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n493), .B1(new_n482), .B2(new_n486), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(G1384), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1037), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G1961), .ZN(new_n1043));
  OAI21_X1  g618(.A(G171), .B1(new_n1034), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1031), .B1(new_n1045), .B2(G2078), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1043), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1030), .A2(new_n1001), .A3(new_n1048), .A4(new_n1032), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1044), .B(KEYINPUT54), .C1(new_n1050), .C2(G171), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1030), .A2(new_n1001), .A3(new_n1048), .ZN(new_n1054));
  INV_X1    g629(.A(G1966), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1042), .A2(new_n721), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n529), .A2(G8), .A3(new_n531), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1059), .B(KEYINPUT125), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1052), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT125), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1059), .B(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1055), .A2(new_n1054), .B1(new_n1042), .B2(new_n721), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1063), .B(KEYINPUT51), .C1(new_n1064), .C2(new_n1053), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1051), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT93), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G288), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n574), .A2(new_n581), .A3(KEYINPUT93), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(G1976), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT120), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n998), .A2(new_n1037), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1053), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1001), .A2(new_n997), .A3(new_n882), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(KEYINPUT119), .A3(G8), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1070), .A2(new_n1080), .A3(G1976), .A4(new_n1071), .ZN(new_n1081));
  INV_X1    g656(.A(G1976), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(G288), .B2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1073), .A2(new_n1079), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G305), .A2(G1981), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n587), .A2(new_n588), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n513), .A2(G86), .ZN(new_n1088));
  OAI21_X1  g663(.A(G1981), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1086), .A2(KEYINPUT49), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(G305), .B2(G1981), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(new_n1079), .A3(new_n1093), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1084), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(G166), .B2(new_n1053), .ZN(new_n1097));
  NAND3_X1  g672(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n829), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT50), .B1(new_n497), .B2(new_n997), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1040), .A2(new_n1039), .A3(G1384), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n763), .B(new_n1001), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G8), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1105), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1100), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1042), .A2(KEYINPUT118), .A3(new_n763), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1101), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT118), .B1(new_n1042), .B2(new_n763), .ZN(new_n1112));
  OAI211_X1 g687(.A(G8), .B(new_n1099), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1075), .A2(new_n1074), .A3(new_n1053), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT119), .B1(new_n1077), .B2(G8), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1081), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1080), .B1(new_n833), .B2(G1976), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT52), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1095), .A2(new_n1109), .A3(new_n1113), .A4(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1068), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT56), .B(G2072), .Z(new_n1121));
  OR3_X1    g696(.A1(new_n1026), .A2(new_n1027), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1001), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1123));
  INV_X1    g698(.A(G1956), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n566), .B2(new_n570), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1122), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1042), .A2(G1348), .B1(G2067), .B2(new_n1077), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(new_n618), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(KEYINPUT124), .B(new_n1130), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1131), .A2(KEYINPUT60), .A3(new_n916), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1026), .A2(new_n1027), .A3(G1996), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT58), .B(G1341), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1075), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n545), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1144), .B(new_n545), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1138), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1130), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(new_n1133), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1131), .A2(new_n618), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT60), .B1(new_n1132), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1129), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(KEYINPUT61), .A3(new_n1130), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1136), .B(new_n1137), .C1(new_n1150), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1033), .A2(new_n1029), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1046), .A2(new_n1160), .A3(G301), .A4(new_n1047), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT126), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1050), .A2(G171), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1161), .A2(KEYINPUT126), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1159), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1120), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1067), .A2(KEYINPUT62), .ZN(new_n1168));
  AND4_X1   g743(.A1(new_n1113), .A2(new_n1118), .A3(new_n1084), .A4(new_n1094), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1061), .A2(new_n1065), .A3(new_n1170), .A4(new_n1066), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1163), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1169), .A2(new_n1109), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1168), .B1(new_n1173), .B2(KEYINPUT127), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1113), .A2(new_n1118), .A3(new_n1084), .A4(new_n1094), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1109), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1176), .A2(new_n1177), .A3(new_n1163), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1175), .B1(new_n1178), .B2(new_n1171), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1167), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(G288), .A2(G1976), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT121), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1094), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1079), .B1(new_n1183), .B2(new_n1085), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1113), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1095), .A2(new_n1185), .A3(new_n1118), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1064), .A2(new_n1053), .A3(G286), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1169), .A2(new_n1190), .A3(new_n1109), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1190), .A2(KEYINPUT63), .ZN(new_n1194));
  OAI21_X1  g769(.A(G8), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1194), .B1(new_n1100), .B2(new_n1195), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1196), .A2(new_n1169), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1188), .B(new_n1189), .C1(new_n1193), .C2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1191), .A2(new_n1192), .B1(new_n1169), .B2(new_n1196), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT123), .B1(new_n1199), .B2(new_n1187), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1180), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1013), .B1(G1986), .B2(G290), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1017), .B(new_n1020), .C1(new_n1002), .C2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1024), .B1(new_n1201), .B2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g779(.A1(new_n708), .A2(G319), .A3(new_n671), .ZN(new_n1206));
  OR2_X1    g780(.A1(new_n1206), .A2(G227), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n984), .A2(new_n988), .ZN(new_n1208));
  NOR3_X1   g782(.A1(new_n1207), .A2(new_n1208), .A3(new_n909), .ZN(G308));
  OR3_X1    g783(.A1(new_n1207), .A2(new_n1208), .A3(new_n909), .ZN(G225));
endmodule


