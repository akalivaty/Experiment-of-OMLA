

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XOR2_X1 U319 ( .A(n442), .B(n441), .Z(n287) );
  XNOR2_X1 U320 ( .A(n384), .B(G204GAT), .ZN(n385) );
  XNOR2_X1 U321 ( .A(n431), .B(n385), .ZN(n387) );
  XNOR2_X1 U322 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U323 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U324 ( .A(KEYINPUT28), .B(n457), .Z(n528) );
  INV_X1 U325 ( .A(G190GAT), .ZN(n447) );
  NOR2_X1 U326 ( .A1(n525), .A2(n446), .ZN(n558) );
  XNOR2_X1 U327 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U328 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT0), .B(G134GAT), .Z(n289) );
  XNOR2_X1 U330 ( .A(KEYINPUT83), .B(G120GAT), .ZN(n288) );
  XNOR2_X1 U331 ( .A(n289), .B(n288), .ZN(n290) );
  XNOR2_X1 U332 ( .A(G113GAT), .B(n290), .ZN(n316) );
  XOR2_X1 U333 ( .A(KEYINPUT86), .B(G71GAT), .Z(n292) );
  XNOR2_X1 U334 ( .A(G183GAT), .B(G176GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n304) );
  XOR2_X1 U336 ( .A(G15GAT), .B(G127GAT), .Z(n407) );
  XOR2_X1 U337 ( .A(KEYINPUT84), .B(G190GAT), .Z(n294) );
  XNOR2_X1 U338 ( .A(G43GAT), .B(G99GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U340 ( .A(n407), .B(n295), .Z(n297) );
  NAND2_X1 U341 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U343 ( .A(n298), .B(KEYINPUT20), .Z(n302) );
  XOR2_X1 U344 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n300) );
  XNOR2_X1 U345 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n432) );
  XNOR2_X1 U347 ( .A(n432), .B(KEYINPUT85), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n305) );
  XOR2_X1 U350 ( .A(n316), .B(n305), .Z(n489) );
  INV_X1 U351 ( .A(n489), .ZN(n525) );
  XOR2_X1 U352 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n445) );
  XOR2_X1 U353 ( .A(G162GAT), .B(G148GAT), .Z(n307) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(G127GAT), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U356 ( .A(G29GAT), .B(G85GAT), .Z(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n324) );
  XOR2_X1 U358 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n311) );
  XNOR2_X1 U359 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U361 ( .A(G57GAT), .B(KEYINPUT4), .Z(n313) );
  XNOR2_X1 U362 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n322) );
  XOR2_X1 U365 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n320) );
  INV_X1 U366 ( .A(n316), .ZN(n318) );
  XNOR2_X1 U367 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n317), .B(KEYINPUT3), .ZN(n341) );
  XNOR2_X1 U369 ( .A(n318), .B(n341), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n326) );
  NAND2_X1 U373 ( .A1(G225GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n482) );
  INV_X1 U375 ( .A(n482), .ZN(n561) );
  XNOR2_X1 U376 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n327), .B(G162GAT), .ZN(n349) );
  XOR2_X1 U378 ( .A(KEYINPUT23), .B(n349), .Z(n329) );
  NAND2_X1 U379 ( .A1(G228GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n345) );
  XOR2_X1 U381 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n331) );
  XNOR2_X1 U382 ( .A(KEYINPUT87), .B(KEYINPUT22), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(n332), .B(KEYINPUT91), .Z(n334) );
  XOR2_X1 U385 ( .A(G141GAT), .B(G22GAT), .Z(n369) );
  XNOR2_X1 U386 ( .A(n369), .B(KEYINPUT88), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n336) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n335), .B(G148GAT), .ZN(n388) );
  XOR2_X1 U390 ( .A(n336), .B(n388), .Z(n343) );
  XNOR2_X1 U391 ( .A(G211GAT), .B(G218GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n337), .B(KEYINPUT89), .ZN(n338) );
  XOR2_X1 U393 ( .A(n338), .B(KEYINPUT21), .Z(n340) );
  XNOR2_X1 U394 ( .A(G197GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n440) );
  XNOR2_X1 U396 ( .A(n440), .B(n341), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n457) );
  AND2_X1 U399 ( .A1(n561), .A2(n457), .ZN(n443) );
  INV_X1 U400 ( .A(KEYINPUT54), .ZN(n442) );
  XOR2_X1 U401 ( .A(G29GAT), .B(G43GAT), .Z(n347) );
  XNOR2_X1 U402 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n373) );
  XNOR2_X1 U404 ( .A(G99GAT), .B(G85GAT), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n348), .B(KEYINPUT73), .ZN(n391) );
  XNOR2_X1 U406 ( .A(n373), .B(n391), .ZN(n362) );
  XOR2_X1 U407 ( .A(G36GAT), .B(G190GAT), .Z(n433) );
  XOR2_X1 U408 ( .A(n433), .B(n349), .Z(n351) );
  XNOR2_X1 U409 ( .A(G134GAT), .B(G218GAT), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U411 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n353) );
  NAND2_X1 U412 ( .A1(G232GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U414 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U415 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n357) );
  XNOR2_X1 U416 ( .A(G106GAT), .B(G92GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n358), .B(KEYINPUT77), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n548) );
  XOR2_X1 U421 ( .A(KEYINPUT69), .B(G8GAT), .Z(n364) );
  XNOR2_X1 U422 ( .A(G15GAT), .B(G113GAT), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U424 ( .A(KEYINPUT29), .B(KEYINPUT71), .Z(n366) );
  XNOR2_X1 U425 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n380) );
  XOR2_X1 U428 ( .A(G36GAT), .B(G50GAT), .Z(n371) );
  XOR2_X1 U429 ( .A(G1GAT), .B(KEYINPUT70), .Z(n413) );
  XNOR2_X1 U430 ( .A(n369), .B(n413), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U432 ( .A(n372), .B(G197GAT), .Z(n378) );
  XOR2_X1 U433 ( .A(n373), .B(KEYINPUT68), .Z(n375) );
  NAND2_X1 U434 ( .A1(G229GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(n376), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n552) );
  XNOR2_X1 U439 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n398) );
  XOR2_X1 U440 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n382) );
  XNOR2_X1 U441 ( .A(KEYINPUT72), .B(KEYINPUT74), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n397) );
  XNOR2_X1 U443 ( .A(G176GAT), .B(G92GAT), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n383), .B(G64GAT), .ZN(n431) );
  AND2_X1 U445 ( .A1(G230GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U446 ( .A(G71GAT), .B(G57GAT), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n386), .B(KEYINPUT13), .ZN(n403) );
  XOR2_X1 U448 ( .A(n387), .B(n403), .Z(n390) );
  XNOR2_X1 U449 ( .A(G120GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n390), .B(n389), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n391), .B(KEYINPUT75), .ZN(n393) );
  INV_X1 U452 ( .A(KEYINPUT32), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n569) );
  XNOR2_X1 U454 ( .A(n398), .B(n569), .ZN(n554) );
  NAND2_X1 U455 ( .A1(n552), .A2(n554), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n399), .B(KEYINPUT46), .ZN(n420) );
  XOR2_X1 U457 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n405) );
  XOR2_X1 U458 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n401) );
  XNOR2_X1 U459 ( .A(KEYINPUT15), .B(KEYINPUT79), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n419) );
  XNOR2_X1 U463 ( .A(G8GAT), .B(G183GAT), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n406), .B(KEYINPUT78), .ZN(n434) );
  XOR2_X1 U465 ( .A(n407), .B(n434), .Z(n409) );
  NAND2_X1 U466 ( .A1(G231GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n417) );
  XOR2_X1 U468 ( .A(KEYINPUT12), .B(G64GAT), .Z(n411) );
  XNOR2_X1 U469 ( .A(G211GAT), .B(G78GAT), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U471 ( .A(n412), .B(G155GAT), .Z(n415) );
  XNOR2_X1 U472 ( .A(G22GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U474 ( .A(n417), .B(n416), .Z(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n534) );
  NAND2_X1 U476 ( .A1(n420), .A2(n534), .ZN(n421) );
  NOR2_X1 U477 ( .A1(n548), .A2(n421), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n422), .B(KEYINPUT47), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n548), .B(KEYINPUT99), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n423), .B(KEYINPUT36), .ZN(n578) );
  NOR2_X1 U481 ( .A1(n578), .A2(n534), .ZN(n424) );
  XOR2_X1 U482 ( .A(KEYINPUT45), .B(n424), .Z(n425) );
  NOR2_X1 U483 ( .A1(n569), .A2(n425), .ZN(n426) );
  INV_X1 U484 ( .A(n552), .ZN(n564) );
  NAND2_X1 U485 ( .A1(n426), .A2(n564), .ZN(n427) );
  NAND2_X1 U486 ( .A1(n428), .A2(n427), .ZN(n430) );
  XOR2_X1 U487 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n523) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n438) );
  XOR2_X1 U490 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U491 ( .A1(G226GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n513) );
  NOR2_X1 U495 ( .A1(n523), .A2(n513), .ZN(n441) );
  NAND2_X1 U496 ( .A1(n443), .A2(n287), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U498 ( .A1(n558), .A2(n548), .ZN(n450) );
  XOR2_X1 U499 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n448) );
  NOR2_X1 U500 ( .A1(n564), .A2(n569), .ZN(n480) );
  NOR2_X1 U501 ( .A1(n548), .A2(n534), .ZN(n451) );
  XNOR2_X1 U502 ( .A(KEYINPUT16), .B(n451), .ZN(n466) );
  XOR2_X1 U503 ( .A(KEYINPUT27), .B(n513), .Z(n460) );
  NAND2_X1 U504 ( .A1(n460), .A2(n482), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n452), .B(KEYINPUT96), .ZN(n522) );
  NOR2_X1 U506 ( .A1(n522), .A2(n528), .ZN(n453) );
  NAND2_X1 U507 ( .A1(n525), .A2(n453), .ZN(n465) );
  INV_X1 U508 ( .A(n457), .ZN(n455) );
  NOR2_X1 U509 ( .A1(n525), .A2(n513), .ZN(n454) );
  NOR2_X1 U510 ( .A1(n455), .A2(n454), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n456), .B(KEYINPUT25), .ZN(n462) );
  NOR2_X1 U512 ( .A1(n489), .A2(n457), .ZN(n458) );
  XOR2_X1 U513 ( .A(KEYINPUT26), .B(n458), .Z(n459) );
  XNOR2_X1 U514 ( .A(KEYINPUT97), .B(n459), .ZN(n562) );
  NAND2_X1 U515 ( .A1(n562), .A2(n460), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND2_X1 U517 ( .A1(n463), .A2(n561), .ZN(n464) );
  NAND2_X1 U518 ( .A1(n465), .A2(n464), .ZN(n475) );
  AND2_X1 U519 ( .A1(n466), .A2(n475), .ZN(n496) );
  NAND2_X1 U520 ( .A1(n480), .A2(n496), .ZN(n473) );
  NOR2_X1 U521 ( .A1(n561), .A2(n473), .ZN(n468) );
  XNOR2_X1 U522 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U524 ( .A(G1GAT), .B(n469), .Z(G1324GAT) );
  NOR2_X1 U525 ( .A1(n513), .A2(n473), .ZN(n470) );
  XOR2_X1 U526 ( .A(G8GAT), .B(n470), .Z(G1325GAT) );
  NOR2_X1 U527 ( .A1(n525), .A2(n473), .ZN(n472) );
  XNOR2_X1 U528 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(G1326GAT) );
  INV_X1 U530 ( .A(n528), .ZN(n518) );
  NOR2_X1 U531 ( .A1(n518), .A2(n473), .ZN(n474) );
  XOR2_X1 U532 ( .A(G22GAT), .B(n474), .Z(G1327GAT) );
  XOR2_X1 U533 ( .A(G29GAT), .B(KEYINPUT39), .Z(n484) );
  NAND2_X1 U534 ( .A1(n534), .A2(n475), .ZN(n476) );
  XNOR2_X1 U535 ( .A(KEYINPUT100), .B(n476), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n578), .A2(n477), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n509) );
  NAND2_X1 U539 ( .A1(n509), .A2(n480), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT38), .B(n481), .Z(n492) );
  NAND2_X1 U541 ( .A1(n482), .A2(n492), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT102), .B(n485), .ZN(G1328GAT) );
  XOR2_X1 U544 ( .A(G36GAT), .B(KEYINPUT103), .Z(n488) );
  INV_X1 U545 ( .A(n513), .ZN(n486) );
  NAND2_X1 U546 ( .A1(n486), .A2(n492), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1329GAT) );
  NAND2_X1 U548 ( .A1(n492), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  NAND2_X1 U551 ( .A1(n492), .A2(n528), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(KEYINPUT104), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  NAND2_X1 U554 ( .A1(n554), .A2(n564), .ZN(n495) );
  XOR2_X1 U555 ( .A(KEYINPUT106), .B(n495), .Z(n508) );
  NAND2_X1 U556 ( .A1(n496), .A2(n508), .ZN(n505) );
  NOR2_X1 U557 ( .A1(n505), .A2(n561), .ZN(n500) );
  XOR2_X1 U558 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n498) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U562 ( .A1(n513), .A2(n505), .ZN(n501) );
  XOR2_X1 U563 ( .A(KEYINPUT108), .B(n501), .Z(n502) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U565 ( .A1(n525), .A2(n505), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1334GAT) );
  NOR2_X1 U568 ( .A1(n518), .A2(n505), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NAND2_X1 U571 ( .A1(n509), .A2(n508), .ZN(n517) );
  NOR2_X1 U572 ( .A1(n561), .A2(n517), .ZN(n512) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(KEYINPUT111), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NOR2_X1 U576 ( .A1(n513), .A2(n517), .ZN(n514) );
  XOR2_X1 U577 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U578 ( .A1(n525), .A2(n517), .ZN(n515) );
  XOR2_X1 U579 ( .A(KEYINPUT112), .B(n515), .Z(n516) );
  XNOR2_X1 U580 ( .A(G99GAT), .B(n516), .ZN(G1338GAT) );
  NOR2_X1 U581 ( .A1(n518), .A2(n517), .ZN(n520) );
  XNOR2_X1 U582 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NOR2_X1 U585 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U586 ( .A(KEYINPUT114), .B(n524), .Z(n541) );
  NOR2_X1 U587 ( .A1(n525), .A2(n541), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(KEYINPUT115), .ZN(n527) );
  NOR2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n537), .A2(n552), .ZN(n529) );
  XNOR2_X1 U591 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U593 ( .A1(n537), .A2(n554), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT116), .Z(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  INV_X1 U597 ( .A(n534), .ZN(n572) );
  NAND2_X1 U598 ( .A1(n537), .A2(n572), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U602 ( .A1(n537), .A2(n548), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  INV_X1 U604 ( .A(n562), .ZN(n540) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n552), .A2(n549), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n544) );
  NAND2_X1 U609 ( .A1(n549), .A2(n554), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n549), .A2(n572), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT118), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  XOR2_X1 U615 ( .A(G162GAT), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n558), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n556) );
  NAND2_X1 U621 ( .A1(n558), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(n557), .ZN(G1349GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT121), .Z(n560) );
  NAND2_X1 U625 ( .A1(n558), .A2(n572), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  AND2_X1 U627 ( .A1(n561), .A2(n287), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n577) );
  NOR2_X1 U629 ( .A1(n577), .A2(n564), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n566) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U635 ( .A(n577), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n573), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n575) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

