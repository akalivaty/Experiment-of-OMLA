//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  INV_X1    g009(.A(G127gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G113gat), .B(G120gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(KEYINPUT64), .A2(KEYINPUT1), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n213), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G120gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G113gat), .ZN(new_n219));
  INV_X1    g018(.A(G113gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G120gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G127gat), .B(G134gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(new_n215), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT71), .B(KEYINPUT2), .Z(new_n230));
  INV_X1    g029(.A(G141gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G148gat), .ZN(new_n232));
  INV_X1    g031(.A(G148gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G141gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n229), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT73), .ZN(new_n237));
  INV_X1    g036(.A(new_n232), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT72), .B(G148gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(G141gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n242), .A2(new_n228), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n237), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n233), .A2(KEYINPUT72), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT72), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G148gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n247), .A3(G141gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n232), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n242), .A2(new_n228), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(KEYINPUT73), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n236), .B1(new_n244), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n253));
  AOI21_X1  g052(.A(new_n225), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n236), .ZN(new_n255));
  AOI221_X4 g054(.A(new_n237), .B1(new_n242), .B2(new_n228), .C1(new_n248), .C2(new_n232), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT73), .B1(new_n249), .B2(new_n250), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n208), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT5), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n255), .B(new_n225), .C1(new_n256), .C2(new_n257), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n252), .A2(new_n264), .A3(new_n225), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT75), .B1(new_n262), .B2(KEYINPUT4), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT75), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n252), .A2(new_n269), .A3(new_n264), .A4(new_n225), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n270), .A3(new_n263), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n271), .A2(new_n260), .ZN(new_n272));
  INV_X1    g071(.A(new_n225), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(KEYINPUT76), .A3(new_n262), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n208), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n206), .B(new_n267), .C1(new_n272), .C2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n271), .A2(new_n260), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(KEYINPUT5), .A3(new_n278), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n206), .B1(new_n284), .B2(new_n267), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AOI211_X1 g085(.A(new_n281), .B(new_n206), .C1(new_n284), .C2(new_n267), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n290));
  INV_X1    g089(.A(G204gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G197gat), .ZN(new_n292));
  INV_X1    g091(.A(G197gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G204gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(new_n292), .B2(new_n294), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n296), .A2(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G211gat), .B(G218gat), .Z(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n302), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n292), .A2(new_n294), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT68), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n298), .B(KEYINPUT69), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n304), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n290), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n301), .A2(new_n302), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n304), .A3(new_n309), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G226gat), .ZN(new_n316));
  INV_X1    g115(.A(G233gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT27), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT27), .B(G183gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT28), .A3(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT26), .ZN(new_n331));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT26), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(new_n330), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n334), .B1(new_n332), .B2(KEYINPUT24), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342));
  INV_X1    g141(.A(G169gat), .ZN(new_n343));
  INV_X1    g142(.A(G176gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n340), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n319), .A2(new_n323), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT24), .A3(new_n332), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT25), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n340), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n341), .ZN(new_n351));
  AND4_X1   g150(.A1(KEYINPUT25), .A2(new_n350), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n339), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n318), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n346), .A2(KEYINPUT25), .A3(new_n348), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n351), .A3(new_n348), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n356), .A2(new_n359), .B1(new_n329), .B2(new_n338), .ZN(new_n360));
  INV_X1    g159(.A(new_n318), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n315), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n360), .B2(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n353), .A2(new_n318), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n314), .A4(new_n311), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  AND3_X1   g168(.A1(new_n363), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n363), .B2(new_n366), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(new_n366), .ZN(new_n374));
  INV_X1    g173(.A(new_n369), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n289), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n371), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n366), .A3(new_n369), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(KEYINPUT30), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n376), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT80), .B1(new_n288), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n285), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(new_n281), .A3(new_n280), .ZN(new_n386));
  INV_X1    g185(.A(new_n287), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n377), .A2(new_n382), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G227gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n339), .B(new_n225), .C1(new_n349), .C2(new_n352), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n356), .A2(new_n359), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n225), .B1(new_n396), .B2(new_n339), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT32), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G15gat), .B(G43gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(KEYINPUT65), .ZN(new_n403));
  XOR2_X1   g202(.A(G71gat), .B(G99gat), .Z(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n399), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n405), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n398), .B(KEYINPUT32), .C1(new_n400), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n353), .A2(new_n273), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(new_n392), .A3(new_n394), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT34), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT67), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(new_n413), .A3(new_n408), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(KEYINPUT67), .A3(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT77), .B(G22gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n354), .B1(new_n303), .B2(new_n310), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n423), .A2(new_n252), .ZN(new_n424));
  NAND2_X1  g223(.A1(G228gat), .A2(G233gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n426));
  INV_X1    g225(.A(new_n315), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT29), .B1(new_n252), .B2(new_n253), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n424), .B(new_n426), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT31), .B(G50gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n255), .B(new_n253), .C1(new_n256), .C2(new_n257), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n311), .A2(new_n314), .B1(new_n434), .B2(new_n354), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n252), .B1(new_n423), .B2(new_n253), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n425), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n429), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n429), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n422), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n429), .A2(new_n437), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n432), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n429), .A2(new_n437), .A3(new_n433), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n421), .A3(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT35), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n420), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n384), .A2(new_n391), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n417), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n413), .B1(new_n406), .B2(new_n408), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI211_X1 g251(.A(new_n449), .B(new_n413), .C1(new_n406), .C2(new_n408), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n445), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI22_X1  g253(.A1(new_n286), .A2(new_n287), .B1(new_n376), .B2(new_n373), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT35), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n444), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT3), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n434), .B(new_n273), .C1(new_n458), .C2(new_n252), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n266), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n208), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n262), .A2(KEYINPUT76), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n252), .A2(new_n225), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n277), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n207), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(KEYINPUT39), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n207), .B1(new_n266), .B2(new_n459), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n205), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n467), .A2(KEYINPUT40), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT40), .B1(new_n467), .B2(new_n470), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n471), .A2(new_n472), .A3(new_n285), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n457), .B1(new_n383), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT79), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n363), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT37), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n363), .A2(new_n366), .A3(new_n475), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT38), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n375), .B1(new_n374), .B2(KEYINPUT37), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n370), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n477), .B1(new_n363), .B2(new_n366), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT38), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n386), .A2(new_n483), .A3(new_n387), .A4(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n418), .A2(new_n419), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT36), .B1(new_n452), .B2(new_n453), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n474), .A2(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n455), .A2(new_n457), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n448), .A2(new_n456), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G190gat), .B(G218gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT99), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT94), .B(KEYINPUT95), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT41), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501));
  INV_X1    g300(.A(G85gat), .ZN(new_n502));
  INV_X1    g301(.A(G92gat), .ZN(new_n503));
  OAI221_X1 g302(.A(KEYINPUT97), .B1(new_n500), .B2(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G99gat), .ZN(new_n505));
  INV_X1    g304(.A(G106gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT8), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G99gat), .B(G106gat), .Z(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT98), .B(G85gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n503), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT97), .B1(new_n500), .B2(new_n501), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n502), .A2(new_n503), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n512), .B(new_n513), .C1(KEYINPUT97), .C2(new_n501), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n508), .A2(new_n509), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n514), .A2(new_n504), .A3(new_n507), .A4(new_n511), .ZN(new_n516));
  INV_X1    g315(.A(new_n509), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G43gat), .ZN(new_n521));
  INV_X1    g320(.A(G43gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G50gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n523), .A3(KEYINPUT15), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  INV_X1    g325(.A(G29gat), .ZN(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT14), .ZN(new_n529));
  NAND2_X1  g328(.A1(G29gat), .A2(G36gat), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n524), .A2(new_n526), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n522), .A2(KEYINPUT83), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G43gat), .ZN(new_n535));
  AOI21_X1  g334(.A(G50gat), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT84), .B1(new_n520), .B2(G43gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT84), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(new_n522), .A3(G50gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n532), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n531), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(KEYINPUT85), .B(new_n532), .C1(new_n536), .C2(new_n540), .ZN(new_n544));
  INV_X1    g343(.A(new_n524), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n526), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT82), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n529), .A2(new_n526), .A3(KEYINPUT82), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(new_n530), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n499), .B1(new_n519), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n515), .A2(new_n518), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n543), .A2(new_n544), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n545), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n552), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n493), .A2(KEYINPUT99), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n498), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n557), .A2(new_n558), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(new_n553), .A3(new_n519), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n557), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n498), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n561), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n566), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n497), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n564), .B1(new_n560), .B2(new_n561), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n571), .A3(new_n566), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n496), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578));
  INV_X1    g377(.A(G1gat), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(KEYINPUT16), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n578), .A2(new_n579), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT87), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT86), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(G8gat), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n578), .A2(new_n579), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n580), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT86), .B1(new_n588), .B2(KEYINPUT87), .ZN(new_n589));
  INV_X1    g388(.A(G8gat), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(new_n588), .B2(KEYINPUT86), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  OR2_X1    g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT9), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n597));
  INV_X1    g396(.A(G57gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(G64gat), .ZN(new_n599));
  INV_X1    g398(.A(G64gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(G57gat), .B2(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n597), .A2(new_n598), .A3(G64gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n596), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n598), .A2(G64gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n600), .A2(G57gat), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT9), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n593), .A3(new_n594), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT92), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n603), .A2(new_n607), .A3(KEYINPUT92), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n592), .B1(KEYINPUT21), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G127gat), .B(G155gat), .Z(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n612), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G183gat), .B(G211gat), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n624), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n627), .B1(new_n625), .B2(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n620), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n634), .A2(new_n619), .A3(new_n618), .A4(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n516), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n608), .B1(new_n638), .B2(new_n517), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n516), .A2(new_n637), .A3(new_n509), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n610), .A2(new_n515), .A3(new_n611), .A4(new_n518), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n612), .A2(new_n554), .A3(KEYINPUT10), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G230gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n317), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n641), .A2(new_n642), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n648), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n650), .B2(new_n652), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n577), .A2(new_n636), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT101), .ZN(new_n661));
  NAND2_X1  g460(.A1(G229gat), .A2(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n592), .A2(new_n557), .ZN(new_n663));
  INV_X1    g462(.A(new_n553), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n583), .A2(new_n584), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n590), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n667), .B(new_n585), .C1(new_n551), .C2(KEYINPUT17), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT88), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT18), .ZN(new_n671));
  INV_X1    g470(.A(new_n592), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n567), .A3(new_n553), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT88), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n673), .A2(new_n674), .A3(new_n662), .A4(new_n663), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n670), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT89), .B1(new_n592), .B2(new_n557), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT89), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n667), .A2(new_n551), .A3(new_n678), .A4(new_n585), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n663), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n662), .B(KEYINPUT13), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n673), .A2(KEYINPUT18), .A3(new_n662), .A4(new_n663), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(G113gat), .B(G141gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G197gat), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT11), .B(G169gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT12), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT81), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n682), .A2(new_n683), .A3(new_n690), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT90), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n693), .A2(new_n694), .A3(new_n676), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n693), .B2(new_n676), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n577), .A2(new_n636), .A3(new_n698), .A4(new_n659), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n661), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n492), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n288), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n383), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n707), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n704), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n709), .A2(new_n710), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n708), .B1(new_n712), .B2(new_n713), .ZN(G1325gat));
  INV_X1    g513(.A(G15gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n701), .A2(new_n715), .A3(new_n420), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n489), .A2(new_n488), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n716), .B1(new_n720), .B2(new_n715), .ZN(G1326gat));
  NAND2_X1  g520(.A1(new_n701), .A2(new_n457), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  NAND2_X1  g523(.A1(new_n448), .A2(new_n456), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n490), .A2(new_n491), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n577), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n693), .A2(new_n676), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT90), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n693), .A2(new_n676), .A3(new_n694), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n729), .A2(new_n730), .B1(new_n685), .B2(new_n691), .ZN(new_n731));
  INV_X1    g530(.A(new_n659), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n731), .A2(new_n636), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n527), .A3(new_n288), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT45), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n492), .B2(new_n577), .ZN(new_n739));
  INV_X1    g538(.A(new_n577), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n386), .A2(new_n387), .B1(new_n381), .B2(new_n380), .ZN(new_n741));
  INV_X1    g540(.A(new_n453), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n415), .A2(new_n449), .A3(new_n417), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n457), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n446), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n420), .A2(new_n445), .A3(new_n446), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n388), .A2(new_n389), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n747), .B2(KEYINPUT80), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n748), .B2(new_n391), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n474), .A2(new_n486), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n750), .A2(new_n491), .A3(new_n717), .ZN(new_n751));
  OAI211_X1 g550(.A(KEYINPUT44), .B(new_n740), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n739), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n733), .ZN(new_n754));
  OAI21_X1  g553(.A(G29gat), .B1(new_n754), .B2(new_n388), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n755), .ZN(G1328gat));
  NOR3_X1   g555(.A1(new_n734), .A2(G36gat), .A3(new_n389), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g557(.A(G36gat), .B1(new_n754), .B2(new_n389), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1329gat));
  NAND2_X1  g559(.A1(new_n533), .A2(new_n535), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n718), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n420), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n734), .A2(new_n763), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n754), .A2(new_n762), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g565(.A1(new_n734), .A2(G50gat), .A3(new_n445), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n739), .A2(new_n752), .A3(new_n457), .A4(new_n733), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G50gat), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(KEYINPUT104), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT104), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n767), .A2(KEYINPUT103), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT103), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n445), .A2(G50gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n734), .B2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n774), .A2(new_n771), .A3(new_n778), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n772), .A2(new_n773), .B1(new_n779), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g579(.A(new_n636), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n740), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n731), .A3(new_n732), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT105), .B1(new_n492), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n783), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n785), .B(new_n786), .C1(new_n749), .C2(new_n751), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n288), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g588(.A(KEYINPUT106), .B1(new_n784), .B2(new_n787), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(KEYINPUT106), .A3(new_n787), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n383), .B(KEYINPUT107), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n795), .B(new_n796), .Z(G1333gat));
  INV_X1    g596(.A(G71gat), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n784), .A2(new_n787), .A3(new_n798), .A4(new_n420), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n784), .A2(KEYINPUT106), .A3(new_n787), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(new_n790), .A3(new_n717), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n801), .B2(new_n798), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(KEYINPUT50), .B(new_n799), .C1(new_n801), .C2(new_n798), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1334gat));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n457), .A3(new_n792), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g607(.A1(new_n697), .A2(new_n636), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n740), .B(new_n809), .C1(new_n749), .C2(new_n751), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n727), .A2(new_n812), .A3(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(new_n288), .A3(new_n510), .A4(new_n732), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n697), .A2(new_n636), .A3(new_n659), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n753), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n388), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n819), .B2(new_n510), .ZN(G1336gat));
  OAI21_X1  g619(.A(G92gat), .B1(new_n818), .B2(new_n793), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n793), .A2(G92gat), .A3(new_n659), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(new_n815), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n812), .A2(KEYINPUT108), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n727), .B2(new_n809), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n739), .A2(new_n752), .A3(new_n383), .A4(new_n817), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G92gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT109), .B1(new_n832), .B2(KEYINPUT52), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT109), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n835));
  AOI211_X1 g634(.A(new_n834), .B(new_n835), .C1(new_n829), .C2(new_n831), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n824), .B1(new_n833), .B2(new_n836), .ZN(G1337gat));
  OAI21_X1  g636(.A(G99gat), .B1(new_n818), .B2(new_n717), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n420), .A2(new_n505), .A3(new_n732), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n814), .B2(new_n839), .ZN(G1338gat));
  NAND4_X1  g639(.A1(new_n739), .A2(new_n752), .A3(new_n457), .A4(new_n817), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(G106gat), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n827), .A2(new_n828), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n445), .A2(G106gat), .A3(new_n659), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846));
  XOR2_X1   g645(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n847));
  INV_X1    g646(.A(new_n844), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n814), .B2(new_n848), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n845), .A2(new_n846), .B1(new_n849), .B2(new_n842), .ZN(G1339gat));
  NAND3_X1  g649(.A1(new_n644), .A2(new_n648), .A3(new_n645), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n648), .B1(new_n644), .B2(new_n645), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n655), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(KEYINPUT55), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n656), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT55), .B1(new_n852), .B2(new_n855), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n697), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n680), .A2(new_n681), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n662), .B1(new_n673), .B2(new_n663), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n689), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT111), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n732), .C1(new_n696), .C2(new_n695), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n740), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n729), .A2(new_n730), .ZN(new_n868));
  AND4_X1   g667(.A1(new_n868), .A2(new_n859), .A3(new_n740), .A4(new_n865), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n781), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n782), .A2(new_n731), .A3(new_n659), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n457), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n793), .A2(new_n288), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n763), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n875), .A2(new_n220), .A3(new_n731), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n388), .B1(new_n870), .B2(new_n871), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n744), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n697), .A3(new_n793), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n879), .B2(new_n220), .ZN(G1340gat));
  OAI21_X1  g679(.A(G120gat), .B1(new_n875), .B2(new_n659), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n793), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n732), .A2(new_n218), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT112), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n885), .B(new_n886), .ZN(G1341gat));
  NOR3_X1   g686(.A1(new_n875), .A2(new_n211), .A3(new_n781), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n882), .A2(KEYINPUT114), .A3(new_n781), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(G127gat), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT114), .B1(new_n882), .B2(new_n781), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(G1342gat));
  NOR3_X1   g691(.A1(new_n383), .A2(G134gat), .A3(new_n577), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n893), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n894), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT115), .B1(new_n894), .B2(KEYINPUT56), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n872), .A2(new_n740), .A3(new_n874), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT56), .B1(new_n897), .B2(G134gat), .ZN(new_n898));
  INV_X1    g697(.A(new_n894), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n895), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(G1343gat));
  NAND2_X1  g699(.A1(new_n717), .A2(new_n457), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n388), .B(new_n901), .C1(new_n870), .C2(new_n871), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n793), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n231), .B1(new_n903), .B2(new_n731), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n873), .A2(new_n718), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n731), .A2(new_n231), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n870), .A2(new_n871), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n457), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n457), .A2(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n852), .A2(new_n855), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n857), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n697), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n740), .B1(new_n913), .B2(new_n866), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n781), .B1(new_n914), .B2(new_n869), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n909), .B1(new_n915), .B2(new_n871), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n905), .B(new_n906), .C1(new_n908), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n904), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(G1344gat));
  NAND2_X1  g719(.A1(new_n732), .A2(new_n239), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n903), .A2(KEYINPUT117), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT117), .B1(new_n903), .B2(new_n921), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n661), .A2(new_n731), .A3(new_n699), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n445), .B1(new_n928), .B2(new_n915), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n909), .B1(new_n870), .B2(new_n871), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n929), .A2(KEYINPUT57), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n732), .B(new_n905), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n925), .B1(new_n934), .B2(G148gat), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n732), .B(new_n905), .C1(new_n908), .C2(new_n916), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(KEYINPUT59), .A3(new_n239), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n924), .B1(new_n935), .B2(new_n938), .ZN(G1345gat));
  OAI21_X1  g738(.A(new_n905), .B1(new_n908), .B2(new_n916), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n636), .A2(G155gat), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT120), .Z(new_n942));
  OR2_X1    g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G155gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n903), .B2(new_n781), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n943), .A2(new_n945), .ZN(G1346gat));
  OAI21_X1  g745(.A(G162gat), .B1(new_n940), .B2(new_n577), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n383), .A2(G162gat), .A3(new_n577), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n902), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(new_n949), .A3(KEYINPUT121), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1347gat));
  AOI21_X1  g753(.A(new_n288), .B1(new_n870), .B2(new_n871), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n793), .A2(new_n454), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n955), .A2(new_n343), .A3(new_n697), .A4(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n288), .A2(new_n389), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(new_n420), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT123), .Z(new_n962));
  NAND2_X1  g761(.A1(new_n872), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(G169gat), .B1(new_n963), .B2(new_n731), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n959), .A2(KEYINPUT124), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1348gat));
  AND2_X1   g768(.A1(new_n955), .A2(new_n956), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n344), .A3(new_n732), .ZN(new_n971));
  OAI21_X1  g770(.A(G176gat), .B1(new_n963), .B2(new_n659), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  NAND3_X1  g772(.A1(new_n970), .A2(new_n327), .A3(new_n636), .ZN(new_n974));
  OAI21_X1  g773(.A(G183gat), .B1(new_n963), .B2(new_n781), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n970), .A2(new_n323), .A3(new_n740), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n872), .A2(new_n740), .A3(new_n962), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n979), .A2(new_n980), .A3(G190gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n979), .B2(G190gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G1351gat));
  AND2_X1   g782(.A1(new_n960), .A2(new_n717), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n731), .A2(new_n293), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n984), .B(new_n985), .C1(new_n932), .C2(new_n933), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n901), .A2(new_n793), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n955), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n293), .B1(new_n988), .B2(new_n731), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n986), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1352gat));
  OR2_X1    g793(.A1(new_n932), .A2(new_n933), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n995), .A2(new_n732), .A3(new_n984), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G204gat), .ZN(new_n997));
  XNOR2_X1  g796(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n999), .A2(KEYINPUT126), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n988), .A2(G204gat), .A3(new_n659), .ZN(new_n1001));
  MUX2_X1   g800(.A(new_n998), .B(new_n1000), .S(new_n1001), .Z(new_n1002));
  NAND2_X1  g801(.A1(new_n997), .A2(new_n1002), .ZN(G1353gat));
  OR3_X1    g802(.A1(new_n988), .A2(G211gat), .A3(new_n781), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n636), .B(new_n984), .C1(new_n932), .C2(new_n933), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  NAND4_X1  g807(.A1(new_n995), .A2(G218gat), .A3(new_n740), .A4(new_n984), .ZN(new_n1009));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1010), .B1(new_n988), .B2(new_n577), .ZN(new_n1011));
  XNOR2_X1  g810(.A(new_n1011), .B(KEYINPUT127), .ZN(new_n1012));
  AND2_X1   g811(.A1(new_n1009), .A2(new_n1012), .ZN(G1355gat));
endmodule


