

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U324 ( .A(n395), .B(KEYINPUT54), .ZN(n419) );
  XNOR2_X1 U325 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U326 ( .A(n300), .B(G106GAT), .ZN(n301) );
  AND2_X1 U327 ( .A1(n419), .A2(n418), .ZN(n421) );
  XNOR2_X1 U328 ( .A(n373), .B(KEYINPUT48), .ZN(n374) );
  XOR2_X1 U329 ( .A(n311), .B(n310), .Z(n569) );
  INV_X1 U330 ( .A(KEYINPUT33), .ZN(n339) );
  XNOR2_X1 U331 ( .A(n340), .B(n339), .ZN(n341) );
  INV_X1 U332 ( .A(n524), .ZN(n418) );
  XNOR2_X1 U333 ( .A(n342), .B(n341), .ZN(n343) );
  INV_X1 U334 ( .A(KEYINPUT66), .ZN(n420) );
  NOR2_X1 U335 ( .A1(n458), .A2(n555), .ZN(n591) );
  NOR2_X1 U336 ( .A1(n461), .A2(n473), .ZN(n577) );
  XOR2_X1 U337 ( .A(KEYINPUT41), .B(n365), .Z(n544) );
  XNOR2_X1 U338 ( .A(n455), .B(KEYINPUT62), .ZN(n456) );
  XNOR2_X1 U339 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U340 ( .A(n457), .B(n456), .ZN(G1355GAT) );
  XNOR2_X1 U341 ( .A(n465), .B(n464), .ZN(G1349GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT73), .B(G134GAT), .Z(n293) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(G190GAT), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U345 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n295) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U348 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n297) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(KEYINPUT74), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U351 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U352 ( .A(G85GAT), .B(G92GAT), .Z(n330) );
  XOR2_X1 U353 ( .A(KEYINPUT72), .B(G162GAT), .Z(n427) );
  XOR2_X1 U354 ( .A(n330), .B(n427), .Z(n302) );
  NAND2_X1 U355 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n311) );
  XOR2_X1 U358 ( .A(KEYINPUT7), .B(G50GAT), .Z(n308) );
  XNOR2_X1 U359 ( .A(G36GAT), .B(G29GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U361 ( .A(KEYINPUT8), .B(n309), .ZN(n359) );
  INV_X1 U362 ( .A(n359), .ZN(n310) );
  INV_X1 U363 ( .A(n569), .ZN(n578) );
  XOR2_X1 U364 ( .A(KEYINPUT36), .B(n578), .Z(n499) );
  XOR2_X1 U365 ( .A(G57GAT), .B(KEYINPUT13), .Z(n329) );
  XOR2_X1 U366 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n313) );
  XNOR2_X1 U367 ( .A(G71GAT), .B(KEYINPUT14), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(n329), .B(n314), .Z(n317) );
  XNOR2_X1 U370 ( .A(G22GAT), .B(G1GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n315), .B(G8GAT), .ZN(n355) );
  XOR2_X1 U372 ( .A(G155GAT), .B(G78GAT), .Z(n426) );
  XNOR2_X1 U373 ( .A(n355), .B(n426), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U375 ( .A(KEYINPUT76), .B(G64GAT), .Z(n319) );
  NAND2_X1 U376 ( .A1(G231GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U378 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U379 ( .A(G211GAT), .B(G127GAT), .Z(n323) );
  XNOR2_X1 U380 ( .A(G15GAT), .B(G183GAT), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n324), .B(KEYINPUT77), .ZN(n325) );
  XOR2_X1 U383 ( .A(n326), .B(n325), .Z(n590) );
  INV_X1 U384 ( .A(n590), .ZN(n564) );
  NOR2_X1 U385 ( .A1(n499), .A2(n564), .ZN(n328) );
  XNOR2_X1 U386 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n345) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n344) );
  XOR2_X1 U389 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n332) );
  NAND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n334) );
  INV_X1 U392 ( .A(KEYINPUT32), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n338) );
  XNOR2_X1 U394 ( .A(G99GAT), .B(G71GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n335), .B(G120GAT), .ZN(n439) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n336), .B(G148GAT), .ZN(n422) );
  XNOR2_X1 U398 ( .A(n439), .B(n422), .ZN(n337) );
  XNOR2_X1 U399 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U400 ( .A(G176GAT), .B(G64GAT), .Z(n389) );
  XNOR2_X1 U401 ( .A(G78GAT), .B(n389), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n362) );
  INV_X1 U403 ( .A(n362), .ZN(n586) );
  NOR2_X1 U404 ( .A1(n345), .A2(n586), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n346), .B(KEYINPUT112), .ZN(n360) );
  XOR2_X1 U406 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n348) );
  XNOR2_X1 U407 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U409 ( .A(G141GAT), .B(G197GAT), .Z(n350) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U412 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U413 ( .A(G15GAT), .B(G113GAT), .Z(n354) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G43GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n441) );
  XNOR2_X1 U416 ( .A(n441), .B(n355), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n359), .B(n358), .Z(n581) );
  INV_X1 U419 ( .A(n581), .ZN(n557) );
  XOR2_X1 U420 ( .A(KEYINPUT70), .B(n557), .Z(n571) );
  INV_X1 U421 ( .A(n571), .ZN(n466) );
  NAND2_X1 U422 ( .A1(n360), .A2(n466), .ZN(n372) );
  INV_X1 U423 ( .A(KEYINPUT65), .ZN(n361) );
  NAND2_X1 U424 ( .A1(n586), .A2(n361), .ZN(n364) );
  NAND2_X1 U425 ( .A1(n362), .A2(KEYINPUT65), .ZN(n363) );
  NAND2_X1 U426 ( .A1(n364), .A2(n363), .ZN(n365) );
  INV_X1 U427 ( .A(n544), .ZN(n559) );
  NOR2_X1 U428 ( .A1(n557), .A2(n559), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n366), .B(KEYINPUT46), .ZN(n367) );
  XOR2_X1 U430 ( .A(n590), .B(KEYINPUT109), .Z(n574) );
  NOR2_X1 U431 ( .A1(n367), .A2(n574), .ZN(n368) );
  NAND2_X1 U432 ( .A1(n368), .A2(n569), .ZN(n370) );
  XOR2_X1 U433 ( .A(KEYINPUT110), .B(KEYINPUT47), .Z(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n371) );
  NAND2_X1 U435 ( .A1(n372), .A2(n371), .ZN(n375) );
  XOR2_X1 U436 ( .A(KEYINPUT64), .B(KEYINPUT113), .Z(n373) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n537) );
  XNOR2_X1 U438 ( .A(KEYINPUT83), .B(KEYINPUT18), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n376), .B(KEYINPUT19), .ZN(n377) );
  XOR2_X1 U440 ( .A(n377), .B(KEYINPUT17), .Z(n379) );
  XNOR2_X1 U441 ( .A(G183GAT), .B(G190GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n440) );
  XOR2_X1 U443 ( .A(KEYINPUT21), .B(G218GAT), .Z(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT88), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U446 ( .A(G197GAT), .B(n382), .Z(n437) );
  XOR2_X1 U447 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n384) );
  XNOR2_X1 U448 ( .A(G169GAT), .B(G8GAT), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n437), .B(n385), .ZN(n393) );
  XOR2_X1 U451 ( .A(KEYINPUT74), .B(G92GAT), .Z(n387) );
  XNOR2_X1 U452 ( .A(G36GAT), .B(G204GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U454 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(n440), .B(n394), .Z(n527) );
  AND2_X1 U459 ( .A1(n537), .A2(n527), .ZN(n395) );
  XOR2_X1 U460 ( .A(G85GAT), .B(G155GAT), .Z(n397) );
  XNOR2_X1 U461 ( .A(G113GAT), .B(G148GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n399) );
  XOR2_X1 U463 ( .A(G29GAT), .B(G162GAT), .Z(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n415) );
  XOR2_X1 U465 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n401) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U468 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n403) );
  XNOR2_X1 U469 ( .A(G120GAT), .B(KEYINPUT1), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U471 ( .A(n405), .B(n404), .ZN(n413) );
  XOR2_X1 U472 ( .A(G57GAT), .B(KEYINPUT89), .Z(n411) );
  XOR2_X1 U473 ( .A(KEYINPUT80), .B(G134GAT), .Z(n407) );
  XNOR2_X1 U474 ( .A(KEYINPUT79), .B(G127GAT), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U476 ( .A(KEYINPUT0), .B(n408), .Z(n438) );
  XNOR2_X1 U477 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n409) );
  XNOR2_X1 U478 ( .A(n409), .B(KEYINPUT3), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n438), .B(n423), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n417) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n524) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n458) );
  XOR2_X1 U486 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n453) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n425) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U491 ( .A(KEYINPUT87), .B(n426), .Z(n429) );
  XNOR2_X1 U492 ( .A(G50GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U494 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n475) );
  XOR2_X1 U499 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n451) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XOR2_X1 U503 ( .A(KEYINPUT82), .B(KEYINPUT85), .Z(n445) );
  XNOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n447) );
  XOR2_X1 U506 ( .A(KEYINPUT84), .B(KEYINPUT81), .Z(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n539) );
  INV_X1 U510 ( .A(n539), .ZN(n473) );
  NAND2_X1 U511 ( .A1(n475), .A2(n473), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n555) );
  INV_X1 U513 ( .A(n591), .ZN(n454) );
  NOR2_X1 U514 ( .A1(n454), .A2(n499), .ZN(n457) );
  INV_X1 U515 ( .A(G218GAT), .ZN(n455) );
  NOR2_X1 U516 ( .A1(n458), .A2(n475), .ZN(n460) );
  XNOR2_X1 U517 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U519 ( .A1(n577), .A2(n544), .ZN(n465) );
  XOR2_X1 U520 ( .A(G176GAT), .B(KEYINPUT56), .Z(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n462) );
  XOR2_X1 U522 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n487) );
  OR2_X1 U523 ( .A1(n466), .A2(n586), .ZN(n501) );
  XOR2_X1 U524 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n468) );
  NAND2_X1 U525 ( .A1(n590), .A2(n569), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n468), .B(n467), .ZN(n485) );
  XOR2_X1 U527 ( .A(KEYINPUT86), .B(n539), .Z(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT28), .B(n475), .ZN(n532) );
  XOR2_X1 U529 ( .A(KEYINPUT27), .B(n527), .Z(n478) );
  INV_X1 U530 ( .A(n478), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n524), .A2(n469), .ZN(n554) );
  NOR2_X1 U532 ( .A1(n532), .A2(n554), .ZN(n538) );
  NAND2_X1 U533 ( .A1(n470), .A2(n538), .ZN(n471) );
  XOR2_X1 U534 ( .A(KEYINPUT94), .B(n471), .Z(n483) );
  INV_X1 U535 ( .A(n527), .ZN(n472) );
  NOR2_X1 U536 ( .A1(n473), .A2(n472), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U538 ( .A(n476), .B(KEYINPUT96), .Z(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT25), .B(n477), .ZN(n480) );
  NOR2_X1 U540 ( .A1(n555), .A2(n478), .ZN(n479) );
  NOR2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n481) );
  NOR2_X1 U542 ( .A1(n524), .A2(n481), .ZN(n482) );
  NOR2_X1 U543 ( .A1(n483), .A2(n482), .ZN(n496) );
  INV_X1 U544 ( .A(n496), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n485), .A2(n484), .ZN(n511) );
  NOR2_X1 U546 ( .A1(n501), .A2(n511), .ZN(n494) );
  NAND2_X1 U547 ( .A1(n494), .A2(n524), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n490) );
  NAND2_X1 U551 ( .A1(n494), .A2(n527), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .Z(n493) );
  NAND2_X1 U555 ( .A1(n494), .A2(n539), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  NAND2_X1 U557 ( .A1(n494), .A2(n532), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n495), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n504) );
  NOR2_X1 U560 ( .A1(n496), .A2(n590), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(KEYINPUT101), .ZN(n498) );
  NOR2_X1 U562 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT37), .B(n500), .ZN(n523) );
  NOR2_X1 U564 ( .A1(n501), .A2(n523), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT38), .ZN(n509) );
  NAND2_X1 U566 ( .A1(n524), .A2(n509), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G29GAT), .B(n505), .ZN(G1328GAT) );
  NAND2_X1 U569 ( .A1(n527), .A2(n509), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n506), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n539), .A2(n509), .ZN(n507) );
  XNOR2_X1 U572 ( .A(KEYINPUT40), .B(n507), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U574 ( .A1(n509), .A2(n532), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT42), .B(KEYINPUT102), .Z(n513) );
  NAND2_X1 U577 ( .A1(n557), .A2(n544), .ZN(n522) );
  NOR2_X1 U578 ( .A1(n522), .A2(n511), .ZN(n518) );
  NAND2_X1 U579 ( .A1(n518), .A2(n524), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n514), .Z(G1332GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n527), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U584 ( .A(G71GAT), .B(KEYINPUT103), .Z(n517) );
  NAND2_X1 U585 ( .A1(n518), .A2(n539), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n520) );
  NAND2_X1 U588 ( .A1(n518), .A2(n532), .ZN(n519) );
  XNOR2_X1 U589 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(n521), .ZN(G1335GAT) );
  XOR2_X1 U591 ( .A(G85GAT), .B(KEYINPUT105), .Z(n526) );
  NOR2_X1 U592 ( .A1(n523), .A2(n522), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n533), .A2(n524), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n530) );
  NAND2_X1 U598 ( .A1(n533), .A2(n539), .ZN(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U600 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n535) );
  NAND2_X1 U602 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U604 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  INV_X1 U605 ( .A(n537), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n550), .A2(n571), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(KEYINPUT114), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U612 ( .A1(n550), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n548) );
  NAND2_X1 U615 ( .A1(n550), .A2(n574), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n552) );
  NAND2_X1 U619 ( .A1(n550), .A2(n578), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n556), .A2(n537), .ZN(n568) );
  NOR2_X1 U624 ( .A1(n557), .A2(n568), .ZN(n558) );
  XOR2_X1 U625 ( .A(G141GAT), .B(n558), .Z(G1344GAT) );
  NOR2_X1 U626 ( .A1(n568), .A2(n559), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n561) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U631 ( .A1(n564), .A2(n568), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G155GAT), .B(n567), .ZN(G1346GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(G162GAT), .B(n570), .Z(G1347GAT) );
  XOR2_X1 U637 ( .A(G169GAT), .B(KEYINPUT121), .Z(n573) );
  NAND2_X1 U638 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1348GAT) );
  XOR2_X1 U640 ( .A(G183GAT), .B(KEYINPUT123), .Z(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1350GAT) );
  XNOR2_X1 U643 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1351GAT) );
  XNOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT124), .ZN(n585) );
  XOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT59), .Z(n583) );
  NAND2_X1 U648 ( .A1(n591), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n588) );
  NAND2_X1 U652 ( .A1(n591), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(n589) );
  XOR2_X1 U654 ( .A(G204GAT), .B(n589), .Z(G1353GAT) );
  XOR2_X1 U655 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n593) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G211GAT), .B(n594), .ZN(G1354GAT) );
endmodule

