//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n208), .A2(new_n209), .B1(G169gat), .B2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(KEYINPUT24), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n207), .A2(new_n210), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n207), .A2(new_n210), .A3(new_n215), .A4(KEYINPUT25), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221));
  INV_X1    g020(.A(G127gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G134gat), .ZN(new_n223));
  INV_X1    g022(.A(G134gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G127gat), .ZN(new_n225));
  OAI22_X1  g024(.A1(new_n221), .A2(KEYINPUT1), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G120gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G113gat), .ZN(new_n228));
  INV_X1    g027(.A(G113gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G120gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT27), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G183gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n212), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(new_n239), .A3(new_n212), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT28), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n203), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n203), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n242), .A2(new_n245), .A3(new_n214), .A4(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n220), .A2(new_n236), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n236), .B1(new_n220), .B2(new_n250), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G227gat), .A2(G233gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(KEYINPUT64), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT34), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT34), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(new_n260), .A3(new_n257), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n202), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G15gat), .B(G43gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G71gat), .B(G99gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n256), .B1(new_n252), .B2(new_n253), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT33), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n220), .A2(new_n250), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n235), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n257), .B1(new_n271), .B2(new_n251), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT32), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT66), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n267), .A2(new_n275), .A3(KEYINPUT32), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n269), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n269), .A2(new_n274), .A3(new_n276), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n266), .A2(new_n268), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n272), .A2(new_n273), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n263), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  AOI211_X1 g084(.A(new_n283), .B(new_n262), .C1(new_n278), .C2(new_n280), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT36), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT36), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n281), .A2(new_n284), .B1(new_n259), .B2(new_n261), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n259), .A2(new_n261), .ZN(new_n291));
  AOI211_X1 g090(.A(new_n283), .B(new_n291), .C1(new_n278), .C2(new_n280), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n288), .A2(new_n293), .A3(KEYINPUT69), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n287), .A2(new_n295), .A3(KEYINPUT36), .ZN(new_n296));
  INV_X1    g095(.A(G141gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G148gat), .ZN(new_n298));
  INV_X1    g097(.A(G148gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT2), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n302), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n301), .A2(new_n303), .B1(new_n307), .B2(KEYINPUT74), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n307), .A2(KEYINPUT74), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n299), .ZN(new_n312));
  NAND2_X1  g111(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(G141gat), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n298), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n302), .B1(new_n306), .B2(KEYINPUT2), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n315), .A2(KEYINPUT76), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT76), .B1(new_n315), .B2(new_n316), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT80), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT80), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n322), .B(new_n310), .C1(new_n317), .C2(new_n318), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n320), .A2(new_n321), .A3(new_n236), .A4(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT82), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(KEYINPUT82), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327));
  INV_X1    g126(.A(new_n298), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n331), .B2(G141gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n316), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n327), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n315), .A2(KEYINPUT76), .A3(new_n316), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n334), .A2(new_n335), .B1(new_n309), .B2(new_n308), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n236), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n325), .A2(new_n326), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342));
  XOR2_X1   g141(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n343));
  OAI211_X1 g142(.A(new_n310), .B(new_n343), .C1(new_n317), .C2(new_n318), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n226), .A2(new_n234), .A3(KEYINPUT77), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT77), .B1(new_n226), .B2(new_n234), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n335), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n310), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n342), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n353), .A2(KEYINPUT79), .A3(new_n347), .A4(new_n344), .ZN(new_n354));
  AOI211_X1 g153(.A(KEYINPUT5), .B(new_n341), .C1(new_n352), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n354), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n321), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n320), .A2(KEYINPUT4), .A3(new_n236), .A4(new_n323), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n356), .A2(new_n340), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  INV_X1    g159(.A(new_n347), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n337), .B1(new_n361), .B2(new_n336), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n362), .B2(new_n341), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n339), .A2(new_n355), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G1gat), .B(G29gat), .Z(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G57gat), .B(G85gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT6), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n339), .A2(new_n355), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n363), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n376), .B2(new_n369), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n372), .B1(new_n377), .B2(new_n371), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n270), .A2(KEYINPUT71), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT71), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n220), .A2(new_n382), .A3(new_n250), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n270), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT72), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n380), .ZN(new_n388));
  XNOR2_X1  g187(.A(G197gat), .B(G204gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT22), .ZN(new_n390));
  INV_X1    g189(.A(G211gat), .ZN(new_n391));
  INV_X1    g190(.A(G218gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(G211gat), .B(G218gat), .Z(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT29), .B1(new_n220), .B2(new_n250), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT72), .B1(new_n397), .B2(new_n381), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n384), .A2(new_n388), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n381), .A2(KEYINPUT29), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n379), .A2(new_n383), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n396), .B(KEYINPUT70), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n220), .A2(new_n381), .A3(new_n250), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  NAND3_X1  g207(.A1(new_n399), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n399), .B2(new_n405), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT73), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n409), .A2(new_n414), .A3(new_n410), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n409), .B2(new_n410), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n378), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  INV_X1    g219(.A(G228gat), .ZN(new_n421));
  INV_X1    g220(.A(G233gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n343), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n396), .B2(new_n385), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n320), .B2(new_n323), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n396), .B1(new_n344), .B2(new_n385), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT83), .B(new_n424), .C1(new_n427), .C2(new_n428), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n344), .A2(new_n385), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n402), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n396), .A2(new_n385), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n353), .B(new_n423), .C1(new_n336), .C2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n420), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  AOI211_X1 g240(.A(G22gat), .B(new_n439), .C1(new_n431), .C2(new_n432), .ZN(new_n442));
  OAI21_X1  g241(.A(G78gat), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n426), .ZN(new_n444));
  INV_X1    g243(.A(new_n323), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n322), .B1(new_n350), .B2(new_n310), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n396), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n434), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT83), .B1(new_n450), .B2(new_n424), .ZN(new_n451));
  INV_X1    g250(.A(new_n432), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n440), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G22gat), .ZN(new_n454));
  INV_X1    g253(.A(G78gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n433), .A2(new_n420), .A3(new_n440), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G50gat), .ZN(new_n458));
  INV_X1    g257(.A(G106gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n443), .B2(new_n457), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n294), .B(new_n296), .C1(new_n419), .C2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n324), .A2(KEYINPUT82), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n338), .B1(new_n324), .B2(KEYINPUT82), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n356), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n341), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n370), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT39), .B1(new_n362), .B2(new_n341), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n469), .B2(new_n341), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n466), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT40), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n469), .A2(new_n341), .ZN(new_n477));
  INV_X1    g276(.A(new_n473), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT84), .A3(new_n370), .A4(new_n471), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n475), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n475), .A2(new_n480), .A3(KEYINPUT85), .A4(new_n476), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n479), .A2(KEYINPUT40), .A3(new_n370), .A4(new_n471), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT86), .B1(new_n364), .B2(new_n370), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n376), .A2(new_n487), .A3(new_n369), .ZN(new_n488));
  AND4_X1   g287(.A1(new_n485), .A2(new_n417), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n483), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT6), .B1(new_n364), .B2(new_n370), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n491), .A3(new_n488), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n399), .A2(new_n405), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n408), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n399), .A2(new_n405), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n493), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n384), .A2(new_n388), .A3(new_n398), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n401), .A2(new_n404), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n500), .A2(new_n448), .B1(new_n501), .B2(new_n402), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n493), .B1(new_n502), .B2(new_n495), .ZN(new_n503));
  INV_X1    g302(.A(new_n408), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n497), .B2(KEYINPUT37), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n409), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n507), .A3(new_n372), .ZN(new_n508));
  INV_X1    g307(.A(new_n460), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n441), .A2(new_n442), .A3(G78gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n455), .B1(new_n454), .B2(new_n456), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n508), .A2(new_n461), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT87), .B1(new_n490), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n508), .A2(new_n461), .A3(new_n512), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT87), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n483), .A2(new_n484), .A3(new_n489), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n465), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  AOI211_X1 g318(.A(KEYINPUT35), .B(new_n417), .C1(new_n492), .C2(new_n372), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n290), .A2(new_n292), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n520), .A2(new_n464), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n512), .A2(new_n287), .A3(new_n461), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n512), .A2(new_n287), .A3(KEYINPUT88), .A4(new_n461), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n419), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n522), .B1(KEYINPUT35), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT89), .B1(new_n519), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n465), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n534));
  INV_X1    g333(.A(new_n522), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n529), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G8gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(G1gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(G1gat), .B2(new_n541), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT14), .B(G29gat), .ZN(new_n550));
  INV_X1    g349(.A(G36gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G29gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G43gat), .B(G50gat), .Z(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n552), .A2(new_n556), .A3(new_n554), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n549), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n549), .B2(new_n558), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT92), .B1(new_n548), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(KEYINPUT17), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n547), .ZN(new_n564));
  MUX2_X1   g363(.A(KEYINPUT92), .B(new_n562), .S(new_n564), .Z(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n569), .A2(KEYINPUT18), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G197gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT11), .B(G169gat), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT12), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n561), .B(new_n547), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(new_n566), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n569), .A2(KEYINPUT18), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n570), .A2(new_n576), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT95), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n582), .A2(new_n581), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(KEYINPUT95), .A3(new_n576), .A4(new_n570), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n570), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n575), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n539), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n378), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n563), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT41), .ZN(new_n605));
  INV_X1    g404(.A(G232gat), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n605), .A2(new_n606), .A3(new_n422), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n561), .B2(new_n602), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(KEYINPUT98), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(KEYINPUT98), .B2(new_n612), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n605), .B1(new_n606), .B2(new_n422), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT97), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n611), .A2(new_n617), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n612), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(KEYINPUT96), .A2(G57gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G64gat), .ZN(new_n624));
  INV_X1    g423(.A(G71gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n455), .ZN(new_n626));
  NOR2_X1   g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n627), .A2(KEYINPUT9), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n624), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  AND2_X1   g429(.A1(G57gat), .A2(G64gat), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G127gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n547), .B1(new_n635), .B2(new_n634), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G155gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n641), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n622), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n595), .A2(new_n601), .A3(new_n599), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n629), .B(new_n633), .C1(new_n649), .C2(KEYINPUT99), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n602), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n603), .A2(new_n654), .A3(new_n634), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n651), .A2(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n653), .B1(new_n658), .B2(new_n652), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT101), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n659), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n648), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT102), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n592), .A2(new_n593), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g470(.A1(new_n592), .A2(new_n669), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n540), .B1(new_n673), .B2(new_n417), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT16), .B(G8gat), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n672), .A2(new_n418), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(KEYINPUT42), .B2(new_n676), .ZN(G1325gat));
  NAND2_X1  g477(.A1(new_n294), .A2(new_n296), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n672), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n521), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n672), .B2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n672), .A2(new_n464), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT103), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NOR3_X1   g487(.A1(new_n622), .A2(new_n647), .A3(new_n666), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n539), .A2(new_n591), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n593), .A2(new_n553), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n690), .A2(KEYINPUT104), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT104), .B1(new_n690), .B2(new_n691), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(KEYINPUT45), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n666), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n591), .A2(new_n646), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n622), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n529), .A2(new_n538), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n514), .A2(new_n518), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT105), .B1(new_n700), .B2(new_n530), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702));
  AOI211_X1 g501(.A(new_n702), .B(new_n465), .C1(new_n514), .C2(new_n518), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n536), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n622), .B(KEYINPUT106), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(KEYINPUT44), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n696), .B1(new_n699), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(new_n593), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n694), .B1(new_n709), .B2(new_n553), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT45), .B1(new_n692), .B2(new_n693), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT107), .ZN(G1328gat));
  INV_X1    g512(.A(new_n690), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n551), .A3(new_n417), .ZN(new_n715));
  AND2_X1   g514(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n708), .A2(new_n417), .ZN(new_n719));
  OAI221_X1 g518(.A(new_n718), .B1(new_n551), .B2(new_n719), .C1(new_n716), .C2(new_n715), .ZN(G1329gat));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n708), .B2(new_n679), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n723), .A2(KEYINPUT109), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(KEYINPUT47), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n690), .A2(G43gat), .A3(new_n682), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT110), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n722), .A2(KEYINPUT110), .A3(new_n726), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n727), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(KEYINPUT47), .B2(new_n724), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1330gat));
  INV_X1    g531(.A(G50gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n464), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n708), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n690), .A2(G50gat), .A3(new_n464), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT111), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n533), .A2(new_n702), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n519), .A2(KEYINPUT105), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n528), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR4_X1   g540(.A1(new_n741), .A2(new_n591), .A3(new_n648), .A4(new_n695), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n593), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g543(.A(new_n418), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT112), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1333gat));
  AOI21_X1  g548(.A(new_n625), .B1(new_n742), .B2(new_n679), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n682), .A2(G71gat), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n742), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n742), .A2(new_n734), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  AOI22_X1  g554(.A1(new_n585), .A2(new_n587), .B1(new_n575), .B2(new_n589), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n646), .A3(new_n666), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n756), .A2(KEYINPUT113), .A3(new_n646), .A4(new_n666), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n699), .B2(new_n707), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G85gat), .B1(new_n763), .B2(new_n378), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n591), .A2(new_n647), .A3(new_n622), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n741), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n704), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n666), .A2(new_n597), .A3(new_n593), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n764), .B1(new_n771), .B2(new_n772), .ZN(G1336gat));
  NOR3_X1   g572(.A1(new_n695), .A2(G92gat), .A3(new_n418), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n768), .B2(new_n769), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n699), .A2(new_n707), .ZN(new_n777));
  INV_X1    g576(.A(new_n761), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n417), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n776), .B1(new_n779), .B2(G92gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n770), .A2(new_n774), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n418), .B(new_n761), .C1(new_n699), .C2(new_n707), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n598), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT114), .B1(new_n786), .B2(KEYINPUT52), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n780), .B2(new_n782), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n598), .B1(new_n762), .B2(new_n417), .ZN(new_n790));
  NOR4_X1   g589(.A1(new_n790), .A2(KEYINPUT115), .A3(KEYINPUT52), .A4(new_n776), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n783), .A2(new_n787), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT115), .B1(new_n786), .B2(KEYINPUT52), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n788), .A3(new_n782), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n797), .B(KEYINPUT116), .C1(new_n787), .C2(new_n783), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(new_n798), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n763), .B2(new_n680), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n695), .A2(G99gat), .A3(new_n682), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n771), .B2(new_n801), .ZN(G1338gat));
  AOI21_X1  g601(.A(new_n459), .B1(new_n762), .B2(new_n734), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n695), .A2(new_n464), .A3(G106gat), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n770), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n803), .B2(KEYINPUT117), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n805), .B(new_n807), .Z(G1339gat));
  NAND2_X1  g607(.A1(new_n756), .A2(new_n667), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n658), .A2(new_n652), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n810), .A2(KEYINPUT54), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n658), .A2(new_n652), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n814), .A2(KEYINPUT118), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(KEYINPUT118), .ZN(new_n816));
  AOI211_X1 g615(.A(new_n662), .B(new_n812), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n664), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(KEYINPUT55), .B2(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n577), .A2(new_n580), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n822), .B1(new_n565), .B2(new_n566), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n574), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n588), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n821), .A2(new_n826), .A3(new_n705), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n821), .A2(new_n756), .B1(new_n826), .B2(new_n695), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n705), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n809), .B1(new_n829), .B2(new_n647), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n830), .A2(new_n464), .A3(new_n521), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n418), .A3(new_n593), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n832), .A2(new_n229), .A3(new_n756), .ZN(new_n833));
  INV_X1    g632(.A(new_n830), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n378), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n525), .A2(new_n526), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n835), .A2(new_n418), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n591), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n838), .B2(new_n229), .ZN(G1340gat));
  NOR3_X1   g638(.A1(new_n832), .A2(new_n227), .A3(new_n695), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n666), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n227), .ZN(G1341gat));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n222), .A3(new_n647), .ZN(new_n843));
  OAI21_X1  g642(.A(G127gat), .B1(new_n832), .B2(new_n646), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1342gat));
  NOR2_X1   g644(.A1(new_n622), .A2(new_n417), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n835), .A2(new_n224), .A3(new_n836), .A4(new_n846), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n832), .B2(new_n622), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(G1343gat));
  XNOR2_X1  g650(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n817), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n756), .A2(new_n819), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n826), .A2(new_n695), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n622), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n827), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n647), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n809), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n734), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n830), .A2(new_n862), .A3(new_n734), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n593), .A2(new_n418), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n679), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n861), .A2(new_n863), .A3(new_n591), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n865), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n860), .B2(KEYINPUT57), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(KEYINPUT121), .A3(new_n591), .A4(new_n863), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n868), .A2(G141gat), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n679), .A2(new_n464), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n830), .A2(new_n593), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n756), .A2(G141gat), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n830), .A2(KEYINPUT120), .A3(new_n593), .A4(new_n873), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n876), .A2(new_n418), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR4_X1   g680(.A1(new_n874), .A2(G141gat), .A3(new_n417), .A4(new_n756), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n882), .B1(G141gat), .B2(new_n866), .ZN(new_n883));
  OAI22_X1  g682(.A1(new_n872), .A2(new_n881), .B1(new_n880), .B2(new_n883), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n870), .A2(new_n863), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(KEYINPUT59), .A3(new_n695), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n830), .A2(new_n734), .ZN(new_n887));
  OR3_X1    g686(.A1(new_n821), .A2(new_n826), .A3(new_n622), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n856), .A2(new_n888), .ZN(new_n889));
  OAI22_X1  g688(.A1(new_n889), .A2(new_n647), .B1(new_n591), .B2(new_n668), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n464), .A2(KEYINPUT57), .ZN(new_n891));
  AOI22_X1  g690(.A1(KEYINPUT57), .A2(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n666), .A3(new_n865), .ZN(new_n893));
  AND2_X1   g692(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n876), .A2(new_n418), .A3(new_n666), .A4(new_n878), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT59), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n331), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n898), .ZN(G1345gat));
  OAI21_X1  g698(.A(G155gat), .B1(new_n885), .B2(new_n646), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n876), .A2(new_n878), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n418), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n647), .A2(new_n304), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(G1346gat));
  NAND3_X1  g703(.A1(new_n901), .A2(new_n305), .A3(new_n846), .ZN(new_n905));
  OAI21_X1  g704(.A(G162gat), .B1(new_n885), .B2(new_n705), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n593), .A2(new_n418), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n831), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(G169gat), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n909), .A2(new_n910), .A3(new_n756), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n834), .A2(new_n593), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n836), .A2(new_n417), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n591), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n910), .B2(new_n914), .ZN(G1348gat));
  INV_X1    g714(.A(G176gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n909), .A2(new_n916), .A3(new_n695), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n912), .A2(new_n913), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n918), .B2(new_n695), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT122), .B(new_n916), .C1(new_n918), .C2(new_n695), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(G1349gat));
  OAI21_X1  g722(.A(G183gat), .B1(new_n909), .B2(new_n646), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n912), .A2(new_n240), .A3(new_n647), .A4(new_n913), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n909), .B2(new_n622), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n705), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n912), .A2(new_n212), .A3(new_n935), .A4(new_n913), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n932), .A2(new_n933), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n938), .A3(new_n939), .ZN(G1351gat));
  NOR3_X1   g739(.A1(new_n679), .A2(new_n418), .A3(new_n464), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n912), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT125), .B(G197gat), .Z(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n591), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n680), .A2(new_n908), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT126), .Z(new_n947));
  NAND2_X1  g746(.A1(new_n892), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n756), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n949), .B2(new_n944), .ZN(G1352gat));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n890), .A2(new_n891), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n666), .A4(new_n947), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(new_n955), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n695), .A2(G204gat), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT62), .B1(new_n942), .B2(new_n959), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n942), .A2(KEYINPUT62), .A3(new_n959), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n960), .A3(new_n961), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n943), .A2(new_n391), .A3(new_n647), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n892), .A2(new_n647), .A3(new_n947), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  OAI21_X1  g766(.A(G218gat), .B1(new_n948), .B2(new_n622), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n943), .A2(new_n392), .A3(new_n935), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1355gat));
endmodule


