//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984;
  AND2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT76), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  INV_X1    g004(.A(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n208));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n204), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OR3_X1    g011(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n213), .A2(new_n214), .B1(G155gat), .B2(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n211), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n217), .B2(new_n218), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n202), .A2(new_n203), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n216), .A2(new_n225), .A3(new_n222), .ZN(new_n226));
  AND2_X1   g025(.A1(G113gat), .A2(G120gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G113gat), .A2(G120gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT66), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G113gat), .ZN(new_n230));
  OR3_X1    g029(.A1(new_n230), .A2(KEYINPUT66), .A3(G120gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n229), .A2(new_n231), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(KEYINPUT65), .A2(G127gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT65), .A2(G127gat), .ZN(new_n236));
  OAI21_X1  g035(.A(G134gat), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G120gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g039(.A1(G113gat), .A2(G120gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G127gat), .ZN(new_n243));
  INV_X1    g042(.A(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n237), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n234), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n224), .A2(new_n226), .A3(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n234), .A2(new_n246), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n212), .A2(new_n215), .B1(new_n221), .B2(new_n220), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n253));
  AOI21_X1  g052(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n248), .B(new_n254), .C1(new_n255), .C2(new_n252), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n223), .A2(new_n247), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n252), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n259), .B2(new_n249), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n252), .A2(new_n253), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n252), .A2(new_n255), .ZN(new_n263));
  INV_X1    g062(.A(new_n257), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(new_n249), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n262), .A2(new_n248), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT0), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G85gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(KEYINPUT6), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT85), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n271), .B1(new_n261), .B2(new_n266), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT6), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT6), .B1(new_n267), .B2(new_n272), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n266), .A3(new_n271), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(KEYINPUT84), .A3(new_n280), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n278), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n289), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n290), .B2(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  AND2_X1   g092(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(G190gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n286), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n289), .A2(G169gat), .A3(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT23), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n297), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n293), .A2(new_n292), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT64), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n305), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT64), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n303), .A2(new_n309), .A3(KEYINPUT25), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n296), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G183gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT27), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G183gat), .ZN(new_n315));
  INV_X1    g114(.A(G190gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT27), .B(G183gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT28), .A3(new_n316), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n300), .A2(new_n323), .A3(new_n301), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n287), .A2(KEYINPUT26), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n324), .A2(new_n292), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(G226gat), .B(G233gat), .C1(new_n311), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G226gat), .A2(G233gat), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n296), .A2(new_n310), .B1(new_n322), .B2(new_n326), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(KEYINPUT29), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G211gat), .A2(G218gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT22), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(KEYINPUT72), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G211gat), .B(G218gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(KEYINPUT72), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n338), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n344), .A2(new_n345), .B1(new_n341), .B2(KEYINPUT72), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n341), .A2(KEYINPUT72), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n339), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n333), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n340), .B1(new_n338), .B2(new_n342), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n339), .A3(new_n347), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(KEYINPUT73), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  NAND3_X1  g157(.A1(new_n328), .A2(new_n331), .A3(new_n353), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n361), .A2(KEYINPUT30), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(new_n359), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n358), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n355), .A2(KEYINPUT74), .A3(new_n359), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(KEYINPUT30), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT88), .B1(new_n285), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n296), .A2(new_n310), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n322), .A2(new_n326), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT68), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n372), .A2(new_n250), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n250), .B2(new_n330), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT34), .ZN(new_n378));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n372), .A2(new_n250), .A3(new_n373), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT68), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n247), .B1(new_n311), .B2(new_n327), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n375), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n379), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT34), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n374), .B1(new_n330), .B2(new_n250), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n385), .B1(new_n376), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT32), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G15gat), .B(G43gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT69), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G71gat), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n394), .A2(KEYINPUT69), .ZN(new_n397));
  INV_X1    g196(.A(G71gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(KEYINPUT69), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n396), .A2(new_n400), .A3(G99gat), .ZN(new_n401));
  AOI21_X1  g200(.A(G99gat), .B1(new_n396), .B2(new_n400), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n391), .A2(new_n393), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT32), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n384), .B2(new_n385), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT33), .B1(new_n384), .B2(new_n385), .ZN(new_n407));
  INV_X1    g206(.A(new_n403), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n388), .B1(new_n404), .B2(new_n409), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(KEYINPUT35), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT29), .B1(new_n251), .B2(new_n225), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT80), .B1(new_n353), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n226), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n352), .A4(new_n349), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n350), .B2(new_n351), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n223), .B1(new_n422), .B2(KEYINPUT3), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT79), .B(new_n223), .C1(new_n422), .C2(KEYINPUT3), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n417), .A2(new_n421), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G228gat), .A2(G233gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n423), .B(new_n430), .C1(new_n353), .C2(new_n416), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT81), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n419), .A2(new_n352), .A3(new_n349), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n430), .A4(new_n423), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G22gat), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n429), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n429), .B2(new_n436), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n440));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT31), .B(G50gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NOR4_X1   g243(.A1(new_n438), .A2(new_n439), .A3(new_n440), .A4(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n438), .A2(new_n439), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n446), .B2(KEYINPUT82), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n440), .B1(new_n438), .B2(new_n439), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND4_X1   g248(.A1(new_n276), .A2(new_n267), .A3(KEYINPUT6), .A4(new_n272), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n276), .B1(new_n275), .B2(KEYINPUT6), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n279), .A2(KEYINPUT84), .A3(new_n280), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT84), .B1(new_n279), .B2(new_n280), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n456));
  INV_X1    g255(.A(new_n370), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n371), .A2(new_n415), .A3(new_n449), .A4(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n281), .A2(new_n273), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(new_n370), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT70), .B1(new_n382), .B2(new_n386), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n404), .A2(new_n462), .A3(new_n409), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n404), .B2(new_n409), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n262), .A2(new_n248), .A3(new_n263), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n249), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(KEYINPUT83), .A3(new_n249), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT39), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n259), .A2(new_n249), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n472), .A2(KEYINPUT39), .A3(new_n473), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n271), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n275), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT40), .A4(new_n271), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n370), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n449), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n355), .A2(new_n486), .A3(new_n359), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n358), .A2(KEYINPUT38), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n363), .A2(KEYINPUT37), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n361), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n452), .B(new_n491), .C1(new_n453), .C2(new_n454), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n365), .A2(KEYINPUT37), .A3(new_n367), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n366), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n496), .A3(new_n366), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n487), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(KEYINPUT86), .A2(new_n492), .B1(new_n498), .B2(KEYINPUT38), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n283), .A2(new_n284), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n500), .A2(new_n501), .A3(new_n452), .A4(new_n491), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n485), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT36), .B1(new_n463), .B2(new_n464), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n505));
  AOI221_X4 g304(.A(new_n405), .B1(new_n403), .B2(KEYINPUT33), .C1(new_n384), .C2(new_n385), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n387), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT36), .B1(new_n507), .B2(new_n410), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI211_X1 g309(.A(KEYINPUT71), .B(KEYINPUT36), .C1(new_n507), .C2(new_n410), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n429), .A2(new_n436), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G22gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n429), .A2(new_n436), .A3(new_n437), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(KEYINPUT82), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n448), .A2(new_n517), .A3(new_n444), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n446), .A2(KEYINPUT82), .A3(new_n443), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n281), .A2(new_n273), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n457), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n513), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n468), .B1(new_n503), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G169gat), .B(G197gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT12), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  INV_X1    g332(.A(G43gat), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT92), .B1(new_n534), .B2(G50gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(G50gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G50gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G43gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(KEYINPUT92), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n533), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT93), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT94), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n539), .A2(new_n536), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n533), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n551), .B2(new_n550), .ZN(new_n553));
  NAND2_X1  g352(.A1(G29gat), .A2(G36gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n542), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n547), .A2(KEYINPUT91), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n557), .A2(new_n546), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n547), .A2(KEYINPUT91), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n558), .A2(new_n559), .B1(G29gat), .B2(G36gat), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n560), .A2(new_n553), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT17), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(G1gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(KEYINPUT16), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  OAI221_X1 g365(.A(new_n565), .B1(new_n566), .B2(G8gat), .C1(new_n564), .C2(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(G8gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n556), .A2(new_n571), .A3(KEYINPUT17), .A4(new_n561), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n561), .B1(new_n542), .B2(new_n555), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT96), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n569), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT97), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(KEYINPUT18), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n573), .B(new_n569), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n578), .B(KEYINPUT13), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n570), .A2(new_n576), .B1(new_n573), .B2(new_n569), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n582), .B1(new_n588), .B2(new_n578), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n532), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n581), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n592), .A2(new_n583), .A3(new_n586), .A4(new_n531), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n525), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT9), .ZN(new_n600));
  INV_X1    g399(.A(G78gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n398), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G57gat), .ZN(new_n603));
  INV_X1    g402(.A(G64gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G57gat), .A2(G64gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n602), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n598), .A2(new_n599), .A3(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(KEYINPUT99), .A2(KEYINPUT100), .A3(G57gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(KEYINPUT99), .A2(G57gat), .ZN(new_n610));
  OAI21_X1  g409(.A(G64gat), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n604), .B1(new_n612), .B2(new_n603), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n611), .A2(new_n596), .A3(new_n602), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n569), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT101), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n243), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n619), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G155gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n624), .B(new_n628), .Z(new_n629));
  NAND2_X1  g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  INV_X1    g429(.A(G85gat), .ZN(new_n631));
  INV_X1    g430(.A(G92gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(KEYINPUT8), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT7), .ZN(new_n634));
  OAI211_X1 g433(.A(KEYINPUT103), .B(new_n634), .C1(new_n631), .C2(new_n632), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G99gat), .B(G106gat), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n638), .A2(G85gat), .A3(G92gat), .A4(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n637), .B1(new_n636), .B2(new_n640), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n562), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n576), .ZN(new_n646));
  AND2_X1   g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n573), .A2(new_n644), .B1(KEYINPUT41), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G190gat), .B(G218gat), .Z(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n646), .B2(new_n648), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n647), .A2(KEYINPUT41), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT102), .ZN(new_n655));
  XOR2_X1   g454(.A(G134gat), .B(G162gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT104), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n651), .A2(new_n653), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660));
  OAI22_X1  g459(.A1(new_n651), .A2(new_n653), .B1(new_n660), .B2(new_n657), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n608), .A2(new_n614), .ZN(new_n663));
  INV_X1    g462(.A(new_n643), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n641), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n615), .B1(new_n642), .B2(new_n643), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n644), .A2(KEYINPUT10), .A3(new_n663), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT105), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT105), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n665), .A2(new_n666), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n672), .ZN(new_n677));
  XNOR2_X1  g476(.A(G120gat), .B(G148gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  NAND3_X1  g479(.A1(new_n675), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n671), .B(KEYINPUT106), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n668), .B2(new_n669), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n677), .ZN(new_n685));
  INV_X1    g484(.A(new_n680), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n629), .A2(new_n662), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n595), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n521), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n564), .ZN(G1324gat));
  XNOR2_X1  g493(.A(KEYINPUT107), .B(KEYINPUT16), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G8gat), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n595), .A2(new_n370), .A3(new_n691), .A4(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G8gat), .B1(new_n692), .B2(new_n457), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n697), .ZN(new_n699));
  MUX2_X1   g498(.A(new_n697), .B(new_n699), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g499(.A(G15gat), .B1(new_n692), .B2(new_n513), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n414), .A2(G15gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n692), .B2(new_n702), .ZN(G1326gat));
  NAND2_X1  g502(.A1(new_n525), .A2(new_n594), .ZN(new_n704));
  OR4_X1    g503(.A1(KEYINPUT108), .A2(new_n704), .A3(new_n449), .A4(new_n690), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT108), .B1(new_n692), .B2(new_n449), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  XNOR2_X1  g508(.A(new_n624), .B(new_n628), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n689), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n704), .A2(new_n662), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n544), .A3(new_n460), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n449), .B2(new_n461), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT109), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n512), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n492), .A2(KEYINPUT86), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n498), .A2(KEYINPUT38), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n502), .A3(new_n721), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n449), .A2(new_n484), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n719), .A2(new_n724), .B1(new_n467), .B2(new_n459), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n715), .B1(new_n725), .B2(new_n662), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n662), .A2(new_n715), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n525), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n711), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n726), .A2(new_n594), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n521), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n731), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n712), .A2(new_n545), .A3(new_n370), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT46), .ZN(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n730), .B2(new_n457), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(KEYINPUT46), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(G1329gat));
  NAND2_X1  g536(.A1(new_n659), .A2(new_n661), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n595), .A2(new_n738), .A3(new_n729), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n534), .B1(new_n739), .B2(new_n414), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n512), .A2(G43gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n730), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT47), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n740), .B(new_n744), .C1(new_n730), .C2(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1330gat));
  OAI21_X1  g545(.A(G50gat), .B1(new_n730), .B2(new_n449), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n449), .A2(G50gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n712), .A2(new_n748), .B1(KEYINPUT110), .B2(new_n749), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n749), .A2(KEYINPUT110), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n747), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n747), .B2(new_n750), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(G1331gat));
  INV_X1    g553(.A(new_n718), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT109), .B1(new_n520), .B2(new_n522), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n513), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n468), .B1(new_n757), .B2(new_n503), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n710), .A2(new_n738), .A3(new_n594), .A4(new_n689), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n521), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT99), .B(G57gat), .Z(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1332gat));
  AND2_X1   g562(.A1(new_n758), .A2(new_n759), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n370), .B(KEYINPUT111), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  OR2_X1    g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1333gat));
  NAND3_X1  g571(.A1(new_n764), .A2(new_n398), .A3(new_n413), .ZN(new_n773));
  OAI21_X1  g572(.A(G71gat), .B1(new_n760), .B2(new_n513), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n449), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n601), .ZN(G1335gat));
  INV_X1    g577(.A(new_n594), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n710), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT114), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n758), .A2(new_n738), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n758), .A2(KEYINPUT51), .A3(new_n738), .A4(new_n781), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(KEYINPUT115), .A3(new_n783), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n689), .A2(G85gat), .A3(new_n521), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n781), .A2(new_n688), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n726), .A2(new_n728), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792), .B2(new_n521), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(G1336gat));
  OAI21_X1  g593(.A(G92gat), .B1(new_n792), .B2(new_n457), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n784), .A2(new_n786), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n766), .A2(G92gat), .A3(new_n689), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n787), .A2(new_n788), .A3(new_n797), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  OAI21_X1  g601(.A(G92gat), .B1(new_n792), .B2(new_n766), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(G1337gat));
  NOR2_X1   g604(.A1(new_n414), .A2(new_n689), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(G99gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n788), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(G99gat), .B1(new_n792), .B2(new_n513), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1338gat));
  NOR3_X1   g610(.A1(new_n449), .A2(G106gat), .A3(new_n689), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n787), .A2(new_n788), .A3(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n726), .A2(new_n520), .A3(new_n728), .A4(new_n791), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT53), .B1(new_n814), .B2(G106gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n814), .A2(new_n817), .A3(G106gat), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n814), .B2(G106gat), .ZN(new_n819));
  INV_X1    g618(.A(new_n812), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n784), .B2(new_n786), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n668), .A2(new_n669), .A3(new_n682), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n673), .B2(new_n674), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n680), .B1(new_n683), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n825), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n674), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n670), .A3(new_n672), .ZN(new_n834));
  OAI211_X1 g633(.A(KEYINPUT55), .B(new_n830), .C1(new_n834), .C2(new_n827), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n681), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n590), .B2(new_n593), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n588), .A2(new_n578), .B1(new_n584), .B2(new_n585), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n530), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n593), .A2(new_n688), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n662), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n593), .A2(new_n839), .ZN(new_n842));
  INV_X1    g641(.A(new_n836), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n738), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n629), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n690), .A2(new_n594), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n521), .A3(new_n520), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n766), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(new_n465), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n230), .A3(new_n594), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n848), .A2(new_n594), .A3(new_n413), .A4(new_n766), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(G113gat), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n853), .A2(new_n852), .A3(G113gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(G1340gat));
  NAND2_X1  g655(.A1(new_n850), .A2(new_n688), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n807), .A2(new_n238), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n857), .A2(new_n238), .B1(new_n849), .B2(new_n858), .ZN(G1341gat));
  NOR2_X1   g658(.A1(new_n235), .A2(new_n236), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n850), .A2(new_n860), .A3(new_n629), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n849), .A2(new_n413), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n710), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n860), .B2(new_n863), .ZN(G1342gat));
  NAND2_X1  g663(.A1(new_n738), .A2(new_n457), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT118), .Z(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n848), .A2(new_n244), .A3(new_n465), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT56), .Z(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n862), .B2(new_n662), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1343gat));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n520), .B1(new_n845), .B2(new_n846), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n513), .A2(new_n460), .A3(new_n766), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n594), .A2(new_n205), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT121), .Z(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n872), .B1(new_n878), .B2(KEYINPUT120), .ZN(new_n879));
  INV_X1    g678(.A(new_n874), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT119), .B1(new_n837), .B2(new_n840), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n594), .A2(new_n843), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n593), .A2(new_n688), .A3(new_n839), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n882), .A2(new_n886), .A3(new_n662), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n629), .B1(new_n887), .B2(new_n844), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n520), .B1(new_n888), .B2(new_n846), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n881), .B1(KEYINPUT57), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n205), .B1(new_n890), .B2(new_n594), .ZN(new_n891));
  INV_X1    g690(.A(new_n878), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n879), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n881), .ZN(new_n894));
  INV_X1    g693(.A(new_n889), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n894), .B(new_n594), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G141gat), .ZN(new_n898));
  INV_X1    g697(.A(new_n879), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n878), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n893), .A2(new_n900), .ZN(G1344gat));
  NAND3_X1  g700(.A1(new_n875), .A2(new_n206), .A3(new_n688), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  INV_X1    g703(.A(new_n846), .ZN(new_n905));
  INV_X1    g704(.A(new_n844), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n837), .A2(new_n840), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n738), .B1(new_n907), .B2(new_n884), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n908), .B2(new_n882), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n904), .B(new_n905), .C1(new_n909), .C2(new_n629), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n888), .B2(new_n846), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n449), .A2(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n913), .A2(new_n688), .A3(new_n880), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n903), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n206), .C1(new_n890), .C2(new_n688), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n902), .B1(new_n916), .B2(new_n917), .ZN(G1345gat));
  NAND2_X1  g717(.A1(new_n875), .A2(new_n629), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n217), .ZN(new_n920));
  INV_X1    g719(.A(new_n890), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n629), .A2(G155gat), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT123), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n926), .B(new_n920), .C1(new_n921), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1346gat));
  AOI21_X1  g727(.A(new_n218), .B1(new_n890), .B2(new_n738), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n513), .A2(new_n460), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n873), .A2(new_n866), .A3(G162gat), .A4(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT125), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n894), .B(new_n738), .C1(new_n895), .C2(new_n896), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G162gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935));
  INV_X1    g734(.A(new_n931), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n932), .A2(new_n937), .ZN(G1347gat));
  NAND2_X1  g737(.A1(new_n765), .A2(new_n521), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n465), .A3(new_n449), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n847), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G169gat), .B1(new_n942), .B2(new_n594), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n414), .A2(new_n460), .A3(new_n457), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n449), .B(new_n944), .C1(new_n845), .C2(new_n846), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n945), .A2(new_n298), .A3(new_n779), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n943), .A2(new_n946), .ZN(G1348gat));
  NAND3_X1  g746(.A1(new_n942), .A2(new_n299), .A3(new_n688), .ZN(new_n948));
  OAI21_X1  g747(.A(G176gat), .B1(new_n945), .B2(new_n689), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1349gat));
  AOI21_X1  g749(.A(KEYINPUT127), .B1(KEYINPUT126), .B2(KEYINPUT60), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n942), .A2(new_n320), .A3(new_n629), .ZN(new_n953));
  OAI21_X1  g752(.A(G183gat), .B1(new_n945), .B2(new_n710), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n957), .B1(new_n952), .B2(new_n955), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n945), .B2(new_n662), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT61), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n316), .A3(new_n738), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1351gat));
  AND2_X1   g761(.A1(new_n913), .A2(new_n914), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n512), .A2(new_n460), .A3(new_n457), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(G197gat), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n779), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n873), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n513), .A3(new_n940), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n969), .A2(new_n779), .ZN(new_n970));
  AOI22_X1  g769(.A1(new_n965), .A2(new_n967), .B1(new_n966), .B2(new_n970), .ZN(G1352gat));
  NAND3_X1  g770(.A1(new_n963), .A2(new_n688), .A3(new_n964), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(G204gat), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n969), .A2(G204gat), .A3(new_n689), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1353gat));
  OR3_X1    g775(.A1(new_n969), .A2(G211gat), .A3(new_n710), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n913), .A2(new_n629), .A3(new_n914), .A4(new_n964), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n738), .A3(new_n964), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G218gat), .ZN(new_n983));
  OR3_X1    g782(.A1(new_n969), .A2(G218gat), .A3(new_n662), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


