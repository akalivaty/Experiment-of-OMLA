//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n203));
  NAND2_X1  g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT7), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G85gat), .ZN(new_n207));
  INV_X1    g006(.A(G92gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n203), .A2(new_n206), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G99gat), .B(G106gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(KEYINPUT8), .A2(new_n202), .B1(new_n207), .B2(new_n208), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n215), .A2(new_n212), .A3(new_n206), .A4(new_n210), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(KEYINPUT101), .A3(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n206), .A2(new_n210), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT101), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n218), .A2(new_n219), .A3(new_n212), .A4(new_n215), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT10), .ZN(new_n222));
  NAND2_X1  g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  INV_X1    g022(.A(G71gat), .ZN(new_n224));
  INV_X1    g023(.A(G78gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G57gat), .B(G64gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n223), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(G71gat), .A2(G78gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G71gat), .A2(G78gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT97), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT97), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n226), .A2(new_n233), .A3(new_n223), .ZN(new_n234));
  INV_X1    g033(.A(G64gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G57gat), .ZN(new_n236));
  INV_X1    g035(.A(G57gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G64gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n234), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT98), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n230), .B2(KEYINPUT9), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n223), .A2(KEYINPUT98), .A3(new_n228), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n229), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n221), .A2(new_n222), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n245), .A3(new_n220), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT105), .ZN(new_n249));
  INV_X1    g048(.A(new_n245), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n216), .A3(new_n214), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT105), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n217), .A2(new_n245), .A3(new_n252), .A4(new_n220), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n249), .A2(new_n222), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n254), .A2(KEYINPUT106), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(KEYINPUT106), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n247), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G230gat), .A2(G233gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT107), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n249), .A2(new_n253), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n262), .A2(new_n251), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n261), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G204gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(new_n269), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT94), .ZN(new_n273));
  XNOR2_X1  g072(.A(G15gat), .B(G22gat), .ZN(new_n274));
  INV_X1    g073(.A(G1gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT16), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n274), .A2(G1gat), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n277), .A2(new_n278), .A3(G8gat), .ZN(new_n279));
  INV_X1    g078(.A(G8gat), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n274), .A2(G1gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n276), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n273), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(G8gat), .B1(new_n277), .B2(new_n278), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n280), .A3(new_n282), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT94), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G43gat), .B(G50gat), .Z(new_n289));
  INV_X1    g088(.A(KEYINPUT15), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(KEYINPUT91), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G43gat), .B(G50gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT15), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G29gat), .A2(G36gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT14), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G29gat), .A2(G36gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT92), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n291), .A2(new_n294), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n295), .B(KEYINPUT14), .ZN(new_n301));
  INV_X1    g100(.A(new_n298), .ZN(new_n302));
  OAI211_X1 g101(.A(KEYINPUT15), .B(new_n292), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G229gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT17), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n304), .B(new_n307), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT93), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT93), .B1(new_n285), .B2(new_n286), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n305), .B(new_n306), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT18), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n300), .A2(new_n303), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n284), .B2(new_n287), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n304), .B(KEYINPUT17), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n309), .A2(new_n310), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT18), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n319), .A3(new_n306), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n306), .B(KEYINPUT13), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n284), .A2(new_n314), .A3(new_n287), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(new_n315), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT95), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT95), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n326), .B(new_n322), .C1(new_n323), .C2(new_n315), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n313), .A2(new_n320), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G113gat), .B(G141gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G169gat), .B(G197gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT90), .B(KEYINPUT12), .Z(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  NOR2_X1   g134(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n313), .A2(new_n320), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n325), .A2(new_n327), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT96), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT96), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n328), .A2(new_n341), .A3(new_n335), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n336), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n272), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n288), .B1(KEYINPUT21), .B2(new_n250), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT100), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n347), .ZN(new_n349));
  NAND2_X1  g148(.A1(G231gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n348), .B2(new_n349), .ZN(new_n354));
  XNOR2_X1  g153(.A(G127gat), .B(G155gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n355), .B(KEYINPUT20), .Z(new_n356));
  NOR3_X1   g155(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G183gat), .B(G211gat), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT99), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT19), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT21), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n245), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n361), .B(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n356), .B1(new_n353), .B2(new_n354), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n358), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n358), .B2(new_n365), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G134gat), .B(G162gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT41), .ZN(new_n370));
  INV_X1    g169(.A(G232gat), .ZN(new_n371));
  INV_X1    g170(.A(G233gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n369), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n316), .A2(new_n221), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n221), .A2(new_n314), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(G190gat), .B(G218gat), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT102), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT102), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n375), .A2(new_n383), .A3(new_n378), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT103), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n374), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n379), .A2(new_n381), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n387), .B(new_n389), .Z(new_n390));
  OAI21_X1  g189(.A(KEYINPUT104), .B1(new_n368), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n366), .A2(new_n367), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT104), .ZN(new_n393));
  INV_X1    g192(.A(new_n390), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n397));
  INV_X1    g196(.A(G226gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(new_n372), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OR2_X1    g199(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT68), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT68), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(new_n405), .A3(new_n402), .ZN(new_n406));
  AOI21_X1  g205(.A(G190gat), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT28), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G190gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n403), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT69), .ZN(new_n415));
  NOR2_X1   g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT66), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT66), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(G169gat), .B2(G176gat), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT26), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n413), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  OR3_X1    g224(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT24), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(G183gat), .B2(G190gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n412), .A2(KEYINPUT24), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n426), .B(new_n427), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT23), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n416), .A2(KEYINPUT23), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n431), .A2(new_n424), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT25), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n412), .A2(KEYINPUT24), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n412), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n428), .A2(G183gat), .A3(G190gat), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n412), .A2(new_n438), .A3(KEYINPUT24), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n441), .B(new_n442), .C1(G183gat), .C2(G190gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n417), .A2(new_n419), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n435), .B1(new_n444), .B2(KEYINPUT23), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n443), .A2(new_n445), .A3(new_n424), .A4(new_n433), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n409), .A2(new_n425), .B1(new_n436), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n400), .B1(new_n447), .B2(KEYINPUT29), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT73), .B(G204gat), .ZN(new_n449));
  INV_X1    g248(.A(G197gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT22), .ZN(new_n452));
  INV_X1    g251(.A(G211gat), .ZN(new_n453));
  INV_X1    g252(.A(G218gat), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(G211gat), .B(G218gat), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(KEYINPUT74), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n451), .B(new_n455), .C1(KEYINPUT74), .C2(new_n458), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n436), .A2(new_n446), .ZN(new_n463));
  INV_X1    g262(.A(new_n420), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n414), .B(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n466), .A3(new_n424), .ZN(new_n467));
  INV_X1    g266(.A(new_n413), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(new_n468), .C1(new_n408), .C2(new_n407), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n400), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n448), .A2(new_n462), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT77), .ZN(new_n473));
  INV_X1    g272(.A(new_n462), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n448), .B2(new_n471), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n463), .A2(new_n469), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT29), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n399), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(KEYINPUT75), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT76), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT75), .B1(new_n479), .B2(new_n470), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n448), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(KEYINPUT76), .A3(new_n474), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n473), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G8gat), .B(G36gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(new_n235), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(new_n208), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT78), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT77), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n472), .B(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT76), .B1(new_n486), .B2(new_n474), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n482), .B(new_n462), .C1(new_n484), .C2(new_n485), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT78), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n491), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT82), .B(G155gat), .Z(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G162gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(G155gat), .A2(G162gat), .ZN(new_n504));
  OR2_X1    g303(.A1(G155gat), .A2(G162gat), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n503), .A2(KEYINPUT2), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G148gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G141gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n509), .A2(KEYINPUT81), .ZN(new_n510));
  INV_X1    g309(.A(G141gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G148gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(KEYINPUT81), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n504), .A2(new_n515), .A3(KEYINPUT2), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n504), .B2(KEYINPUT2), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n512), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(new_n509), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n504), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT79), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n506), .A2(new_n514), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G113gat), .B(G120gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT1), .ZN(new_n525));
  XNOR2_X1  g324(.A(G127gat), .B(G134gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G134gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n525), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT1), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n523), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n506), .A2(new_n514), .ZN(new_n535));
  INV_X1    g334(.A(new_n522), .ZN(new_n536));
  INV_X1    g335(.A(new_n520), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT3), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n531), .A2(new_n532), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT3), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n535), .B(new_n541), .C1(new_n536), .C2(new_n537), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G225gat), .A2(G233gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n533), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n534), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT5), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n538), .A2(new_n540), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n533), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n543), .A3(new_n548), .A4(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT0), .B(G57gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G85gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(G1gat), .B(G29gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n552), .A2(new_n558), .A3(new_n553), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n554), .A2(KEYINPUT6), .A3(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n498), .A2(new_n491), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT30), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n488), .A2(new_n492), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n501), .A2(new_n565), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n542), .A2(new_n478), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n474), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT29), .B1(new_n460), .B2(new_n461), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n538), .B1(new_n574), .B2(KEYINPUT3), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n573), .A2(new_n575), .A3(G228gat), .A4(G233gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(G228gat), .A2(G233gat), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n462), .B1(new_n542), .B2(new_n478), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n456), .A2(new_n458), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n451), .A2(new_n457), .A3(new_n455), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n478), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n523), .B1(new_n581), .B2(new_n541), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n577), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G50gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G78gat), .ZN(new_n587));
  INV_X1    g386(.A(G106gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(G22gat), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G22gat), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n576), .A2(new_n583), .A3(new_n592), .A4(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(new_n590), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(new_n595), .A3(new_n596), .A4(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n571), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT34), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT71), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n477), .B(new_n540), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n602), .A2(KEYINPUT72), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(G227gat), .A2(G233gat), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT72), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n603), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT71), .B(new_n602), .C1(new_n604), .C2(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n604), .A2(new_n607), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G15gat), .B(G43gat), .Z(new_n617));
  XNOR2_X1  g416(.A(G71gat), .B(G99gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n614), .A2(KEYINPUT32), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n616), .A3(new_n619), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n613), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n612), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n625), .A2(new_n628), .A3(KEYINPUT36), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT36), .B1(new_n625), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n601), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n634), .B(new_n495), .C1(new_n496), .C2(new_n497), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT87), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n483), .A2(new_n487), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n638), .A2(KEYINPUT87), .A3(new_n634), .A4(new_n495), .ZN(new_n639));
  AND4_X1   g438(.A1(new_n633), .A2(new_n637), .A3(new_n491), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n486), .A2(new_n462), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n448), .A2(new_n474), .A3(new_n471), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(KEYINPUT37), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n565), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n498), .A2(KEYINPUT37), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n637), .A2(new_n645), .A3(new_n639), .A4(new_n491), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n566), .B1(new_n646), .B2(KEYINPUT38), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n600), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT39), .B1(new_n550), .B2(new_n545), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT85), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n534), .A2(new_n543), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n651), .B(new_n652), .C1(new_n653), .C2(new_n544), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n544), .B1(new_n534), .B2(new_n543), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n559), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT86), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT40), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n567), .A2(new_n570), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n493), .A2(new_n500), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n560), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n632), .B1(new_n648), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n568), .B(KEYINPUT30), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n600), .B1(new_n628), .B2(new_n625), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n664), .A2(new_n665), .A3(new_n565), .A4(new_n501), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT35), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n397), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n600), .ZN(new_n670));
  INV_X1    g469(.A(new_n565), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n637), .A2(new_n639), .A3(new_n633), .A4(new_n491), .ZN(new_n672));
  INV_X1    g471(.A(new_n643), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n646), .A2(KEYINPUT38), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n568), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n662), .B(new_n670), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n601), .A3(new_n631), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n666), .B(KEYINPUT35), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(KEYINPUT88), .A3(new_n679), .ZN(new_n680));
  AOI211_X1 g479(.A(new_n345), .B(new_n396), .C1(new_n669), .C2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n671), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  INV_X1    g482(.A(new_n681), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n660), .A2(new_n661), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT42), .B1(new_n686), .B2(new_n280), .ZN(new_n687));
  INV_X1    g486(.A(new_n685), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT108), .B(G8gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT16), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n681), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  MUX2_X1   g490(.A(KEYINPUT42), .B(new_n687), .S(new_n691), .Z(G1325gat));
  INV_X1    g491(.A(new_n625), .ZN(new_n693));
  INV_X1    g492(.A(new_n628), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(G15gat), .B1(new_n681), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n684), .A2(new_n631), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(new_n698), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n600), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NAND2_X1  g501(.A1(new_n669), .A2(new_n680), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n390), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n345), .A2(new_n392), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(G29gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n671), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n678), .A2(new_n679), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n390), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n394), .B1(new_n669), .B2(new_n680), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(new_n565), .A3(new_n706), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n710), .B1(new_n708), .B2(new_n717), .ZN(G1328gat));
  INV_X1    g517(.A(G36gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n707), .A2(new_n719), .A3(new_n688), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT46), .Z(new_n721));
  NOR3_X1   g520(.A1(new_n716), .A2(new_n685), .A3(new_n706), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n719), .B2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(new_n631), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n715), .A2(new_n724), .A3(new_n705), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G43gat), .ZN(new_n726));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n727), .A3(new_n696), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1330gat));
  NOR4_X1   g530(.A1(new_n704), .A2(G50gat), .A3(new_n670), .A4(new_n706), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n715), .A2(new_n600), .A3(new_n705), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT109), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G50gat), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n734), .A2(KEYINPUT109), .ZN(new_n737));
  OAI211_X1 g536(.A(KEYINPUT48), .B(new_n733), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n734), .A2(G50gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n732), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(G1331gat));
  INV_X1    g541(.A(new_n343), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n743), .B(new_n396), .C1(new_n678), .C2(new_n679), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n272), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n565), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n237), .ZN(G1332gat));
  INV_X1    g546(.A(new_n745), .ZN(new_n748));
  NAND2_X1  g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(new_n688), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT110), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n751), .B(new_n753), .ZN(G1333gat));
  NAND3_X1  g553(.A1(new_n748), .A2(G71gat), .A3(new_n724), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n748), .A2(KEYINPUT111), .A3(new_n696), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n745), .B2(new_n695), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n755), .B1(new_n759), .B2(G71gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n670), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n225), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n392), .A2(new_n743), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n711), .A2(new_n390), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n272), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n671), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n764), .A2(new_n272), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n716), .A2(new_n207), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n772), .B1(new_n671), .B2(new_n774), .ZN(G1336gat));
  OAI211_X1 g574(.A(new_n208), .B(new_n272), .C1(new_n767), .C2(new_n768), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n685), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(KEYINPUT52), .ZN(new_n778));
  INV_X1    g577(.A(new_n773), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n712), .B1(new_n703), .B2(new_n390), .ZN(new_n780));
  INV_X1    g579(.A(new_n713), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n688), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n715), .A2(new_n784), .A3(new_n688), .A4(new_n779), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n785), .A3(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n782), .A2(new_n788), .A3(G92gat), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n782), .B2(G92gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n789), .A2(new_n790), .A3(new_n777), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(G1337gat));
  NOR3_X1   g592(.A1(new_n716), .A2(new_n631), .A3(new_n773), .ZN(new_n794));
  INV_X1    g593(.A(G99gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n695), .A2(G99gat), .A3(new_n770), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT114), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n794), .A2(new_n795), .B1(new_n769), .B2(new_n797), .ZN(G1338gat));
  NOR4_X1   g597(.A1(new_n769), .A2(G106gat), .A3(new_n770), .A4(new_n670), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n716), .A2(new_n670), .A3(new_n773), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n800), .B(new_n801), .C1(new_n588), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n716), .A2(new_n773), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n588), .B1(new_n804), .B2(new_n600), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n805), .B2(new_n799), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1339gat));
  INV_X1    g606(.A(KEYINPUT106), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n262), .A2(new_n808), .A3(new_n222), .A4(new_n251), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n254), .A2(KEYINPUT106), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n246), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n259), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n261), .A2(new_n812), .A3(KEYINPUT54), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n257), .A2(new_n814), .A3(new_n260), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n815), .A2(KEYINPUT115), .A3(new_n269), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT115), .B1(new_n815), .B2(new_n269), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n343), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT55), .B(new_n813), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT116), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n811), .A2(KEYINPUT54), .A3(new_n259), .ZN(new_n824));
  INV_X1    g623(.A(new_n269), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n815), .A2(KEYINPUT115), .A3(new_n269), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT55), .A4(new_n813), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n820), .A2(new_n822), .A3(new_n270), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n340), .A2(new_n342), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n318), .A2(new_n306), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n323), .A2(new_n315), .A3(new_n322), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n333), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT117), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n272), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n394), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n818), .A2(new_n819), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n390), .A2(new_n841), .A3(new_n832), .A4(new_n836), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n822), .A2(new_n830), .A3(new_n270), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n390), .B1(new_n831), .B2(new_n837), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT118), .B1(new_n847), .B2(new_n844), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n368), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n391), .A2(new_n395), .A3(new_n770), .A4(new_n343), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n688), .A2(new_n565), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n851), .A2(new_n665), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n743), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n272), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n392), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(G127gat), .ZN(G1342gat));
  AND2_X1   g658(.A1(new_n853), .A2(new_n390), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n529), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n862), .B(new_n863), .C1(new_n529), .C2(new_n860), .ZN(G1343gat));
  NOR2_X1   g663(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n600), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(KEYINPUT119), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n670), .B1(new_n849), .B2(new_n850), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(KEYINPUT57), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n392), .B1(new_n839), .B2(new_n845), .ZN(new_n873));
  INV_X1    g672(.A(new_n850), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT57), .B(new_n600), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n852), .A2(new_n631), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n743), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G141gat), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n871), .A2(new_n511), .A3(new_n743), .A4(new_n878), .ZN(new_n881));
  NAND2_X1  g680(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n866), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n865), .B(new_n883), .C1(new_n879), .C2(G141gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1344gat));
  XOR2_X1   g686(.A(new_n850), .B(KEYINPUT121), .Z(new_n888));
  AOI21_X1  g687(.A(KEYINPUT122), .B1(new_n839), .B2(new_n845), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n847), .A2(new_n890), .A3(new_n844), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n889), .A2(new_n891), .A3(new_n392), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n868), .B(new_n600), .C1(new_n888), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n894), .A3(new_n272), .ZN(new_n895));
  OAI21_X1  g694(.A(G148gat), .B1(new_n895), .B2(new_n877), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT59), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n876), .A2(new_n878), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n770), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(new_n507), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n871), .A2(new_n878), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n507), .A3(new_n272), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1345gat));
  AOI21_X1  g704(.A(new_n502), .B1(new_n903), .B2(new_n392), .ZN(new_n906));
  INV_X1    g705(.A(new_n899), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n392), .A2(new_n502), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(G1346gat));
  AOI21_X1  g708(.A(G162gat), .B1(new_n903), .B2(new_n390), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n907), .A2(G162gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n390), .ZN(G1347gat));
  NOR3_X1   g711(.A1(new_n685), .A2(new_n600), .A3(new_n695), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(new_n849), .B2(new_n850), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n913), .A2(new_n914), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(G169gat), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n918), .A2(new_n919), .A3(new_n565), .A4(new_n743), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n685), .A2(new_n671), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n696), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT124), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n600), .B1(new_n922), .B2(KEYINPUT124), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n851), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(new_n743), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n920), .B1(new_n928), .B2(new_n919), .ZN(G1348gat));
  NAND2_X1  g728(.A1(new_n918), .A2(new_n565), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n266), .B1(new_n930), .B2(new_n770), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n927), .A2(G176gat), .A3(new_n272), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G1349gat));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n404), .A2(new_n406), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n918), .A2(new_n565), .A3(new_n392), .A4(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n927), .A2(new_n392), .ZN(new_n939));
  INV_X1    g738(.A(G183gat), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n936), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n927), .B2(new_n392), .ZN(new_n942));
  INV_X1    g741(.A(new_n938), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT60), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n944), .ZN(G1350gat));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n390), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(G190gat), .ZN(new_n948));
  AOI211_X1 g747(.A(KEYINPUT61), .B(new_n410), .C1(new_n927), .C2(new_n390), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n390), .A2(new_n410), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n948), .A2(new_n949), .B1(new_n930), .B2(new_n950), .ZN(G1351gat));
  AND2_X1   g750(.A1(new_n893), .A2(new_n894), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n921), .A2(new_n631), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n343), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n867), .A2(new_n953), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n957), .A2(new_n450), .A3(new_n743), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1352gat));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n955), .B2(new_n770), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n952), .A2(KEYINPUT127), .A3(new_n272), .A4(new_n954), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(G204gat), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n957), .A2(new_n268), .A3(new_n272), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1353gat));
  NAND3_X1  g765(.A1(new_n957), .A2(new_n453), .A3(new_n392), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n392), .A3(new_n954), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n955), .B2(new_n394), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n454), .A3(new_n390), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


