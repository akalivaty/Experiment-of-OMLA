//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G50), .ZN(new_n206));
  INV_X1    g0006(.A(G226), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g0010(.A1(G77), .A2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT65), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n210), .B(new_n211), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n219), .B1(new_n218), .B2(new_n217), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NOR2_X1   g0025(.A1(new_n223), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(G50), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n225), .B(new_n228), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n207), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n221), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n206), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n220), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n253), .A2(new_n250), .A3(G13), .A4(G20), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(KEYINPUT8), .B(G58), .Z(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n229), .ZN(new_n260));
  AOI211_X1 g0060(.A(new_n260), .B(new_n255), .C1(new_n250), .C2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n258), .B1(new_n262), .B2(new_n257), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G223), .A2(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT77), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT77), .B1(new_n270), .B2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(G33), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n266), .B(new_n273), .C1(new_n207), .C2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G87), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n265), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n230), .B1(new_n268), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n283), .A2(new_n278), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G232), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n277), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G190), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT16), .ZN(new_n290));
  INV_X1    g0090(.A(G58), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n208), .ZN(new_n292));
  OAI21_X1  g0092(.A(G20), .B1(new_n292), .B2(new_n202), .ZN(new_n293));
  XOR2_X1   g0093(.A(new_n293), .B(KEYINPUT80), .Z(new_n294));
  INV_X1    g0094(.A(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n268), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G159), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT7), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n270), .A2(KEYINPUT77), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n267), .B1(new_n268), .B2(KEYINPUT3), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n300), .B1(new_n304), .B2(G20), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n295), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(KEYINPUT78), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT78), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n300), .C1(new_n304), .C2(G20), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(G68), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT79), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n307), .A2(KEYINPUT79), .A3(G68), .A4(new_n309), .ZN(new_n313));
  AOI211_X1 g0113(.A(new_n290), .B(new_n299), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n270), .A2(G33), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n302), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT7), .B1(new_n316), .B2(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n302), .A2(new_n315), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(new_n300), .A3(new_n295), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n208), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n290), .B1(new_n299), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n260), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n264), .B(new_n289), .C1(new_n314), .C2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n286), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT17), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n312), .A2(new_n313), .ZN(new_n329));
  INV_X1    g0129(.A(new_n299), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n323), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n263), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT17), .ZN(new_n334));
  INV_X1    g0134(.A(new_n327), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .A4(new_n289), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n328), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT18), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n299), .B1(new_n312), .B2(new_n313), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n323), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT81), .B1(new_n341), .B2(new_n263), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT81), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(new_n264), .C1(new_n314), .C2(new_n323), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n286), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(G169), .B2(new_n286), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n339), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  AOI211_X1 g0150(.A(KEYINPUT18), .B(new_n348), .C1(new_n342), .C2(new_n344), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n338), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n353));
  INV_X1    g0153(.A(G150), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n268), .A2(G20), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n353), .B1(new_n354), .B2(new_n296), .C1(new_n257), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n260), .ZN(new_n358));
  XOR2_X1   g0158(.A(new_n358), .B(KEYINPUT67), .Z(new_n359));
  NAND2_X1  g0159(.A1(new_n261), .A2(G50), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n252), .A2(new_n254), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n360), .C1(G50), .C2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n316), .A2(KEYINPUT66), .A3(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT66), .ZN(new_n364));
  INV_X1    g0164(.A(G1698), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n318), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(G223), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G77), .ZN(new_n368));
  INV_X1    g0168(.A(G222), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n316), .A2(new_n365), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n367), .B1(new_n368), .B2(new_n316), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n265), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n284), .A2(G226), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n281), .ZN(new_n374));
  INV_X1    g0174(.A(G169), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n362), .B(new_n376), .C1(G179), .C2(new_n374), .ZN(new_n377));
  XOR2_X1   g0177(.A(new_n377), .B(KEYINPUT69), .Z(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n262), .B2(new_n368), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n255), .A2(new_n368), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n261), .A2(KEYINPUT71), .A3(G77), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n257), .A2(new_n296), .B1(new_n295), .B2(new_n368), .ZN(new_n384));
  XOR2_X1   g0184(.A(KEYINPUT15), .B(G87), .Z(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n356), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n260), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n381), .A2(new_n382), .A3(new_n383), .A4(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n363), .A2(G238), .A3(new_n366), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n316), .A2(G232), .A3(new_n365), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n318), .A2(G107), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n393), .A2(KEYINPUT70), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(KEYINPUT70), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n265), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n280), .B1(new_n284), .B2(G244), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n389), .B1(new_n398), .B2(G200), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n287), .B2(new_n398), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n352), .A2(new_n379), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n362), .B(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n374), .A2(G200), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT10), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n405), .B1(KEYINPUT72), .B2(KEYINPUT9), .C1(new_n287), .C2(new_n374), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n404), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT10), .B(new_n407), .C1(new_n403), .C2(new_n409), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n316), .A2(G232), .A3(G1698), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n414), .B1(new_n268), .B2(new_n213), .C1(new_n370), .C2(new_n207), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n265), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n284), .A2(G238), .ZN(new_n417));
  XOR2_X1   g0217(.A(new_n280), .B(KEYINPUT74), .Z(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT13), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n416), .A2(new_n422), .A3(new_n417), .A4(new_n418), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n419), .A2(KEYINPUT75), .A3(KEYINPUT13), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(G169), .A3(new_n425), .ZN(new_n426));
  XOR2_X1   g0226(.A(KEYINPUT76), .B(KEYINPUT14), .Z(new_n427));
  AND2_X1   g0227(.A1(new_n420), .A2(new_n423), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n426), .A2(new_n427), .B1(G179), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT14), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n424), .A2(G169), .A3(new_n425), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n261), .A2(G68), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n356), .A2(new_n368), .B1(new_n206), .B2(new_n296), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n295), .A2(G68), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n260), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT11), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n255), .A2(new_n208), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT12), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n437), .A2(new_n438), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n434), .A2(new_n439), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n428), .A2(G190), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n424), .A2(G200), .A3(new_n425), .ZN(new_n446));
  INV_X1    g0246(.A(new_n443), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n398), .A2(new_n375), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n396), .A2(new_n346), .A3(new_n397), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(new_n389), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n413), .A2(new_n444), .A3(new_n448), .A4(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n401), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n318), .A2(G20), .A3(new_n275), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(KEYINPUT22), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  NAND2_X1  g0257(.A1(KEYINPUT22), .A2(G87), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n273), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n295), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n295), .A2(G107), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT23), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n456), .A2(new_n460), .A3(KEYINPUT24), .A4(new_n462), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n260), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT88), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n361), .A2(G107), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT25), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n260), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n250), .A2(G33), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n361), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT82), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n361), .A2(new_n477), .A3(new_n473), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n472), .B1(new_n479), .B2(G107), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n469), .A2(new_n470), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n468), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n215), .B1(new_n476), .B2(new_n478), .ZN(new_n484));
  NOR4_X1   g0284(.A1(new_n484), .A2(new_n472), .A3(KEYINPUT88), .A4(new_n481), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n467), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G45), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(G1), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n265), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G264), .ZN(new_n491));
  INV_X1    g0291(.A(new_n488), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n279), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n489), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT89), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n304), .A2(new_n496), .A3(G250), .A4(new_n365), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n365), .B(new_n269), .C1(new_n271), .C2(new_n272), .ZN(new_n498));
  INV_X1    g0298(.A(G250), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT89), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n304), .A2(G257), .A3(G1698), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT90), .B(G294), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G33), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n497), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n495), .B1(new_n504), .B2(new_n265), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G179), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n506), .A2(KEYINPUT91), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(KEYINPUT91), .C1(new_n375), .C2(new_n505), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n486), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n479), .A2(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n482), .A3(new_n471), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n480), .A2(new_n468), .A3(new_n482), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n505), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G200), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n505), .A2(G190), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n514), .A2(new_n467), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n509), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n295), .C1(G33), .C2(new_n213), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n220), .A2(G20), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n260), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n521), .A2(new_n260), .A3(KEYINPUT20), .A4(new_n522), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n526), .B1(new_n255), .B2(new_n220), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n361), .A2(G116), .A3(new_n473), .A4(new_n474), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n214), .A2(new_n365), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n269), .B(new_n531), .C1(new_n271), .C2(new_n272), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n365), .A2(G264), .ZN(new_n533));
  INV_X1    g0333(.A(G303), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n316), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n265), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n490), .A2(G270), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n494), .A3(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n530), .A2(new_n538), .A3(new_n346), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT21), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n375), .B1(new_n527), .B2(new_n528), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n540), .A3(new_n538), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n539), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n536), .A2(new_n537), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(G190), .A3(new_n494), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n529), .B1(new_n538), .B2(G200), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT87), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT87), .B1(new_n547), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(new_n269), .C1(new_n271), .C2(new_n272), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(G1698), .ZN(new_n555));
  AND2_X1   g0355(.A1(KEYINPUT4), .A2(G244), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n302), .A2(new_n315), .A3(new_n556), .A4(new_n365), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n302), .A2(new_n315), .A3(G250), .A4(G1698), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n557), .A2(new_n558), .A3(new_n520), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n265), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT83), .ZN(new_n562));
  XOR2_X1   g0362(.A(KEYINPUT5), .B(G41), .Z(new_n563));
  OAI21_X1  g0363(.A(new_n283), .B1(new_n563), .B2(new_n492), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n564), .B2(new_n214), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n490), .A2(KEYINPUT83), .A3(G257), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(new_n567), .A3(new_n494), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n255), .A2(new_n213), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n297), .A2(G77), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n215), .A2(KEYINPUT6), .A3(G97), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n213), .A2(new_n215), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n572), .B1(new_n575), .B2(KEYINPUT6), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G20), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n571), .B(new_n577), .C1(new_n320), .C2(new_n215), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n260), .B1(new_n479), .B2(G97), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n561), .A2(new_n567), .A3(G190), .A4(new_n494), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n569), .A2(new_n570), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n260), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n479), .A2(G97), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n570), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n568), .A2(new_n375), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n561), .A2(new_n567), .A3(new_n346), .A4(new_n494), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n552), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT84), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n457), .B1(new_n554), .B2(new_n365), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n498), .A2(new_n209), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n303), .A2(new_n302), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n594), .A2(G238), .A3(new_n365), .A4(new_n269), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(G244), .A3(G1698), .A4(new_n269), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT84), .A4(new_n457), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n265), .ZN(new_n599));
  INV_X1    g0399(.A(new_n493), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n283), .A2(G250), .A3(new_n492), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT85), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n283), .B1(new_n593), .B2(new_n597), .ZN(new_n605));
  INV_X1    g0405(.A(new_n601), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n605), .A2(new_n493), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT85), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n604), .A2(new_n608), .A3(new_n375), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n493), .B1(new_n598), .B2(new_n265), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT85), .B1(new_n610), .B2(new_n601), .ZN(new_n611));
  NOR4_X1   g0411(.A1(new_n605), .A2(new_n603), .A3(new_n493), .A4(new_n606), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n346), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n295), .A2(new_n614), .B1(new_n574), .B2(new_n275), .ZN(new_n615));
  XOR2_X1   g0415(.A(new_n615), .B(KEYINPUT86), .Z(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n356), .B2(new_n213), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n304), .A2(new_n295), .A3(G68), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(new_n260), .B1(new_n255), .B2(new_n386), .ZN(new_n621));
  INV_X1    g0421(.A(new_n479), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n386), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n609), .A2(new_n613), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n604), .A2(new_n608), .A3(G200), .ZN(new_n625));
  OAI21_X1  g0425(.A(G190), .B1(new_n611), .B2(new_n612), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n479), .A2(G87), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n519), .A2(new_n589), .A3(new_n624), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n454), .A2(new_n630), .ZN(G372));
  INV_X1    g0431(.A(KEYINPUT92), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n628), .B(new_n632), .C1(new_n326), .C2(new_n607), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n326), .B1(new_n610), .B2(new_n601), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n621), .A2(new_n627), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT92), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n626), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n602), .A2(new_n375), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n613), .A2(new_n623), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  INV_X1    g0441(.A(new_n587), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n639), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n624), .A2(new_n629), .A3(new_n642), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n509), .A2(new_n545), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n637), .A2(new_n647), .A3(new_n518), .A4(new_n639), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n643), .B(new_n646), .C1(new_n588), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n453), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(KEYINPUT18), .B(new_n349), .C1(new_n341), .C2(new_n263), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n339), .B1(new_n333), .B2(new_n348), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n447), .B1(new_n429), .B2(new_n432), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT93), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n451), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n449), .A2(KEYINPUT93), .A3(new_n450), .A4(new_n389), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n337), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n448), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n653), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n378), .B1(new_n661), .B2(new_n413), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n650), .A2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(G330), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n546), .A2(G179), .A3(new_n494), .A4(new_n529), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n541), .A2(new_n540), .A3(new_n538), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n542), .ZN(new_n667));
  INV_X1    g0467(.A(new_n551), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n549), .ZN(new_n669));
  INV_X1    g0469(.A(G13), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G20), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n250), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n669), .B1(new_n530), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n667), .A2(new_n529), .A3(new_n677), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n664), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n509), .A2(new_n518), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n678), .B1(new_n514), .B2(new_n467), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n509), .B2(new_n678), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT94), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n545), .A2(new_n677), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n519), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n509), .A2(new_n677), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n686), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n226), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n574), .A2(new_n275), .A3(new_n220), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n694), .A2(new_n695), .A3(new_n250), .ZN(new_n696));
  INV_X1    g0496(.A(new_n232), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT28), .Z(new_n699));
  NAND2_X1  g0499(.A1(new_n649), .A2(new_n678), .ZN(new_n700));
  XOR2_X1   g0500(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n637), .A2(new_n642), .A3(new_n639), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT26), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n624), .A2(new_n629), .A3(new_n641), .A4(new_n642), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n639), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT98), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n588), .B(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n648), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT29), .B(new_n678), .C1(new_n706), .C2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n702), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT96), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT95), .B1(new_n630), .B2(new_n677), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n624), .A2(new_n629), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n581), .A2(new_n587), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n669), .A2(new_n509), .A3(new_n518), .A4(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n678), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n568), .B1(new_n604), .B2(new_n608), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n505), .A2(G179), .A3(new_n546), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(KEYINPUT30), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n568), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n724), .B(new_n722), .C1(new_n611), .C2(new_n612), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n607), .A2(G179), .A3(new_n724), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n515), .A3(new_n538), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n723), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n677), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT31), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n730), .A2(new_n733), .A3(new_n677), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n714), .A2(new_n720), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n713), .B1(new_n735), .B2(new_n664), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n719), .B1(new_n718), .B2(new_n678), .ZN(new_n737));
  NOR4_X1   g0537(.A1(new_n715), .A2(new_n717), .A3(KEYINPUT95), .A4(new_n677), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n733), .B1(new_n730), .B2(new_n677), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n730), .A2(new_n733), .A3(new_n677), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT96), .A3(G330), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n712), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n699), .B1(new_n744), .B2(G1), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT99), .Z(G364));
  INV_X1    g0546(.A(new_n694), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n250), .B1(new_n671), .B2(G45), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT100), .Z(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n295), .A2(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n275), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n295), .A2(new_n346), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n754), .B1(G50), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n755), .A2(new_n287), .A3(G200), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n208), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT32), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n760), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n755), .A2(G190), .A3(new_n326), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G58), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n752), .A2(new_n287), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT101), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G107), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n287), .A2(G179), .A3(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n295), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n765), .A2(new_n761), .B1(new_n213), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n755), .A2(new_n762), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n318), .B(new_n779), .C1(G77), .C2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n766), .A2(new_n769), .A3(new_n776), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n756), .B(KEYINPUT102), .ZN(new_n784));
  INV_X1    g0584(.A(new_n778), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n784), .A2(G326), .B1(new_n502), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT103), .Z(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  NOR2_X1   g0588(.A1(new_n759), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n318), .B1(new_n763), .B2(new_n790), .C1(new_n791), .C2(new_n780), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n789), .B(new_n792), .C1(G322), .C2(new_n768), .ZN(new_n793));
  INV_X1    g0593(.A(G283), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n787), .B(new_n793), .C1(new_n794), .C2(new_n774), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n753), .A2(new_n534), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n783), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n229), .B1(G20), .B2(new_n375), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n798), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n304), .A2(new_n693), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n697), .A2(new_n487), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(new_n245), .C2(new_n487), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n316), .A2(G355), .A3(new_n226), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(G116), .C2(new_n226), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n797), .A2(new_n798), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n679), .A2(new_n680), .ZN(new_n809));
  INV_X1    g0609(.A(new_n801), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n751), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n681), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n749), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n809), .A2(G330), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(G396));
  NAND3_X1  g0615(.A1(new_n658), .A2(new_n389), .A3(new_n677), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n389), .A2(new_n677), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n400), .A2(new_n451), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n700), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n649), .A2(new_n678), .A3(new_n819), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n743), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n749), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n798), .A2(new_n799), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT104), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n368), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n304), .B1(new_n206), .B2(new_n753), .C1(new_n829), .C2(new_n763), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n774), .A2(new_n208), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n757), .A2(G137), .B1(new_n781), .B2(G159), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n768), .A2(G143), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n354), .C2(new_n759), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT34), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n830), .B(new_n831), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n835), .B2(new_n834), .C1(new_n291), .C2(new_n778), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n756), .A2(new_n534), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n778), .A2(new_n213), .B1(new_n753), .B2(new_n215), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n318), .B1(new_n763), .B2(new_n791), .C1(new_n767), .C2(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(G116), .C2(new_n781), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n775), .A2(G87), .ZN(new_n843));
  INV_X1    g0643(.A(new_n759), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n844), .A2(KEYINPUT105), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(KEYINPUT105), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n842), .B(new_n843), .C1(new_n794), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n837), .B1(new_n838), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n750), .B1(new_n849), .B2(new_n798), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n828), .B(new_n850), .C1(new_n819), .C2(new_n800), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n825), .A2(new_n851), .ZN(G384));
  NOR2_X1   g0652(.A1(new_n447), .A2(new_n678), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n444), .A2(new_n448), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n654), .B2(new_n660), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n735), .A2(new_n857), .A3(new_n820), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n340), .A2(KEYINPUT16), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n473), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n263), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n861), .A2(new_n675), .B1(new_n327), .B2(new_n324), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n348), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n331), .A2(new_n332), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n343), .B1(new_n865), .B2(new_n264), .ZN(new_n866));
  AOI211_X1 g0666(.A(KEYINPUT81), .B(new_n263), .C1(new_n331), .C2(new_n332), .ZN(new_n867));
  INV_X1    g0667(.A(new_n675), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n866), .A2(new_n867), .B1(new_n349), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n324), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT37), .B1(new_n870), .B2(new_n335), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n861), .A2(new_n675), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(KEYINPUT38), .B(new_n873), .C1(new_n352), .C2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n675), .B1(new_n342), .B2(new_n344), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n324), .A2(new_n327), .B1(new_n333), .B2(new_n348), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(new_n872), .ZN(new_n881));
  INV_X1    g0681(.A(new_n878), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n337), .B2(new_n653), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n858), .A2(new_n885), .A3(KEYINPUT40), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n349), .B1(new_n866), .B2(new_n867), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT18), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n345), .A2(new_n339), .A3(new_n349), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n337), .A3(new_n889), .ZN(new_n890));
  AOI221_X4 g0690(.A(new_n877), .B1(new_n864), .B2(new_n872), .C1(new_n890), .C2(new_n874), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n874), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n892), .B2(new_n873), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT107), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n350), .A2(new_n351), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n875), .B1(new_n895), .B2(new_n337), .ZN(new_n896));
  INV_X1    g0696(.A(new_n873), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n877), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT107), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(new_n876), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n894), .A2(new_n900), .A3(new_n858), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n886), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n454), .A2(new_n735), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n903), .B(new_n904), .Z(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(G330), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT39), .B1(new_n891), .B2(new_n893), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n876), .A2(new_n884), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n444), .A2(new_n677), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n651), .A2(new_n652), .A3(new_n675), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n451), .A2(new_n677), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n857), .B1(new_n822), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n894), .A2(new_n900), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(new_n913), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n702), .A2(new_n711), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n662), .B1(new_n454), .B2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  XNOR2_X1  g0721(.A(new_n906), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n250), .B2(new_n671), .ZN(new_n923));
  OAI211_X1 g0723(.A(G20), .B(new_n230), .C1(new_n576), .C2(KEYINPUT35), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n220), .B(new_n924), .C1(KEYINPUT35), .C2(new_n576), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT36), .Z(new_n926));
  NOR2_X1   g0726(.A1(new_n201), .A2(new_n208), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT106), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n232), .A2(new_n368), .A3(new_n292), .ZN(new_n929));
  OAI211_X1 g0729(.A(G1), .B(new_n670), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n923), .A2(new_n926), .A3(new_n930), .ZN(G367));
  INV_X1    g0731(.A(new_n744), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n584), .A2(new_n677), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n708), .A2(new_n933), .B1(new_n642), .B2(new_n677), .ZN(new_n934));
  XOR2_X1   g0734(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n935));
  AND3_X1   g0735(.A1(new_n690), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n690), .B2(new_n934), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n934), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n691), .A2(new_n939), .A3(KEYINPUT45), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT45), .B1(new_n691), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n686), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n681), .A2(KEYINPUT110), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n684), .A2(new_n687), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n945), .A2(new_n688), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n946), .B2(new_n688), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n919), .A2(new_n949), .A3(new_n736), .A4(new_n742), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT111), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n942), .B(new_n686), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT111), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(new_n744), .A4(new_n949), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n932), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n694), .B(KEYINPUT41), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n748), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n708), .A2(new_n933), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT42), .B1(new_n959), .B2(new_n688), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n690), .A2(new_n961), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n960), .B1(new_n587), .B2(new_n677), .C1(new_n962), .C2(new_n959), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT108), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n628), .A2(new_n678), .ZN(new_n966));
  MUX2_X1   g0766(.A(new_n640), .B(new_n644), .S(new_n966), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n965), .A2(new_n970), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n686), .A2(new_n934), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n958), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n775), .A2(G97), .ZN(new_n978));
  INV_X1    g0778(.A(G317), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n273), .C1(new_n979), .C2(new_n763), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  INV_X1    g0781(.A(new_n847), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n982), .A2(new_n502), .B1(G311), .B2(new_n784), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n785), .A2(G107), .B1(new_n768), .B2(G303), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n753), .A2(new_n220), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(KEYINPUT46), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(KEYINPUT46), .B2(new_n985), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n981), .A2(new_n983), .A3(new_n987), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(KEYINPUT112), .B2(new_n980), .C1(new_n794), .C2(new_n780), .ZN(new_n989));
  INV_X1    g0789(.A(new_n201), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n780), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n982), .A2(G159), .B1(G143), .B2(new_n784), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n775), .A2(G77), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n778), .A2(new_n208), .ZN(new_n994));
  INV_X1    g0794(.A(G137), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n316), .B1(new_n763), .B2(new_n995), .C1(new_n767), .C2(new_n354), .ZN(new_n996));
  INV_X1    g0796(.A(new_n753), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n994), .B(new_n996), .C1(G58), .C2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n992), .A2(new_n993), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n989), .B1(new_n991), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n750), .B1(new_n1001), .B2(new_n798), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n967), .A2(new_n810), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n803), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n802), .B1(new_n226), .B2(new_n386), .C1(new_n241), .C2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n977), .A2(new_n1006), .ZN(G387));
  INV_X1    g0807(.A(new_n949), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n932), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(new_n694), .A3(new_n950), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n784), .A2(G322), .B1(G303), .B2(new_n781), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n979), .B2(new_n767), .C1(new_n791), .C2(new_n847), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT48), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n997), .A2(new_n502), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n794), .C2(new_n778), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT49), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n763), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(G326), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n304), .B1(new_n775), .B2(G116), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n767), .A2(new_n206), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n780), .A2(new_n208), .B1(new_n763), .B2(new_n354), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n273), .B(new_n1022), .C1(G159), .C2(new_n757), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n778), .A2(new_n386), .B1(new_n257), .B2(new_n759), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n753), .A2(new_n368), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n978), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1020), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n256), .A2(new_n206), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n695), .B1(new_n1029), .B2(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(G68), .A2(G77), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n487), .A4(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n803), .B(new_n1033), .C1(new_n238), .C2(new_n487), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n316), .A2(new_n695), .A3(new_n226), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G107), .C2(new_n226), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1038), .A2(new_n801), .A3(new_n798), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1028), .A2(new_n798), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n751), .C1(new_n684), .C2(new_n810), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1010), .B(new_n1041), .C1(new_n748), .C2(new_n1008), .ZN(G393));
  OAI22_X1  g0842(.A1(new_n767), .A2(new_n791), .B1(new_n756), .B2(new_n979), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  NAND2_X1  g0844(.A1(new_n982), .A2(G303), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n785), .A2(G116), .B1(new_n997), .B2(G283), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n316), .B1(new_n1017), .B2(G322), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1045), .A2(new_n776), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1044), .B(new_n1048), .C1(G294), .C2(new_n781), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n767), .A2(new_n764), .B1(new_n756), .B2(new_n354), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT51), .Z(new_n1051));
  NAND2_X1  g0851(.A1(new_n1017), .A2(G143), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n785), .A2(G77), .B1(new_n997), .B2(G68), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n273), .B1(new_n781), .B2(new_n256), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n843), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1051), .B(new_n1055), .C1(new_n201), .C2(new_n982), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n798), .B1(new_n1049), .B2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n802), .B1(new_n213), .B2(new_n226), .C1(new_n248), .C2(new_n1004), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n751), .A3(new_n1058), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT114), .Z(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n810), .B2(new_n939), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n944), .B2(new_n748), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT115), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n747), .B1(new_n951), .B2(new_n954), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n944), .A2(new_n950), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n1065), .A2(KEYINPUT116), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT116), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(G390));
  NOR4_X1   g0869(.A1(new_n735), .A2(new_n857), .A3(new_n664), .A4(new_n820), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n907), .B(new_n909), .C1(new_n911), .C2(new_n916), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n911), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n819), .B(new_n678), .C1(new_n706), .C2(new_n710), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1073), .A2(new_n915), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n885), .B(new_n1072), .C1(new_n1074), .C2(new_n857), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n820), .B(new_n857), .C1(new_n736), .C2(new_n742), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n916), .A2(new_n911), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1075), .C1(new_n910), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n822), .A2(new_n915), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1070), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n820), .B1(new_n736), .B2(new_n742), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n857), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n735), .A2(new_n664), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n1086), .B2(new_n819), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1081), .A2(new_n1085), .B1(new_n1088), .B2(new_n1074), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n453), .A2(G330), .A3(new_n741), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n662), .C1(new_n454), .C2(new_n919), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1077), .B(new_n1080), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n735), .A2(new_n713), .A3(new_n664), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT96), .B1(new_n741), .B2(G330), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n819), .B(new_n1084), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1086), .A2(new_n819), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n857), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1074), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n819), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1070), .B1(new_n1099), .B2(new_n857), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1081), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1091), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1080), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1102), .B(new_n1103), .C1(new_n1104), .C2(new_n1076), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1092), .A2(new_n694), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n653), .A2(new_n337), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n878), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n880), .A2(new_n872), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT38), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n890), .A2(new_n874), .B1(new_n864), .B2(new_n872), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(KEYINPUT38), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n857), .B1(new_n1073), .B2(new_n915), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1112), .A2(new_n1113), .A3(new_n911), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n908), .B1(new_n898), .B2(new_n876), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n876), .A2(new_n884), .A3(new_n908), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n916), .A2(new_n911), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1114), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1080), .B1(new_n1119), .B2(new_n1070), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n748), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n316), .B1(new_n768), .B2(G116), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n213), .B2(new_n780), .C1(new_n840), .C2(new_n763), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n754), .B(new_n1124), .C1(G283), .C2(new_n757), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n831), .B1(new_n982), .B2(G107), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n368), .C2(new_n778), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n774), .A2(new_n990), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n778), .A2(new_n764), .B1(new_n756), .B2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT54), .B(G143), .Z(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n316), .B1(new_n1132), .B2(new_n780), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1017), .A2(G125), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1128), .A2(new_n1130), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n829), .B2(new_n767), .C1(new_n995), .C2(new_n847), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n753), .A2(new_n354), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT53), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1127), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n798), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n750), .B1(new_n257), .B2(new_n827), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT117), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(new_n910), .C2(new_n800), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1106), .A2(new_n1122), .A3(new_n1145), .ZN(G378));
  AOI21_X1  g0946(.A(new_n1025), .B1(G97), .B2(new_n844), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n220), .B2(new_n756), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n282), .B1(new_n767), .B2(new_n215), .C1(new_n386), .C2(new_n780), .ZN(new_n1149));
  NOR4_X1   g0949(.A1(new_n1148), .A2(new_n304), .A3(new_n1149), .A4(new_n994), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n291), .B2(new_n774), .C1(new_n794), .C2(new_n763), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT58), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1132), .A2(new_n753), .B1(new_n829), .B2(new_n759), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n768), .A2(G128), .B1(new_n757), .B2(G125), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n995), .B2(new_n780), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(G150), .C2(new_n785), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G33), .B1(new_n1017), .B2(G124), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G41), .B1(new_n775), .B2(G159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G41), .B1(new_n304), .B2(G33), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1152), .B(new_n1161), .C1(G50), .C2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n749), .B1(new_n1163), .B2(new_n798), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n413), .A2(new_n377), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n362), .A2(new_n868), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n1167));
  XNOR2_X1  g0967(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1165), .B(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1164), .B1(new_n1171), .B2(new_n800), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n990), .B2(new_n826), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n901), .A2(new_n902), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n886), .ZN(new_n1175));
  AND4_X1   g0975(.A1(G330), .A2(new_n1174), .A3(new_n1175), .A4(new_n1171), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1171), .B1(new_n903), .B2(G330), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n918), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(G330), .A3(new_n1175), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1171), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n918), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n903), .A2(G330), .A3(new_n1171), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1173), .B1(new_n1185), .B2(new_n1121), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1091), .B1(new_n1120), .B2(new_n1102), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n694), .B1(new_n1188), .B2(KEYINPUT57), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1190), .B(new_n1187), .C1(new_n1184), .C2(new_n1178), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1186), .B1(new_n1189), .B2(new_n1191), .ZN(G375));
  NAND2_X1  g0992(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1091), .B(new_n1098), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n956), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n857), .A2(new_n799), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n798), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n785), .A2(new_n385), .B1(new_n997), .B2(G97), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n316), .B1(new_n1017), .B2(G303), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n993), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n982), .A2(G116), .B1(G107), .B2(new_n781), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n840), .B2(new_n756), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT123), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1200), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n1203), .B2(new_n1202), .C1(new_n794), .C2(new_n767), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n982), .A2(new_n1131), .B1(G132), .B2(new_n757), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n995), .B2(new_n767), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT124), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n781), .A2(G150), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(KEYINPUT124), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n778), .A2(new_n206), .B1(new_n753), .B2(new_n764), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n304), .B1(new_n1129), .B2(new_n763), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n775), .C2(G58), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1197), .B1(new_n1205), .B2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n750), .B(new_n1215), .C1(new_n208), .C2(new_n827), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT125), .Z(new_n1217));
  AOI22_X1  g1017(.A1(new_n1102), .A2(new_n1121), .B1(new_n1196), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1195), .A2(new_n1218), .ZN(G381));
  INV_X1    g1019(.A(new_n1187), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1176), .A2(new_n1177), .A3(new_n918), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1182), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1190), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1188), .A2(KEYINPUT57), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n694), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n748), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(G378), .A2(new_n1227), .A3(new_n1173), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1229), .A2(G384), .A3(G381), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1006), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n958), .B2(new_n976), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .ZN(G407));
  OAI211_X1 g1034(.A(G407), .B(G213), .C1(G343), .C2(new_n1229), .ZN(G409));
  NAND2_X1  g1035(.A1(G375), .A2(G378), .ZN(new_n1236));
  INV_X1    g1036(.A(G213), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(G343), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1188), .A2(new_n956), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1228), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT126), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1194), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1085), .A2(new_n1081), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1244), .A2(KEYINPUT60), .A3(new_n1091), .A4(new_n1098), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(new_n1193), .A3(new_n694), .A4(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1246), .A2(G384), .A3(new_n1218), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G384), .B1(new_n1246), .B2(new_n1218), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1241), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1218), .ZN(new_n1250));
  INV_X1    g1050(.A(G384), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1246), .A2(G384), .A3(new_n1218), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(KEYINPUT126), .A3(new_n1253), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1249), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1236), .A2(new_n1240), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1238), .A2(G2897), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1249), .A2(new_n1254), .A3(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1261), .A2(new_n1259), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1106), .A2(new_n1122), .A3(new_n1145), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1226), .B2(new_n1186), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1186), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1239), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1265), .A2(new_n1266), .B1(new_n1237), .B2(G343), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1260), .B(new_n1262), .C1(new_n1264), .C2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1236), .A2(new_n1240), .A3(new_n1255), .A4(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1257), .A2(new_n1258), .A3(new_n1268), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT127), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n951), .A2(new_n954), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n694), .A3(new_n1066), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT116), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1065), .A2(KEYINPUT116), .A3(new_n1066), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1063), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(G387), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(G390), .A2(new_n1232), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1272), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(G396), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1272), .B(new_n1282), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1271), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1286), .B1(new_n1288), .B2(new_n1256), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1262), .A2(new_n1260), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1256), .A2(new_n1288), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1289), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1287), .A2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(new_n1249), .A2(new_n1254), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1236), .A2(new_n1229), .A3(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1236), .A2(new_n1229), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1261), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1286), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1300), .B(new_n1301), .ZN(G402));
endmodule


