//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  INV_X1    g002(.A(G71gat), .ZN(new_n204));
  INV_X1    g003(.A(G78gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(KEYINPUT97), .B2(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n206), .A2(KEYINPUT97), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G71gat), .B(G78gat), .Z(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n209), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G231gat), .A2(G233gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n212), .A2(new_n213), .ZN(new_n219));
  XOR2_X1   g018(.A(G15gat), .B(G22gat), .Z(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G1gat), .ZN(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT16), .ZN(new_n223));
  OAI221_X1 g022(.A(new_n221), .B1(KEYINPUT95), .B2(G8gat), .C1(new_n220), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(KEYINPUT95), .A2(G8gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n218), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT98), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(G155gat), .ZN(new_n231));
  XOR2_X1   g030(.A(G183gat), .B(G211gat), .Z(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n218), .A2(new_n227), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n227), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G85gat), .A2(G92gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT7), .ZN(new_n242));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243));
  INV_X1    g042(.A(G85gat), .ZN(new_n244));
  INV_X1    g043(.A(G92gat), .ZN(new_n245));
  AOI22_X1  g044(.A1(KEYINPUT8), .A2(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G99gat), .B(G106gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT99), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n242), .A2(KEYINPUT99), .A3(new_n248), .A4(new_n246), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT10), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n253), .A2(new_n254), .A3(new_n212), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n212), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n212), .B2(new_n249), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n255), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT101), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G120gat), .B(G148gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G176gat), .B(G204gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n261), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n262), .B(new_n265), .C1(new_n266), .C2(new_n258), .ZN(new_n267));
  INV_X1    g066(.A(new_n265), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n259), .A2(new_n261), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n258), .A2(new_n266), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n267), .A2(KEYINPUT102), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT102), .B1(new_n267), .B2(new_n271), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT14), .ZN(new_n275));
  OR3_X1    g074(.A1(new_n275), .A2(G29gat), .A3(G36gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(G29gat), .B2(G36gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n278), .A2(KEYINPUT94), .ZN(new_n279));
  NAND2_X1  g078(.A1(G29gat), .A2(G36gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n280), .B(KEYINPUT92), .Z(new_n281));
  INV_X1    g080(.A(G50gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G43gat), .ZN(new_n283));
  INV_X1    g082(.A(G43gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G50gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT15), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n278), .A2(KEYINPUT94), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n279), .A2(new_n281), .A3(new_n286), .A4(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT93), .B1(new_n284), .B2(G50gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n289), .B1(G43gat), .B2(new_n282), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n284), .A2(KEYINPUT93), .A3(G50gat), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT15), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n278), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n293), .A2(new_n281), .ZN(new_n294));
  OAI22_X1  g093(.A1(new_n288), .A2(new_n292), .B1(new_n294), .B2(new_n286), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT17), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n296), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(new_n253), .ZN(new_n299));
  AND2_X1   g098(.A1(G232gat), .A2(G233gat), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n256), .A2(new_n295), .B1(KEYINPUT41), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G190gat), .B(G218gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(G134gat), .B(G162gat), .Z(new_n305));
  NOR2_X1   g104(.A1(new_n300), .A2(KEYINPUT41), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT100), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n307), .A2(KEYINPUT100), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n304), .A2(new_n308), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n240), .A2(new_n274), .A3(new_n313), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n314), .A2(KEYINPUT103), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(KEYINPUT103), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G148gat), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT80), .B1(new_n318), .B2(G141gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT80), .ZN(new_n320));
  INV_X1    g119(.A(G141gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(G148gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(G141gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT81), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT81), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G155gat), .ZN(new_n329));
  INV_X1    g128(.A(G162gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n321), .A2(G148gat), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT2), .B1(new_n338), .B2(new_n323), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n339), .A2(new_n331), .A3(new_n333), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n336), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n217), .A2(G134gat), .ZN(new_n344));
  INV_X1    g143(.A(G134gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(G127gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n343), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(G127gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n217), .A2(G134gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT72), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(G113gat), .B2(G120gat), .ZN(new_n352));
  AND2_X1   g151(.A1(G113gat), .A2(G120gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n347), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G127gat), .B(G134gat), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n356), .B(KEYINPUT72), .C1(new_n353), .C2(new_n352), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n334), .B1(new_n326), .B2(new_n327), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT3), .B1(new_n359), .B2(new_n340), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n357), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n336), .A2(new_n362), .A3(new_n341), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n340), .B1(new_n328), .B2(new_n335), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n361), .A2(new_n365), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(KEYINPUT5), .ZN(new_n370));
  INV_X1    g169(.A(new_n366), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n358), .A2(new_n359), .A3(new_n340), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n362), .B1(new_n336), .B2(new_n341), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT82), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(new_n371), .C1(new_n372), .C2(new_n373), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n375), .A2(new_n369), .A3(KEYINPUT5), .A4(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n374), .B2(KEYINPUT82), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n382), .A2(KEYINPUT83), .A3(new_n369), .A4(new_n377), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n370), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G1gat), .B(G29gat), .Z(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT6), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n370), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n357), .B(new_n355), .C1(new_n359), .C2(new_n340), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n366), .B1(new_n363), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT5), .B1(new_n394), .B2(new_n376), .ZN(new_n395));
  AOI211_X1 g194(.A(KEYINPUT82), .B(new_n366), .C1(new_n363), .C2(new_n393), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT83), .B1(new_n397), .B2(new_n369), .ZN(new_n398));
  AND4_X1   g197(.A1(KEYINPUT83), .A2(new_n382), .A3(new_n369), .A4(new_n377), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n392), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n389), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n226), .B1(new_n296), .B2(new_n295), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n406), .A2(new_n297), .B1(new_n226), .B2(new_n295), .ZN(new_n407));
  NAND2_X1  g206(.A1(G229gat), .A2(G233gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n411), .A2(KEYINPUT96), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n226), .B(new_n295), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n408), .B(KEYINPUT13), .Z(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n409), .B2(new_n410), .ZN(new_n416));
  XNOR2_X1  g215(.A(G113gat), .B(G141gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G197gat), .ZN(new_n418));
  XOR2_X1   g217(.A(KEYINPUT11), .B(G169gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n420), .B(KEYINPUT12), .Z(new_n421));
  NOR2_X1   g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n411), .A2(KEYINPUT96), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n412), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n411), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n425), .B2(new_n416), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n430), .B(KEYINPUT79), .Z(new_n431));
  NAND2_X1  g230(.A1(G183gat), .A2(G190gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT24), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT24), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(G183gat), .A3(G190gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G183gat), .ZN(new_n437));
  INV_X1    g236(.A(G190gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT68), .ZN(new_n440));
  OR3_X1    g239(.A1(KEYINPUT68), .A2(G183gat), .A3(G190gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n436), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G169gat), .A2(G176gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(KEYINPUT23), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT66), .B1(new_n444), .B2(KEYINPUT23), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT23), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n450), .B(new_n451), .C1(G169gat), .C2(G176gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n442), .A2(new_n443), .A3(new_n448), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT25), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT25), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n444), .A2(KEYINPUT23), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n456), .B(new_n443), .C1(new_n457), .C2(KEYINPUT65), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n457), .A2(KEYINPUT65), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n436), .A2(new_n439), .B1(new_n449), .B2(new_n452), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n447), .A2(KEYINPUT71), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT26), .ZN(new_n465));
  NAND2_X1  g264(.A1(KEYINPUT71), .A2(KEYINPUT26), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT67), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n464), .A2(new_n465), .B1(new_n444), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n443), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n432), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n437), .A2(KEYINPUT27), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G183gat), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT69), .A4(new_n438), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT28), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT27), .B(G183gat), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT69), .B1(new_n477), .B2(new_n438), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n471), .A2(new_n473), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT70), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT28), .A4(new_n438), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n470), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n431), .B1(new_n463), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G197gat), .ZN(new_n487));
  INV_X1    g286(.A(G204gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G197gat), .A2(G204gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT22), .ZN(new_n491));
  NAND2_X1  g290(.A1(G211gat), .A2(G218gat), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n489), .A2(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G211gat), .ZN(new_n495));
  INV_X1    g294(.A(G218gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT78), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n492), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n497), .B2(new_n492), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n494), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n501), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n493), .A3(new_n499), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n484), .B1(new_n478), .B2(new_n476), .ZN(new_n507));
  INV_X1    g306(.A(new_n470), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n454), .A2(KEYINPUT25), .B1(new_n460), .B2(new_n461), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT29), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n430), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n486), .B(new_n506), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT29), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n463), .B2(new_n485), .ZN(new_n515));
  INV_X1    g314(.A(new_n431), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(new_n510), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n512), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n513), .B1(new_n518), .B2(new_n506), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n429), .B1(new_n519), .B2(KEYINPUT37), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n512), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n431), .B2(new_n511), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n505), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n523), .A2(KEYINPUT91), .A3(new_n524), .A4(new_n513), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G8gat), .B(G36gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(G64gat), .B(G92gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n527), .B(new_n528), .Z(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n519), .B2(KEYINPUT37), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT38), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n523), .A2(new_n529), .A3(new_n513), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n524), .B1(new_n522), .B2(new_n506), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n486), .B(new_n505), .C1(new_n511), .C2(new_n512), .ZN(new_n536));
  AOI211_X1 g335(.A(KEYINPUT38), .B(new_n529), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n534), .B1(new_n526), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n402), .A2(new_n403), .A3(new_n532), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(new_n282), .ZN(new_n541));
  XOR2_X1   g340(.A(G78gat), .B(G106gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n543), .B(new_n544), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(G228gat), .ZN(new_n548));
  INV_X1    g347(.A(G233gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n506), .B1(new_n342), .B2(new_n514), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n502), .A2(new_n514), .A3(new_n504), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n367), .B1(new_n337), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n551), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n337), .ZN(new_n556));
  INV_X1    g355(.A(new_n367), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT29), .B1(new_n367), .B2(new_n337), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n558), .B(new_n550), .C1(new_n559), .C2(new_n506), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n547), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT88), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n560), .A3(new_n547), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI211_X1 g363(.A(KEYINPUT88), .B(new_n547), .C1(new_n555), .C2(new_n560), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n546), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT89), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT89), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n568), .B(new_n546), .C1(new_n564), .C2(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n561), .A2(new_n546), .ZN(new_n571));
  INV_X1    g370(.A(new_n563), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n529), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n519), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(new_n533), .A3(KEYINPUT30), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT30), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n523), .A2(new_n578), .A3(new_n529), .A4(new_n513), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n361), .A2(new_n365), .A3(new_n368), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n371), .ZN(new_n582));
  NOR4_X1   g381(.A1(new_n358), .A2(new_n359), .A3(new_n364), .A4(new_n340), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT4), .B1(new_n367), .B2(new_n362), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n366), .B1(new_n585), .B2(new_n361), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n363), .A2(new_n393), .A3(new_n366), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT39), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n582), .B(new_n390), .C1(new_n586), .C2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT40), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n577), .A2(new_n579), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT90), .B1(new_n589), .B2(new_n590), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n389), .B1(new_n586), .B2(new_n581), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n371), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT39), .A3(new_n587), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT40), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n570), .A2(new_n574), .B1(new_n600), .B2(new_n401), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n577), .A2(new_n579), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n380), .A2(new_n383), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n390), .B1(new_n603), .B2(new_n392), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n370), .B(new_n389), .C1(new_n380), .C2(new_n383), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT6), .ZN(new_n606));
  INV_X1    g405(.A(new_n403), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n602), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n573), .B1(new_n567), .B2(new_n569), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n539), .A2(new_n601), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT34), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n362), .B1(new_n463), .B2(new_n485), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n509), .A2(new_n510), .A3(new_n358), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT75), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n614), .A2(new_n615), .B1(G227gat), .B2(G233gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(KEYINPUT75), .A3(new_n613), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G227gat), .A2(G233gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT64), .Z(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT34), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT76), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT76), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n624), .A3(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT32), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n620), .A3(new_n613), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT73), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT73), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n612), .A2(new_n631), .A3(new_n620), .A4(new_n613), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n628), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT33), .B1(new_n630), .B2(new_n632), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT74), .B(G71gat), .ZN(new_n635));
  INV_X1    g434(.A(G99gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G15gat), .B(G43gat), .Z(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n633), .A2(new_n634), .A3(new_n640), .ZN(new_n641));
  AOI221_X4 g440(.A(new_n628), .B1(KEYINPUT33), .B2(new_n639), .C1(new_n630), .C2(new_n632), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n627), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n633), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n630), .A2(new_n632), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(new_n647), .A3(new_n639), .ZN(new_n648));
  INV_X1    g447(.A(new_n642), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n618), .A2(new_n626), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n643), .A2(KEYINPUT77), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT36), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT77), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n627), .B(new_n654), .C1(new_n641), .C2(new_n642), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n643), .A2(KEYINPUT36), .A3(new_n651), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n610), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n570), .A2(new_n574), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n651), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT35), .B1(new_n663), .B2(new_n608), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n609), .A2(KEYINPUT35), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n652), .A2(new_n655), .ZN(new_n666));
  INV_X1    g465(.A(new_n602), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n402), .B2(new_n403), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n428), .B1(new_n659), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n317), .A2(new_n405), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g472(.A1(new_n317), .A2(new_n671), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND4_X1  g474(.A1(new_n674), .A2(KEYINPUT42), .A3(new_n667), .A4(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(G8gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n667), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT104), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n679), .A2(new_n675), .ZN(new_n680));
  OAI221_X1 g479(.A(new_n676), .B1(new_n677), .B2(new_n679), .C1(new_n680), .C2(KEYINPUT42), .ZN(G1325gat));
  AND2_X1   g480(.A1(new_n671), .A2(new_n666), .ZN(new_n682));
  INV_X1    g481(.A(G15gat), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n317), .ZN(new_n684));
  INV_X1    g483(.A(new_n658), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n674), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n686), .B2(new_n683), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n674), .A2(new_n609), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  AOI21_X1  g489(.A(new_n313), .B1(new_n659), .B2(new_n670), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n274), .A2(new_n239), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n428), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n404), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n312), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT105), .B1(new_n610), .B2(new_n658), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n608), .A2(new_n609), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n600), .A2(new_n401), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n539), .A2(new_n660), .A3(new_n701), .ZN(new_n702));
  AND4_X1   g501(.A1(KEYINPUT105), .A2(new_n658), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT35), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n609), .A2(new_n661), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n668), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT106), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n664), .A2(new_n710), .A3(new_n669), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n698), .B1(new_n704), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n691), .A2(new_n697), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n693), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n404), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n716), .ZN(G1328gat));
  NOR3_X1   g516(.A1(new_n694), .A2(G36gat), .A3(new_n602), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT46), .ZN(new_n719));
  OAI21_X1  g518(.A(G36gat), .B1(new_n715), .B2(new_n602), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1329gat));
  OAI211_X1 g520(.A(new_n685), .B(new_n693), .C1(new_n713), .C2(new_n714), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n284), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n723), .B2(new_n722), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n692), .A2(G43gat), .A3(new_n313), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n682), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(KEYINPUT47), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n722), .A2(G43gat), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n729), .A2(KEYINPUT107), .B1(new_n682), .B2(new_n726), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n722), .A2(new_n731), .A3(G43gat), .ZN(new_n732));
  AOI211_X1 g531(.A(KEYINPUT108), .B(KEYINPUT47), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(KEYINPUT107), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n732), .A3(new_n727), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n728), .B1(new_n733), .B2(new_n738), .ZN(G1330gat));
  OAI21_X1  g538(.A(G50gat), .B1(new_n715), .B2(new_n660), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n609), .A2(new_n282), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n694), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g542(.A1(new_n704), .A2(new_n712), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n274), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n240), .A3(new_n313), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n745), .A2(new_n427), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g547(.A(new_n404), .B(KEYINPUT110), .Z(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n667), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT49), .B(G64gat), .Z(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n752), .B2(new_n754), .ZN(G1333gat));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n658), .A2(new_n204), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n748), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n748), .B2(new_n757), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n748), .A2(new_n666), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(G71gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n748), .A2(new_n609), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n274), .A2(G85gat), .A3(new_n404), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n240), .A2(new_n427), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n312), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n745), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n744), .A2(KEYINPUT51), .A3(new_n312), .A4(new_n767), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n769), .A2(KEYINPUT112), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT112), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n765), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n240), .A2(new_n274), .A3(new_n427), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n713), .ZN(new_n776));
  INV_X1    g575(.A(new_n714), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n404), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n773), .A2(new_n780), .ZN(G1336gat));
  NAND2_X1  g580(.A1(new_n769), .A2(new_n770), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n667), .A3(new_n746), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n245), .ZN(new_n784));
  NAND2_X1  g583(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n602), .A2(new_n245), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n784), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n785), .B1(new_n784), .B2(new_n788), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(G1337gat));
  NAND3_X1  g590(.A1(new_n746), .A2(new_n636), .A3(new_n666), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT114), .Z(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n771), .B2(new_n772), .ZN(new_n794));
  OAI21_X1  g593(.A(G99gat), .B1(new_n779), .B2(new_n658), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1338gat));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n779), .B2(new_n660), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n778), .A2(KEYINPUT115), .A3(new_n609), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(G106gat), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(G106gat), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n782), .A2(new_n801), .A3(new_n609), .A4(new_n746), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n802), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n801), .B1(new_n778), .B2(new_n609), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1339gat));
  NAND2_X1  g607(.A1(new_n259), .A2(new_n261), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n262), .A2(KEYINPUT54), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n265), .B1(new_n269), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(KEYINPUT55), .A3(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n813), .A2(new_n267), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n812), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n427), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n407), .A2(new_n408), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n413), .A2(new_n414), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n420), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n424), .B(new_n821), .C1(new_n272), .C2(new_n273), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n312), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n818), .A2(new_n822), .A3(KEYINPUT116), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n424), .A2(new_n821), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n817), .A2(new_n267), .A3(new_n813), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n313), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n825), .A2(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g629(.A1(new_n830), .A2(new_n240), .B1(new_n427), .B2(new_n314), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n749), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n602), .A3(new_n707), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n427), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n823), .A2(new_n824), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n313), .A3(new_n826), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n829), .A2(new_n827), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n240), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n314), .A2(new_n427), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n666), .A2(new_n660), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n405), .A2(new_n602), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(KEYINPUT117), .A3(new_n845), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n427), .A2(G113gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n835), .B1(new_n850), .B2(new_n851), .ZN(G1340gat));
  AOI21_X1  g651(.A(G120gat), .B1(new_n834), .B2(new_n746), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n746), .A2(G120gat), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n850), .B2(new_n854), .ZN(G1341gat));
  NOR2_X1   g654(.A1(new_n833), .A2(new_n239), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT118), .ZN(new_n857));
  AOI21_X1  g656(.A(G127gat), .B1(new_n856), .B2(KEYINPUT118), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n239), .A2(new_n217), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n857), .A2(new_n858), .B1(new_n850), .B2(new_n859), .ZN(G1342gat));
  NOR2_X1   g659(.A1(new_n313), .A2(new_n667), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n832), .A2(new_n345), .A3(new_n707), .A4(new_n861), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT56), .Z(new_n863));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n312), .A3(new_n849), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(G134gat), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1343gat));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n831), .A2(new_n867), .A3(new_n609), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n845), .A2(new_n658), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n823), .A2(new_n313), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n240), .B1(new_n870), .B2(new_n838), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n609), .B1(new_n871), .B2(new_n840), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n869), .B1(new_n872), .B2(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G141gat), .B1(new_n874), .B2(new_n428), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT119), .B1(new_n831), .B2(new_n749), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n685), .A2(new_n660), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n831), .A2(KEYINPUT119), .A3(new_n749), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n877), .A2(new_n602), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n427), .A2(new_n321), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT58), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n875), .B(new_n884), .C1(new_n880), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1344gat));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n869), .A2(new_n274), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n609), .A2(new_n867), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT120), .B1(new_n828), .B2(new_n313), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n814), .A2(new_n892), .A3(new_n312), .A4(new_n817), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n891), .A2(new_n827), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n870), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n239), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n315), .A2(new_n316), .A3(new_n428), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n890), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n609), .B1(new_n839), .B2(new_n840), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n889), .B(new_n898), .C1(new_n899), .C2(KEYINPUT57), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n318), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(KEYINPUT57), .ZN(new_n903));
  INV_X1    g702(.A(new_n898), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT121), .B1(new_n905), .B2(new_n889), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n887), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n874), .A2(new_n274), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(KEYINPUT59), .A3(new_n318), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n746), .A2(new_n318), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n907), .A2(new_n909), .B1(new_n880), .B2(new_n910), .ZN(G1345gat));
  NOR3_X1   g710(.A1(new_n874), .A2(new_n329), .A3(new_n239), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n879), .A2(new_n878), .ZN(new_n913));
  NOR4_X1   g712(.A1(new_n913), .A2(new_n876), .A3(new_n667), .A4(new_n239), .ZN(new_n914));
  AOI21_X1  g713(.A(G155gat), .B1(new_n914), .B2(KEYINPUT122), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n880), .B2(new_n239), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n912), .B1(new_n915), .B2(new_n917), .ZN(G1346gat));
  NAND3_X1  g717(.A1(new_n868), .A2(new_n312), .A3(new_n873), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n330), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n861), .A2(new_n330), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n913), .A2(new_n876), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G1347gat));
  OR2_X1    g726(.A1(new_n749), .A2(new_n602), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n843), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(G169gat), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n930), .A2(new_n931), .A3(new_n428), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n841), .A2(new_n405), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n663), .A2(new_n602), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n427), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n931), .B2(new_n935), .ZN(G1348gat));
  INV_X1    g735(.A(G176gat), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n930), .A2(new_n937), .A3(new_n274), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n933), .A2(new_n934), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n937), .B1(new_n939), .B2(new_n274), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(KEYINPUT125), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1349gat));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT60), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n944), .A2(KEYINPUT60), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n843), .A2(new_n240), .A3(new_n929), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G183gat), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n481), .A2(new_n483), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n933), .A2(new_n949), .A3(new_n240), .A4(new_n934), .ZN(new_n950));
  AOI211_X1 g749(.A(new_n945), .B(new_n946), .C1(new_n948), .C2(new_n950), .ZN(new_n951));
  AND4_X1   g750(.A1(new_n944), .A2(new_n948), .A3(KEYINPUT60), .A4(new_n950), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n843), .A2(new_n312), .A3(new_n929), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n954), .A2(new_n955), .A3(G190gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n954), .B2(G190gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n312), .A2(new_n438), .ZN(new_n958));
  OAI22_X1  g757(.A1(new_n956), .A2(new_n957), .B1(new_n939), .B2(new_n958), .ZN(G1351gat));
  NOR3_X1   g758(.A1(new_n685), .A2(new_n602), .A3(new_n660), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n933), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n427), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n928), .A2(new_n685), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n905), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n428), .A2(new_n487), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1352gat));
  NAND4_X1  g766(.A1(new_n933), .A2(new_n488), .A3(new_n746), .A4(new_n960), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT62), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n488), .B1(new_n965), .B2(new_n746), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n969), .A2(new_n970), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n961), .A2(new_n495), .A3(new_n240), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n903), .A2(new_n240), .A3(new_n904), .A4(new_n963), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G211gat), .ZN(new_n974));
  NOR2_X1   g773(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n974), .A2(new_n975), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  NAND3_X1  g779(.A1(new_n961), .A2(new_n496), .A3(new_n312), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n905), .A2(new_n313), .A3(new_n964), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n496), .ZN(G1355gat));
endmodule


