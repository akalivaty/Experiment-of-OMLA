//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT74), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT74), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G140), .ZN(new_n193));
  INV_X1    g007(.A(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT73), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT73), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n194), .A3(G125), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n193), .A2(KEYINPUT16), .A3(new_n196), .A4(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n190), .A2(new_n192), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n194), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(G146), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT77), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n199), .A2(new_n205), .A3(new_n202), .A4(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n189), .A2(G140), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n195), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G119), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT24), .B(G110), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT76), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n220));
  INV_X1    g034(.A(G110), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n213), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n214), .A2(new_n215), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n204), .A2(new_n206), .A3(new_n209), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n225), .A2(new_n209), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n229), .A2(KEYINPUT78), .A3(new_n204), .A4(new_n206), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n199), .A2(new_n202), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n208), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT75), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n203), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(KEYINPUT75), .A3(new_n208), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n214), .A2(new_n215), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n219), .A2(new_n220), .A3(new_n213), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(G110), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G137), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n241), .B(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n231), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n244), .B1(new_n231), .B2(new_n240), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G902), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n188), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n231), .A2(new_n240), .ZN(new_n251));
  INV_X1    g065(.A(new_n244), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n253), .A2(new_n188), .A3(new_n249), .A4(new_n245), .ZN(new_n254));
  INV_X1    g068(.A(G234), .ZN(new_n255));
  OAI21_X1  g069(.A(G217), .B1(new_n255), .B2(G902), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT72), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n187), .B1(new_n250), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n245), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT25), .B1(new_n261), .B2(G902), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n262), .A2(KEYINPUT79), .A3(new_n258), .A4(new_n254), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n258), .A2(G902), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n248), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n260), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT80), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  OR2_X1    g082(.A1(G472), .A2(G902), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n242), .A3(G210), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n270), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G137), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n276), .A2(G137), .ZN(new_n279));
  OAI21_X1  g093(.A(G131), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n281), .B1(new_n276), .B2(G137), .ZN(new_n282));
  INV_X1    g096(.A(G137), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT11), .A3(G134), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n282), .A2(new_n284), .A3(new_n285), .A4(new_n277), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n208), .A2(G143), .ZN(new_n288));
  INV_X1    g102(.A(G143), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G146), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT1), .B1(new_n289), .B2(G146), .ZN(new_n292));
  OAI21_X1  g106(.A(G128), .B1(new_n292), .B2(KEYINPUT65), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(G143), .B2(new_n208), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT65), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n291), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G143), .B(G146), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n294), .A3(G128), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n287), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n282), .A2(new_n277), .A3(new_n284), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G131), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n304), .A2(new_n286), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT0), .A2(G128), .ZN(new_n306));
  OR2_X1    g120(.A1(KEYINPUT0), .A2(G128), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n291), .A2(KEYINPUT64), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n306), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT64), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n299), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n302), .B1(new_n305), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n308), .A2(new_n311), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n304), .A2(new_n286), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(KEYINPUT67), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n301), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT66), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(G116), .B2(new_n212), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n320), .A2(KEYINPUT66), .A3(G119), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n212), .A2(G116), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT2), .B(G113), .Z(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n287), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n210), .B1(new_n295), .B2(new_n296), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n299), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n300), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n314), .A2(new_n315), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n305), .A2(new_n302), .A3(new_n312), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT67), .B1(new_n314), .B2(new_n315), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n333), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n336), .B1(new_n339), .B2(KEYINPUT30), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n275), .B(new_n327), .C1(new_n340), .C2(new_n326), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI211_X1 g157(.A(new_n301), .B(new_n325), .C1(new_n313), .C2(new_n316), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n317), .B2(new_n335), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n346), .B2(new_n325), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT31), .A3(new_n275), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g163(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n350));
  AND2_X1   g164(.A1(new_n333), .A2(new_n334), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(new_n326), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT28), .B1(new_n351), .B2(new_n326), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n275), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n269), .B1(new_n349), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT71), .B1(new_n358), .B2(KEYINPUT32), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n356), .B1(new_n343), .B2(new_n348), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT71), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n362));
  NOR4_X1   g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(new_n269), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n347), .ZN(new_n365));
  INV_X1    g179(.A(new_n275), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n353), .A2(new_n275), .A3(new_n355), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n339), .A2(new_n325), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n327), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n354), .B1(new_n372), .B2(KEYINPUT28), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n366), .A2(new_n368), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G472), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n362), .B1(new_n360), .B2(new_n269), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT70), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT70), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n380), .B(new_n362), .C1(new_n360), .C2(new_n269), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n364), .A2(new_n377), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G214), .B1(G237), .B2(G902), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT88), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n387), .A2(KEYINPUT3), .A3(G107), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  AND2_X1   g203(.A1(KEYINPUT83), .A2(G104), .ZN(new_n390));
  NOR2_X1   g204(.A1(KEYINPUT83), .A2(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n388), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n393));
  XOR2_X1   g207(.A(KEYINPUT85), .B(G101), .Z(new_n394));
  NOR2_X1   g208(.A1(new_n390), .A2(new_n391), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT84), .B1(new_n395), .B2(G107), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n397));
  NOR4_X1   g211(.A1(new_n390), .A2(new_n391), .A3(new_n397), .A4(new_n389), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n393), .B(new_n394), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  OR2_X1    g215(.A1(KEYINPUT83), .A2(G104), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT83), .A2(G104), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(G107), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n397), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n395), .A2(KEYINPUT84), .A3(G107), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n401), .B1(new_n407), .B2(new_n393), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT86), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n393), .B1(new_n396), .B2(new_n398), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G101), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT4), .A4(new_n399), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n415), .A3(G101), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n408), .A2(KEYINPUT87), .A3(new_n415), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n326), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n392), .B1(G104), .B2(new_n389), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G101), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n399), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n320), .A2(KEYINPUT5), .A3(G119), .ZN(new_n427));
  INV_X1    g241(.A(G113), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n426), .A2(new_n429), .B1(new_n324), .B2(new_n323), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G122), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT89), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n298), .A2(new_n300), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n190), .A3(new_n192), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n314), .A2(new_n200), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n242), .A2(G224), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n421), .A2(new_n431), .A3(new_n434), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT6), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n436), .B1(new_n421), .B2(new_n431), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n438), .B(new_n444), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n434), .B(KEYINPUT8), .ZN(new_n449));
  INV_X1    g263(.A(new_n431), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n425), .A2(new_n430), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n443), .A2(KEYINPUT7), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT90), .B1(new_n442), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n440), .A2(new_n456), .A3(new_n441), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n442), .A2(new_n454), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n452), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(G902), .B1(new_n460), .B2(new_n445), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n448), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n448), .B2(new_n461), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n386), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  OAI21_X1  g280(.A(G221), .B1(new_n466), .B2(G902), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT81), .Z(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G140), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n242), .A2(G227), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n439), .A2(new_n399), .A3(KEYINPUT10), .A4(new_n423), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n291), .B1(new_n295), .B2(new_n210), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n300), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n399), .A2(new_n423), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n476), .B2(KEYINPUT10), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n312), .B1(new_n418), .B2(new_n419), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n414), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n305), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n315), .B(new_n477), .C1(new_n414), .C2(new_n478), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n472), .B1(new_n479), .B2(new_n305), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n439), .B1(new_n399), .B2(new_n423), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n315), .B1(new_n484), .B2(new_n476), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(KEYINPUT12), .B(new_n315), .C1(new_n484), .C2(new_n476), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  AOI211_X1 g304(.A(G469), .B(G902), .C1(new_n482), .C2(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n472), .B(KEYINPUT82), .Z(new_n492));
  AND2_X1   g306(.A1(new_n487), .A2(new_n488), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n481), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n414), .A2(new_n478), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n315), .B1(new_n495), .B2(new_n477), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n483), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n497), .A3(G469), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(new_n249), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n469), .B1(new_n491), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G478), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G122), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G116), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n389), .B1(new_n508), .B2(KEYINPUT14), .ZN(new_n509));
  XNOR2_X1  g323(.A(G116), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT98), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n210), .B2(G143), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n289), .A2(KEYINPUT98), .A3(G128), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n210), .A2(G143), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n276), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n276), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n511), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n517), .A2(KEYINPUT99), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n510), .A2(new_n389), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n510), .A2(new_n389), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(KEYINPUT99), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n515), .A2(new_n527), .B1(new_n210), .B2(G143), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n513), .A2(KEYINPUT13), .A3(new_n514), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n276), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n520), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G217), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n466), .A2(new_n532), .A3(G953), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n520), .B(new_n533), .C1(new_n526), .C2(new_n530), .ZN(new_n536));
  AOI21_X1  g350(.A(G902), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT100), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(KEYINPUT100), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n506), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI211_X1 g356(.A(new_n249), .B(new_n242), .C1(G234), .C2(G237), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT21), .B(G898), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g359(.A1(KEYINPUT101), .A2(G952), .ZN(new_n546));
  NAND2_X1  g360(.A1(KEYINPUT101), .A2(G952), .ZN(new_n547));
  AOI21_X1  g361(.A(G953), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n255), .B2(new_n271), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n505), .B1(new_n538), .B2(new_n539), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n542), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n387), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n271), .A2(new_n242), .A3(G214), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n289), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n271), .A2(new_n242), .A3(G143), .A4(G214), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n556), .B(new_n557), .C1(new_n558), .C2(new_n285), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n196), .A2(new_n198), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n208), .B1(new_n562), .B2(new_n193), .ZN(new_n563));
  INV_X1    g377(.A(new_n209), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT91), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n193), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n196), .A2(new_n198), .ZN(new_n567));
  OAI21_X1  g381(.A(G146), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT91), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n209), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n556), .A2(new_n557), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G131), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT18), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n561), .A2(new_n565), .A3(new_n570), .A4(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n576));
  INV_X1    g390(.A(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n285), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n572), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n576), .B1(new_n579), .B2(KEYINPUT17), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n578), .A2(new_n572), .A3(KEYINPUT95), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(KEYINPUT17), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n235), .A2(new_n236), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n554), .B(new_n575), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT19), .B1(new_n566), .B2(new_n567), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT19), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n195), .A2(new_n207), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n588), .A2(new_n208), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n579), .A2(new_n594), .A3(new_n204), .A4(new_n206), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n575), .A2(new_n587), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n554), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n587), .B1(new_n575), .B2(new_n595), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n586), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT20), .ZN(new_n601));
  NOR2_X1   g415(.A1(G475), .A2(G902), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT96), .Z(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT97), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n600), .A2(new_n606), .A3(new_n601), .A4(new_n603), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n603), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT20), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n605), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n575), .B1(new_n584), .B2(new_n585), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n597), .ZN(new_n612));
  INV_X1    g426(.A(new_n586), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n249), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G475), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n552), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n465), .A2(new_n503), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n268), .A2(new_n383), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(new_n394), .Z(G3));
  NAND2_X1  g433(.A1(new_n479), .A2(new_n305), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n489), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n621), .A2(new_n492), .B1(new_n483), .B2(new_n496), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n500), .B1(new_n622), .B2(G469), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n482), .A2(new_n490), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n499), .A3(new_n249), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n468), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n349), .A2(new_n357), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n249), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n358), .B1(new_n628), .B2(G472), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n268), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n550), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n534), .A2(KEYINPUT104), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n531), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n536), .A2(KEYINPUT104), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n634), .B1(new_n531), .B2(new_n633), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT33), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n535), .A2(new_n536), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n640), .A2(KEYINPUT33), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n504), .A2(G902), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n642), .A2(new_n643), .B1(new_n504), .B2(new_n538), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n610), .B2(new_n615), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n646));
  INV_X1    g460(.A(new_n464), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n448), .A2(new_n461), .A3(new_n462), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n649), .B2(new_n386), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n646), .B(new_n386), .C1(new_n463), .C2(new_n464), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n632), .B(new_n645), .C1(new_n650), .C2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n631), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT34), .B(G104), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NAND2_X1  g470(.A1(new_n465), .A2(KEYINPUT102), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n651), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n609), .A2(new_n604), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n540), .A2(new_n541), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n505), .ZN(new_n663));
  INV_X1    g477(.A(new_n551), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n609), .A2(KEYINPUT105), .A3(new_n604), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n661), .A2(new_n615), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n658), .A2(new_n632), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n631), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT35), .B(G107), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NOR2_X1   g486(.A1(new_n252), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n251), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n264), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n260), .A2(new_n263), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n503), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n465), .A2(new_n616), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n629), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  AND2_X1   g496(.A1(new_n383), .A2(new_n678), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n684));
  OR2_X1    g498(.A1(KEYINPUT106), .A2(G900), .ZN(new_n685));
  NAND2_X1  g499(.A1(KEYINPUT106), .A2(G900), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n543), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n549), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n667), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n683), .A2(new_n684), .A3(new_n658), .A4(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n658), .A2(new_n383), .A3(new_n678), .A4(new_n690), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT107), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  XNOR2_X1  g509(.A(new_n688), .B(KEYINPUT39), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n626), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT108), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT40), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n649), .B(KEYINPUT38), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n610), .A2(new_n615), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(new_n665), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n386), .A3(new_n677), .A4(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n364), .A2(new_n382), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n347), .A2(new_n366), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n249), .B1(new_n372), .B2(new_n275), .ZN(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n699), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n289), .ZN(G45));
  AOI211_X1 g526(.A(new_n689), .B(new_n644), .C1(new_n610), .C2(new_n615), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n658), .A2(new_n383), .A3(new_n678), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  NAND2_X1  g529(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n716));
  INV_X1    g530(.A(new_n266), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n267), .ZN(new_n718));
  INV_X1    g532(.A(new_n472), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n496), .B2(new_n620), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n620), .A2(new_n719), .A3(new_n489), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n249), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(G469), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n723), .A2(new_n467), .A3(new_n625), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n383), .A2(new_n716), .A3(new_n718), .A4(new_n724), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n725), .A2(new_n653), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT41), .B(G113), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT109), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n726), .B(new_n728), .ZN(G15));
  NOR2_X1   g543(.A1(new_n669), .A2(new_n725), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n320), .ZN(G18));
  AND2_X1   g545(.A1(new_n260), .A2(new_n263), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n616), .B1(new_n732), .B2(new_n675), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n658), .A2(new_n383), .A3(new_n724), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NAND4_X1  g549(.A1(new_n723), .A2(new_n632), .A3(new_n467), .A4(new_n625), .ZN(new_n736));
  OAI21_X1  g550(.A(G472), .B1(new_n360), .B2(G902), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n373), .A2(new_n275), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n349), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n739), .B2(new_n269), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n736), .A2(new_n266), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n658), .A2(new_n741), .A3(new_n702), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  AOI21_X1  g557(.A(new_n269), .B1(new_n349), .B2(new_n738), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n628), .B2(G472), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n645), .A2(new_n745), .A3(new_n676), .A4(new_n688), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n658), .A3(new_n724), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G125), .ZN(G27));
  NAND2_X1  g562(.A1(new_n623), .A2(new_n625), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n467), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n647), .A2(new_n386), .A3(new_n648), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n644), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n701), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n689), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n268), .A2(new_n383), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n463), .A2(new_n464), .A3(new_n385), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n713), .A2(new_n757), .A3(new_n467), .A4(new_n749), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n358), .A2(KEYINPUT32), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n377), .A2(new_n759), .A3(new_n378), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n717), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT42), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n285), .ZN(G33));
  AND3_X1   g578(.A1(new_n383), .A2(new_n716), .A3(new_n718), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(KEYINPUT110), .A3(new_n690), .A4(new_n752), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n268), .A2(new_n383), .A3(new_n690), .A4(new_n752), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  NOR2_X1   g585(.A1(new_n677), .A2(new_n629), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n701), .A2(new_n644), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT43), .Z(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n772), .B(KEYINPUT44), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n757), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n779));
  OAI21_X1  g593(.A(G469), .B1(new_n622), .B2(KEYINPUT45), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(KEYINPUT45), .B2(new_n622), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n500), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n625), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n467), .B(new_n696), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n779), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(KEYINPUT113), .B(G137), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(G39));
  OAI21_X1  g607(.A(new_n467), .B1(new_n783), .B2(new_n784), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT47), .Z(new_n795));
  NAND2_X1  g609(.A1(new_n713), .A2(new_n757), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n268), .A2(new_n383), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n774), .B2(new_n549), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n773), .B(KEYINPUT43), .ZN(new_n802));
  INV_X1    g616(.A(new_n549), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(KEYINPUT120), .A3(new_n803), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n266), .B(new_n740), .C1(new_n801), .C2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n658), .A3(new_n724), .ZN(new_n806));
  INV_X1    g620(.A(new_n724), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n807), .A2(new_n549), .A3(new_n751), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n709), .A2(new_n268), .A3(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n806), .B(new_n548), .C1(new_n754), .C2(new_n809), .ZN(new_n810));
  AOI211_X1 g624(.A(new_n807), .B(new_n751), .C1(new_n801), .C2(new_n804), .ZN(new_n811));
  INV_X1    g625(.A(new_n761), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n810), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(KEYINPUT121), .A2(KEYINPUT50), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n700), .A2(new_n386), .A3(new_n807), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n805), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n805), .B2(new_n819), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n723), .A2(new_n625), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n469), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n757), .B(new_n805), .C1(new_n795), .C2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n809), .A2(new_n701), .A3(new_n753), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n677), .A2(new_n740), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n811), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n822), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(KEYINPUT122), .A3(new_n820), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n821), .B2(new_n822), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n832), .A2(new_n834), .A3(new_n826), .A4(new_n829), .ZN(new_n835));
  OAI221_X1 g649(.A(new_n816), .B1(new_n823), .B2(new_n830), .C1(new_n835), .C2(KEYINPUT51), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n714), .A2(new_n747), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n658), .A2(new_n702), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n750), .A2(new_n676), .A3(new_n689), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n708), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n692), .A2(KEYINPUT107), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n692), .A2(KEYINPUT107), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n838), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n714), .A2(new_n747), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n691), .B2(new_n693), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n841), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n746), .A2(new_n752), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n663), .A2(new_n664), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT116), .B1(new_n542), .B2(new_n551), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n689), .B1(new_n614), .B2(G475), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n666), .A2(new_n855), .A3(new_n661), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n383), .A2(new_n678), .A3(new_n857), .A4(new_n757), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n756), .A2(new_n762), .A3(new_n851), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n770), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n386), .B(new_n632), .C1(new_n463), .C2(new_n464), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n853), .A2(new_n610), .A3(new_n854), .A4(new_n615), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n862), .B1(new_n754), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n268), .A2(new_n630), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n865), .A2(new_n734), .A3(new_n742), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n669), .A2(new_n725), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n618), .A2(new_n680), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n726), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n861), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT117), .B1(new_n861), .B2(new_n869), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n859), .B1(new_n769), .B2(new_n766), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n618), .B(new_n680), .C1(new_n725), .C2(new_n653), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n865), .A2(new_n734), .A3(new_n742), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n874), .A2(new_n875), .A3(new_n730), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n850), .ZN(new_n880));
  XOR2_X1   g694(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n881));
  AOI21_X1  g695(.A(KEYINPUT119), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n883));
  INV_X1    g697(.A(new_n881), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n883), .B(new_n884), .C1(new_n879), .C2(new_n850), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n837), .B(new_n871), .C1(new_n882), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n845), .A2(new_n849), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n872), .B2(new_n878), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT53), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n884), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n886), .B1(new_n890), .B2(new_n837), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n836), .A2(new_n891), .B1(G952), .B2(G953), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n717), .A2(new_n386), .A3(new_n469), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n773), .B1(new_n893), .B2(KEYINPUT114), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(KEYINPUT114), .B2(new_n893), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT115), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n824), .B(KEYINPUT49), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n708), .A2(new_n700), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n892), .A2(new_n901), .ZN(G75));
  OAI21_X1  g716(.A(new_n871), .B1(new_n882), .B2(new_n885), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(G210), .A3(G902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n438), .B1(new_n446), .B2(new_n447), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n444), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT123), .B(KEYINPUT55), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n904), .A2(new_n905), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n909), .B1(new_n904), .B2(new_n905), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n242), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(new_n500), .B(KEYINPUT57), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n883), .B1(new_n888), .B2(new_n884), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n877), .B1(new_n873), .B2(new_n876), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(KEYINPUT119), .B(new_n881), .C1(new_n918), .C2(new_n887), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n837), .B1(new_n920), .B2(new_n871), .ZN(new_n921));
  INV_X1    g735(.A(new_n871), .ZN(new_n922));
  AOI211_X1 g736(.A(KEYINPUT54), .B(new_n922), .C1(new_n915), .C2(new_n919), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n914), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n624), .B(KEYINPUT124), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n922), .B1(new_n915), .B2(new_n919), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n249), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n781), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n912), .B1(new_n926), .B2(new_n929), .ZN(G54));
  AND2_X1   g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n903), .A2(G902), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n600), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT125), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n912), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n928), .A2(new_n936), .A3(new_n600), .A4(new_n931), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(G60));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n642), .B1(new_n891), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n642), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n886), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n942), .A2(new_n912), .A3(new_n945), .ZN(G63));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT126), .Z(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT60), .Z(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n261), .B1(new_n927), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n903), .A2(new_n674), .A3(new_n949), .ZN(new_n952));
  INV_X1    g766(.A(new_n912), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT61), .A4(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  INV_X1    g772(.A(G224), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n544), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n876), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n906), .B1(G898), .B2(new_n242), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  NAND3_X1  g777(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n340), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(G900), .A2(G953), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n839), .A2(new_n812), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n785), .A2(new_n967), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n763), .B(new_n968), .C1(new_n795), .C2(new_n797), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n791), .A2(new_n770), .A3(new_n847), .A4(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n965), .B(new_n966), .C1(new_n970), .C2(G953), .ZN(new_n971));
  INV_X1    g785(.A(new_n798), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n751), .B1(new_n754), .B2(new_n863), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n698), .A2(new_n765), .A3(new_n973), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n972), .B(new_n974), .C1(new_n789), .C2(new_n790), .ZN(new_n975));
  INV_X1    g789(.A(new_n711), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n847), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT62), .Z(new_n978));
  AOI21_X1  g792(.A(G953), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n971), .B1(new_n979), .B2(new_n965), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n242), .B1(G227), .B2(G900), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G72));
  NAND3_X1  g796(.A1(new_n975), .A2(new_n978), .A3(new_n876), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n705), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n367), .B(KEYINPUT127), .Z(new_n988));
  INV_X1    g802(.A(new_n341), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n890), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n985), .B1(new_n970), .B2(new_n869), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n365), .A2(new_n275), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n912), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n987), .A2(new_n991), .A3(new_n994), .ZN(G57));
endmodule


