

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U326 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U327 ( .A(G92GAT), .B(G218GAT), .Z(n294) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n519) );
  XNOR2_X1 U329 ( .A(n520), .B(n519), .ZN(n550) );
  XNOR2_X1 U330 ( .A(n345), .B(n344), .ZN(n512) );
  NOR2_X1 U331 ( .A1(n583), .A2(n535), .ZN(n533) );
  XOR2_X1 U332 ( .A(G197GAT), .B(G113GAT), .Z(n296) );
  XNOR2_X1 U333 ( .A(G50GAT), .B(G43GAT), .ZN(n295) );
  XNOR2_X1 U334 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U335 ( .A(n297), .B(G15GAT), .Z(n299) );
  XOR2_X1 U336 ( .A(G141GAT), .B(G22GAT), .Z(n381) );
  XNOR2_X1 U337 ( .A(G169GAT), .B(n381), .ZN(n298) );
  XNOR2_X1 U338 ( .A(n299), .B(n298), .ZN(n304) );
  XNOR2_X1 U339 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n300) );
  XNOR2_X1 U340 ( .A(n300), .B(G8GAT), .ZN(n349) );
  XOR2_X1 U341 ( .A(n349), .B(KEYINPUT66), .Z(n302) );
  NAND2_X1 U342 ( .A1(G229GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U343 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U344 ( .A(n304), .B(n303), .Z(n312) );
  XOR2_X1 U345 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U346 ( .A(G36GAT), .B(G29GAT), .ZN(n305) );
  XNOR2_X1 U347 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U348 ( .A(KEYINPUT68), .B(n307), .Z(n343) );
  XOR2_X1 U349 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n309) );
  XNOR2_X1 U350 ( .A(KEYINPUT29), .B(KEYINPUT70), .ZN(n308) );
  XNOR2_X1 U351 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U352 ( .A(n343), .B(n310), .ZN(n311) );
  XNOR2_X1 U353 ( .A(n312), .B(n311), .ZN(n576) );
  INV_X1 U354 ( .A(n576), .ZN(n478) );
  XOR2_X1 U355 ( .A(G78GAT), .B(G148GAT), .Z(n314) );
  XNOR2_X1 U356 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n313) );
  XNOR2_X1 U357 ( .A(n314), .B(n313), .ZN(n366) );
  XOR2_X1 U358 ( .A(G99GAT), .B(G71GAT), .Z(n315) );
  XOR2_X1 U359 ( .A(G120GAT), .B(n315), .Z(n392) );
  XOR2_X1 U360 ( .A(n366), .B(n392), .Z(n329) );
  XNOR2_X1 U361 ( .A(G85GAT), .B(KEYINPUT74), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n316), .B(KEYINPUT75), .ZN(n340) );
  XOR2_X1 U363 ( .A(n340), .B(KEYINPUT76), .Z(n318) );
  NAND2_X1 U364 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U366 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n320) );
  XNOR2_X1 U367 ( .A(G176GAT), .B(KEYINPUT33), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U369 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U370 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n324) );
  XNOR2_X1 U371 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n346) );
  XNOR2_X1 U373 ( .A(G204GAT), .B(G92GAT), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n325), .B(G64GAT), .ZN(n406) );
  XNOR2_X1 U375 ( .A(n346), .B(n406), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n580) );
  NAND2_X1 U378 ( .A1(n478), .A2(n580), .ZN(n466) );
  XNOR2_X1 U379 ( .A(G190GAT), .B(G99GAT), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n294), .B(n330), .ZN(n334) );
  XOR2_X1 U381 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n332) );
  XNOR2_X1 U382 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U384 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U385 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n336) );
  NAND2_X1 U386 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(n337), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U390 ( .A(n341), .B(n340), .Z(n345) );
  XOR2_X1 U391 ( .A(G43GAT), .B(G134GAT), .Z(n393) );
  XOR2_X1 U392 ( .A(G50GAT), .B(G162GAT), .Z(n380) );
  XNOR2_X1 U393 ( .A(n393), .B(n380), .ZN(n342) );
  XOR2_X1 U394 ( .A(n346), .B(G71GAT), .Z(n348) );
  XOR2_X1 U395 ( .A(G15GAT), .B(G127GAT), .Z(n400) );
  XNOR2_X1 U396 ( .A(G183GAT), .B(n400), .ZN(n347) );
  XNOR2_X1 U397 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U398 ( .A(n349), .B(KEYINPUT15), .Z(n351) );
  NAND2_X1 U399 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U400 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U401 ( .A(n353), .B(n352), .Z(n361) );
  XOR2_X1 U402 ( .A(G211GAT), .B(G78GAT), .Z(n355) );
  XNOR2_X1 U403 ( .A(G22GAT), .B(G155GAT), .ZN(n354) );
  XNOR2_X1 U404 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U405 ( .A(G64GAT), .B(KEYINPUT80), .Z(n357) );
  XNOR2_X1 U406 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U408 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U409 ( .A(n361), .B(n360), .ZN(n511) );
  INV_X1 U410 ( .A(n511), .ZN(n583) );
  NOR2_X1 U411 ( .A1(n512), .A2(n583), .ZN(n362) );
  XNOR2_X1 U412 ( .A(KEYINPUT16), .B(n362), .ZN(n451) );
  XOR2_X1 U413 ( .A(KEYINPUT2), .B(KEYINPUT92), .Z(n364) );
  XNOR2_X1 U414 ( .A(KEYINPUT91), .B(G155GAT), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U416 ( .A(KEYINPUT3), .B(n365), .Z(n434) );
  XOR2_X1 U417 ( .A(n366), .B(G204GAT), .Z(n368) );
  NAND2_X1 U418 ( .A1(G228GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U420 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n370) );
  XNOR2_X1 U421 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n369) );
  XNOR2_X1 U422 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U423 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U424 ( .A(KEYINPUT93), .B(KEYINPUT87), .Z(n374) );
  XNOR2_X1 U425 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U427 ( .A(n376), .B(n375), .ZN(n379) );
  XOR2_X1 U428 ( .A(G211GAT), .B(KEYINPUT21), .Z(n378) );
  XNOR2_X1 U429 ( .A(G197GAT), .B(G218GAT), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n378), .B(n377), .ZN(n408) );
  XOR2_X1 U431 ( .A(n379), .B(n408), .Z(n383) );
  XNOR2_X1 U432 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U433 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U434 ( .A(n434), .B(n384), .ZN(n555) );
  XOR2_X1 U435 ( .A(KEYINPUT84), .B(KEYINPUT18), .Z(n386) );
  XNOR2_X1 U436 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U438 ( .A(n387), .B(KEYINPUT19), .Z(n389) );
  XNOR2_X1 U439 ( .A(G190GAT), .B(G183GAT), .ZN(n388) );
  XNOR2_X1 U440 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U441 ( .A(G169GAT), .B(G176GAT), .Z(n390) );
  XOR2_X1 U442 ( .A(n391), .B(n390), .Z(n411) );
  XOR2_X1 U443 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U444 ( .A1(G227GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U445 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U446 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n397) );
  XNOR2_X1 U447 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n396) );
  XNOR2_X1 U448 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U449 ( .A(n399), .B(n398), .Z(n402) );
  XOR2_X1 U450 ( .A(G113GAT), .B(KEYINPUT0), .Z(n430) );
  XNOR2_X1 U451 ( .A(n400), .B(n430), .ZN(n401) );
  XNOR2_X1 U452 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U453 ( .A(n411), .B(n403), .ZN(n566) );
  XOR2_X1 U454 ( .A(G8GAT), .B(KEYINPUT100), .Z(n405) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U456 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U457 ( .A(n407), .B(n406), .Z(n410) );
  XNOR2_X1 U458 ( .A(G36GAT), .B(n408), .ZN(n409) );
  XNOR2_X1 U459 ( .A(n410), .B(n409), .ZN(n412) );
  XNOR2_X1 U460 ( .A(n412), .B(n411), .ZN(n495) );
  NAND2_X1 U461 ( .A1(n566), .A2(n495), .ZN(n413) );
  NAND2_X1 U462 ( .A1(n555), .A2(n413), .ZN(n414) );
  XOR2_X1 U463 ( .A(KEYINPUT25), .B(n414), .Z(n444) );
  XOR2_X1 U464 ( .A(KEYINPUT1), .B(KEYINPUT97), .Z(n416) );
  XNOR2_X1 U465 ( .A(KEYINPUT5), .B(KEYINPUT98), .ZN(n415) );
  XNOR2_X1 U466 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U467 ( .A(G148GAT), .B(G120GAT), .Z(n418) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(G127GAT), .ZN(n417) );
  XNOR2_X1 U469 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U470 ( .A(n420), .B(n419), .ZN(n438) );
  XOR2_X1 U471 ( .A(G57GAT), .B(KEYINPUT94), .Z(n422) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n421) );
  XNOR2_X1 U473 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U474 ( .A(KEYINPUT99), .B(KEYINPUT4), .Z(n424) );
  XNOR2_X1 U475 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U477 ( .A(n426), .B(n425), .Z(n436) );
  XOR2_X1 U478 ( .A(G85GAT), .B(G162GAT), .Z(n428) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(G134GAT), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U481 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U485 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U486 ( .A(n438), .B(n437), .ZN(n554) );
  NOR2_X1 U487 ( .A1(n555), .A2(n566), .ZN(n439) );
  XNOR2_X1 U488 ( .A(n439), .B(KEYINPUT26), .ZN(n574) );
  INV_X1 U489 ( .A(n574), .ZN(n441) );
  INV_X1 U490 ( .A(n495), .ZN(n549) );
  XOR2_X1 U491 ( .A(n549), .B(KEYINPUT101), .Z(n440) );
  XNOR2_X1 U492 ( .A(KEYINPUT27), .B(n440), .ZN(n521) );
  NOR2_X1 U493 ( .A1(n441), .A2(n521), .ZN(n442) );
  NOR2_X1 U494 ( .A1(n554), .A2(n442), .ZN(n443) );
  NAND2_X1 U495 ( .A1(n444), .A2(n443), .ZN(n449) );
  XNOR2_X1 U496 ( .A(KEYINPUT28), .B(n555), .ZN(n527) );
  XNOR2_X1 U497 ( .A(KEYINPUT86), .B(n566), .ZN(n445) );
  NOR2_X1 U498 ( .A1(n521), .A2(n445), .ZN(n446) );
  NAND2_X1 U499 ( .A1(n527), .A2(n446), .ZN(n447) );
  NAND2_X1 U500 ( .A1(n554), .A2(n447), .ZN(n448) );
  NAND2_X1 U501 ( .A1(n449), .A2(n448), .ZN(n462) );
  INV_X1 U502 ( .A(n462), .ZN(n450) );
  NAND2_X1 U503 ( .A1(n451), .A2(n450), .ZN(n479) );
  NOR2_X1 U504 ( .A1(n466), .A2(n479), .ZN(n460) );
  NAND2_X1 U505 ( .A1(n460), .A2(n554), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n453) );
  XNOR2_X1 U507 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(G1324GAT) );
  NAND2_X1 U510 ( .A1(n495), .A2(n460), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n456), .B(KEYINPUT104), .ZN(n457) );
  XNOR2_X1 U512 ( .A(G8GAT), .B(n457), .ZN(G1325GAT) );
  XOR2_X1 U513 ( .A(G15GAT), .B(KEYINPUT35), .Z(n459) );
  NAND2_X1 U514 ( .A1(n460), .A2(n566), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n459), .B(n458), .ZN(G1326GAT) );
  INV_X1 U516 ( .A(n527), .ZN(n501) );
  NAND2_X1 U517 ( .A1(n501), .A2(n460), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U519 ( .A(G29GAT), .B(KEYINPUT39), .Z(n470) );
  NOR2_X1 U520 ( .A1(n511), .A2(n462), .ZN(n464) );
  INV_X1 U521 ( .A(n512), .ZN(n568) );
  XNOR2_X1 U522 ( .A(n568), .B(KEYINPUT105), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT36), .ZN(n586) );
  NAND2_X1 U524 ( .A1(n464), .A2(n586), .ZN(n465) );
  XOR2_X1 U525 ( .A(KEYINPUT37), .B(n465), .Z(n491) );
  NOR2_X1 U526 ( .A1(n491), .A2(n466), .ZN(n468) );
  XNOR2_X1 U527 ( .A(KEYINPUT38), .B(KEYINPUT106), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n468), .B(n467), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n475), .A2(n554), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(n469), .ZN(G1328GAT) );
  NAND2_X1 U531 ( .A1(n495), .A2(n475), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n471), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n473) );
  NAND2_X1 U534 ( .A1(n475), .A2(n566), .ZN(n472) );
  XNOR2_X1 U535 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U536 ( .A(G43GAT), .B(n474), .ZN(G1330GAT) );
  NAND2_X1 U537 ( .A1(n475), .A2(n501), .ZN(n476) );
  XNOR2_X1 U538 ( .A(G50GAT), .B(n476), .ZN(G1331GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n477), .B(n580), .ZN(n558) );
  OR2_X1 U542 ( .A1(n478), .A2(n558), .ZN(n490) );
  NOR2_X1 U543 ( .A1(n490), .A2(n479), .ZN(n486) );
  NAND2_X1 U544 ( .A1(n486), .A2(n554), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U546 ( .A(G57GAT), .B(n482), .Z(G1332GAT) );
  NAND2_X1 U547 ( .A1(n495), .A2(n486), .ZN(n483) );
  XNOR2_X1 U548 ( .A(n483), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U549 ( .A(G71GAT), .B(KEYINPUT109), .Z(n485) );
  NAND2_X1 U550 ( .A1(n486), .A2(n566), .ZN(n484) );
  XNOR2_X1 U551 ( .A(n485), .B(n484), .ZN(G1334GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n488) );
  NAND2_X1 U553 ( .A1(n486), .A2(n501), .ZN(n487) );
  XNOR2_X1 U554 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U555 ( .A(G78GAT), .B(n489), .ZN(G1335GAT) );
  NOR2_X1 U556 ( .A1(n491), .A2(n490), .ZN(n492) );
  XOR2_X1 U557 ( .A(KEYINPUT111), .B(n492), .Z(n500) );
  NAND2_X1 U558 ( .A1(n554), .A2(n500), .ZN(n493) );
  XNOR2_X1 U559 ( .A(KEYINPUT112), .B(n493), .ZN(n494) );
  XNOR2_X1 U560 ( .A(G85GAT), .B(n494), .ZN(G1336GAT) );
  XOR2_X1 U561 ( .A(G92GAT), .B(KEYINPUT113), .Z(n497) );
  NAND2_X1 U562 ( .A1(n500), .A2(n495), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n497), .B(n496), .ZN(G1337GAT) );
  NAND2_X1 U564 ( .A1(n566), .A2(n500), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n498), .B(KEYINPUT114), .ZN(n499) );
  XNOR2_X1 U566 ( .A(G99GAT), .B(n499), .ZN(G1338GAT) );
  NAND2_X1 U567 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n502), .B(KEYINPUT44), .ZN(n503) );
  XNOR2_X1 U569 ( .A(G106GAT), .B(n503), .ZN(G1339GAT) );
  AND2_X1 U570 ( .A1(n576), .A2(n580), .ZN(n507) );
  NAND2_X1 U571 ( .A1(n586), .A2(n511), .ZN(n505) );
  XNOR2_X1 U572 ( .A(KEYINPUT45), .B(KEYINPUT117), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(n506) );
  AND2_X1 U574 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U575 ( .A(KEYINPUT118), .B(n508), .ZN(n518) );
  NOR2_X1 U576 ( .A1(n576), .A2(n558), .ZN(n510) );
  XNOR2_X1 U577 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n514) );
  NOR2_X1 U579 ( .A1(n512), .A2(n511), .ZN(n513) );
  NAND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(KEYINPUT116), .B(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(KEYINPUT47), .B(n516), .ZN(n517) );
  NOR2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n520) );
  INV_X1 U584 ( .A(n521), .ZN(n522) );
  NAND2_X1 U585 ( .A1(n554), .A2(n522), .ZN(n523) );
  OR2_X1 U586 ( .A1(n550), .A2(n523), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n524), .B(KEYINPUT119), .ZN(n539) );
  NAND2_X1 U588 ( .A1(n539), .A2(n566), .ZN(n526) );
  INV_X1 U589 ( .A(KEYINPUT120), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n528) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n535) );
  NOR2_X1 U592 ( .A1(n576), .A2(n535), .ZN(n529) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n529), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n558), .A2(n535), .ZN(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT121), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(n533), .Z(n534) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U600 ( .A1(n568), .A2(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT122), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n539), .A2(n574), .ZN(n546) );
  NOR2_X1 U605 ( .A1(n576), .A2(n546), .ZN(n540) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  NOR2_X1 U607 ( .A1(n546), .A2(n558), .ZN(n544) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n542) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n583), .A2(n546), .ZN(n545) );
  XOR2_X1 U613 ( .A(G155GAT), .B(n545), .Z(G1346GAT) );
  NOR2_X1 U614 ( .A1(n568), .A2(n546), .ZN(n547) );
  XOR2_X1 U615 ( .A(KEYINPUT124), .B(n547), .Z(n548) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n548), .ZN(G1347GAT) );
  INV_X1 U617 ( .A(KEYINPUT54), .ZN(n552) );
  NOR2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n575) );
  NAND2_X1 U621 ( .A1(n575), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT55), .ZN(n570) );
  NAND2_X1 U623 ( .A1(n570), .A2(n566), .ZN(n564) );
  NOR2_X1 U624 ( .A1(n576), .A2(n564), .ZN(n557) );
  XOR2_X1 U625 ( .A(G169GAT), .B(n557), .Z(G1348GAT) );
  NOR2_X1 U626 ( .A1(n558), .A2(n564), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT57), .B(KEYINPUT126), .Z(n560) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT125), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(KEYINPUT56), .B(n561), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n583), .A2(n564), .ZN(n565) );
  XOR2_X1 U633 ( .A(G183GAT), .B(n565), .Z(G1350GAT) );
  INV_X1 U634 ( .A(n566), .ZN(n567) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n573), .ZN(G1351GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n585) );
  NOR2_X1 U641 ( .A1(n576), .A2(n585), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n585), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  INV_X1 U650 ( .A(n585), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

