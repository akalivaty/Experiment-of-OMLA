//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n635, new_n638, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n453), .A2(G2106), .B1(KEYINPUT67), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n465), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(G137), .ZN(new_n477));
  NAND2_X1  g052(.A1(G101), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n471), .A2(new_n472), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n472), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(G160));
  NAND2_X1  g059(.A1(new_n474), .A2(new_n476), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND4_X1  g068(.A1(new_n474), .A2(new_n476), .A3(G138), .A4(new_n465), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n466), .A2(new_n496), .A3(G138), .A4(new_n465), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n465), .A2(G102), .A3(G2104), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n474), .A2(new_n476), .A3(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n498), .A2(new_n503), .A3(KEYINPUT71), .A4(new_n499), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G75), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n510), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n517), .A2(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n519), .A2(G62), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n521), .A2(new_n528), .ZN(G166));
  INV_X1    g104(.A(new_n512), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n531));
  OAI211_X1 g106(.A(G89), .B(new_n530), .C1(new_n519), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n525), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n513), .B2(new_n515), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  NOR4_X1   g111(.A1(new_n535), .A2(new_n536), .A3(new_n510), .A4(new_n512), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT7), .Z(new_n539));
  NOR3_X1   g114(.A1(new_n534), .A2(new_n537), .A3(new_n539), .ZN(G168));
  XNOR2_X1  g115(.A(KEYINPUT5), .B(G543), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n530), .B(new_n541), .C1(new_n519), .C2(new_n531), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n541), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n516), .ZN(new_n546));
  NOR3_X1   g121(.A1(new_n535), .A2(new_n510), .A3(new_n512), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G52), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NOR2_X1   g125(.A1(new_n514), .A2(G651), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n511), .A2(KEYINPUT72), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT6), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n553), .A2(G81), .A3(new_n530), .A4(new_n541), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n553), .A2(G43), .A3(G543), .A4(new_n530), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n522), .A2(new_n524), .A3(G56), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(new_n519), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT73), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n554), .A2(new_n555), .A3(new_n559), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  NAND2_X1  g145(.A1(new_n517), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(KEYINPUT74), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n525), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n573), .A2(new_n575), .B1(G651), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n575), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n574), .A2(KEYINPUT74), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n580), .B(new_n581), .C1(new_n571), .C2(new_n572), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n543), .A2(new_n583), .A3(G91), .ZN(new_n584));
  INV_X1    g159(.A(G91), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT75), .B1(new_n542), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n579), .A2(new_n582), .A3(new_n587), .ZN(G299));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n532), .A2(new_n533), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(new_n541), .B1(new_n547), .B2(G51), .ZN(new_n591));
  INV_X1    g166(.A(new_n539), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR4_X1   g168(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT76), .A4(new_n539), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(G286));
  INV_X1    g170(.A(G166), .ZN(G303));
  OAI21_X1  g171(.A(G651), .B1(new_n541), .B2(G74), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n543), .A2(G87), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n547), .A2(G49), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(G288));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n603));
  INV_X1    g178(.A(G86), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n542), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n517), .A2(KEYINPUT78), .A3(G86), .A4(new_n541), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G73), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G61), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n525), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n547), .A2(G48), .B1(new_n519), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(G305));
  AOI22_X1  g187(.A1(new_n541), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(new_n516), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(new_n615));
  INV_X1    g190(.A(G47), .ZN(new_n616));
  INV_X1    g191(.A(G85), .ZN(new_n617));
  OAI221_X1 g192(.A(new_n615), .B1(new_n616), .B2(new_n571), .C1(new_n617), .C2(new_n542), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT80), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n541), .A2(G66), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n511), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n547), .A2(G54), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G92), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n542), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(KEYINPUT10), .ZN(new_n629));
  AOI211_X1 g204(.A(new_n623), .B(new_n625), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n620), .B1(G868), .B2(new_n630), .ZN(G284));
  OAI21_X1  g206(.A(new_n620), .B1(G868), .B2(new_n630), .ZN(G321));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(G299), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G286), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n633), .ZN(G297));
  OAI21_X1  g211(.A(new_n634), .B1(new_n635), .B2(new_n633), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n630), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n630), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n486), .A2(G123), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT83), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n488), .A2(G135), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT82), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n650), .B(new_n651), .C1(G111), .C2(new_n465), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2096), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n465), .A2(G2104), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n485), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT13), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n660), .ZN(G156));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT15), .B(G2435), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT14), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT85), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1341), .B(G1348), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(G14), .ZN(G401));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2072), .B(G2078), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  XOR2_X1   g255(.A(new_n677), .B(KEYINPUT86), .Z(new_n681));
  OAI21_X1  g256(.A(KEYINPUT17), .B1(new_n681), .B2(new_n676), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(new_n678), .Z(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n676), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT89), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n691), .B(new_n693), .Z(new_n700));
  AOI211_X1 g275(.A(new_n697), .B(new_n699), .C1(new_n690), .C2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1986), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1991), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n703), .B(new_n706), .ZN(G229));
  NAND2_X1  g282(.A1(G299), .A2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G20), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n708), .A2(KEYINPUT23), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(KEYINPUT23), .B2(new_n710), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT102), .B(G1956), .Z(new_n713));
  XOR2_X1   g288(.A(new_n712), .B(new_n713), .Z(new_n714));
  AOI22_X1  g289(.A1(G129), .A2(new_n486), .B1(new_n488), .B2(G141), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  INV_X1    g292(.A(G105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n717), .C1(new_n718), .C2(new_n655), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT98), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G29), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT27), .B(G1996), .Z(new_n726));
  OAI211_X1 g301(.A(new_n725), .B(new_n726), .C1(G29), .C2(G32), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n725), .B1(G29), .B2(G32), .ZN(new_n728));
  INV_X1    g303(.A(new_n726), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G5), .A2(G16), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G171), .B2(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G1961), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G35), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n734), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT29), .Z(new_n737));
  INV_X1    g312(.A(G2090), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND4_X1   g314(.A1(new_n727), .A2(new_n730), .A3(new_n733), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G11), .ZN(new_n741));
  INV_X1    g316(.A(G28), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n743), .A2(new_n744), .A3(new_n734), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n741), .B(new_n745), .C1(new_n653), .C2(new_n734), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT99), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n734), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n734), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT100), .B(G2078), .Z(new_n750));
  AND2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n709), .A2(G21), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G168), .B2(new_n709), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1966), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n747), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n749), .A2(new_n750), .ZN(new_n756));
  INV_X1    g331(.A(G1961), .ZN(new_n757));
  INV_X1    g332(.A(new_n732), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n734), .A2(G33), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(new_n465), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G139), .B2(new_n488), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT25), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n734), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n757), .A2(new_n758), .B1(new_n767), .B2(G2072), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n740), .A2(new_n755), .A3(new_n756), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n767), .A2(G2072), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n737), .A2(new_n738), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT101), .ZN(new_n772));
  NAND2_X1  g347(.A1(G160), .A2(G29), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G34), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n775), .A2(new_n776), .A3(new_n734), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n769), .A2(new_n770), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n486), .A2(G128), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n488), .A2(G140), .ZN(new_n783));
  OR2_X1    g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n784), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n734), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n734), .A2(G26), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT28), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(KEYINPUT28), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT96), .B(G2067), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n709), .A2(G4), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n630), .B2(new_n709), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT94), .B(G1348), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G16), .A2(G19), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n564), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G1341), .Z(new_n802));
  NAND3_X1  g377(.A1(new_n795), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT97), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n781), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT92), .B1(G16), .B2(G23), .ZN(new_n806));
  OR3_X1    g381(.A1(KEYINPUT92), .A2(G16), .A3(G23), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n806), .B(new_n807), .C1(G288), .C2(new_n709), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT33), .B(G1976), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n709), .A2(G22), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G166), .B2(new_n709), .ZN(new_n812));
  INV_X1    g387(.A(G1971), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n709), .A2(G6), .ZN(new_n816));
  INV_X1    g391(.A(G305), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n709), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT32), .B(G1981), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT93), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n734), .A2(G25), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n486), .A2(G119), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n488), .A2(G131), .ZN(new_n827));
  NOR2_X1   g402(.A1(G95), .A2(G2105), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT90), .Z(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n734), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT35), .B(G1991), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT91), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n709), .A2(G24), .ZN(new_n837));
  INV_X1    g412(.A(G290), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n709), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(G1986), .Z(new_n840));
  NAND4_X1  g415(.A1(new_n824), .A2(new_n835), .A3(new_n836), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT36), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n836), .A2(new_n840), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n843), .A2(new_n844), .A3(new_n835), .A4(new_n824), .ZN(new_n845));
  AOI211_X1 g420(.A(new_n714), .B(new_n805), .C1(new_n842), .C2(new_n845), .ZN(G311));
  AOI21_X1  g421(.A(new_n805), .B1(new_n842), .B2(new_n845), .ZN(new_n847));
  INV_X1    g422(.A(new_n714), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(G150));
  NAND3_X1  g424(.A1(new_n522), .A2(new_n524), .A3(G67), .ZN(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n852), .A2(KEYINPUT103), .A3(new_n519), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT103), .B1(new_n852), .B2(new_n519), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND4_X1   g430(.A1(G55), .A2(new_n553), .A3(G543), .A4(new_n530), .ZN(new_n856));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  NOR4_X1   g432(.A1(new_n535), .A2(new_n525), .A3(new_n857), .A4(new_n512), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n856), .A2(new_n858), .A3(KEYINPUT104), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n517), .A2(G55), .A3(G543), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n517), .A2(G93), .A3(new_n541), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n855), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT107), .B(KEYINPUT37), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(new_n624), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(new_n638), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT39), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n561), .A2(new_n563), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n853), .A2(new_n854), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT104), .B1(new_n856), .B2(new_n858), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n861), .A2(new_n862), .A3(new_n860), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT105), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n560), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n864), .A2(new_n879), .A3(new_n564), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n871), .B(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n867), .B1(new_n884), .B2(G860), .ZN(G145));
  INV_X1    g460(.A(new_n766), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n486), .A2(G130), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n488), .A2(G142), .ZN(new_n888));
  OR2_X1    g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n723), .A2(new_n788), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n723), .A2(new_n788), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  INV_X1    g471(.A(new_n891), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n892), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n886), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n831), .B(new_n504), .Z(new_n901));
  NAND3_X1  g476(.A1(new_n895), .A2(new_n898), .A3(new_n886), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(new_n904));
  XNOR2_X1  g479(.A(G160), .B(new_n492), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n653), .B(new_n658), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  OR3_X1    g482(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g487(.A(new_n881), .B(new_n640), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n579), .A2(new_n587), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n630), .A2(new_n914), .A3(new_n582), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n869), .A2(G299), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT41), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT41), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n916), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT42), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G166), .B(G288), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n817), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n924), .A2(new_n817), .ZN(new_n927));
  OAI21_X1  g502(.A(G290), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n838), .A3(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n913), .A2(new_n919), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n932), .B(new_n933), .C1(new_n913), .C2(new_n921), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n923), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n931), .B1(new_n923), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n864), .A2(new_n633), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G295));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n937), .A2(new_n940), .A3(new_n938), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(new_n937), .B2(new_n938), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(G331));
  OAI21_X1  g518(.A(G171), .B1(new_n593), .B2(new_n594), .ZN(new_n944));
  NAND2_X1  g519(.A1(G168), .A2(G301), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n878), .A3(new_n877), .A4(new_n880), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n944), .A2(new_n945), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n881), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n919), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n921), .B1(new_n949), .B2(new_n947), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n930), .B(new_n928), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n947), .ZN(new_n955));
  INV_X1    g530(.A(new_n921), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT109), .B(new_n921), .C1(new_n949), .C2(new_n947), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n931), .B(new_n950), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(new_n909), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT111), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n953), .A2(new_n962), .A3(new_n959), .A4(new_n909), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n952), .B(new_n954), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n931), .B1(new_n965), .B2(new_n950), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n959), .A2(new_n909), .ZN(new_n967));
  OR3_X1    g542(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT43), .B1(new_n966), .B2(new_n967), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n953), .A2(new_n972), .A3(new_n959), .A4(new_n909), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g551(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n971), .C2(new_n973), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n504), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(G40), .B1(new_n480), .B2(new_n482), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n833), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n831), .B(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT112), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n723), .B(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G2067), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n787), .B(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(G290), .B(G1986), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n984), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n517), .A2(G86), .A3(new_n541), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n610), .A2(new_n519), .ZN(new_n998));
  INV_X1    g573(.A(G48), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n997), .B(new_n998), .C1(new_n571), .C2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT116), .B1(new_n1000), .B2(G1981), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n607), .A2(new_n1003), .A3(new_n611), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(G1981), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT49), .B(new_n1002), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n980), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n504), .A2(KEYINPUT113), .A3(new_n979), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G40), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n468), .B(KEYINPUT68), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n474), .A2(new_n476), .A3(G125), .ZN(new_n1016));
  OAI21_X1  g591(.A(G2105), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n477), .A2(new_n478), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n465), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(KEYINPUT69), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1014), .B1(new_n1020), .B2(new_n481), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1009), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1007), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n1001), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1008), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  INV_X1    g602(.A(G288), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1004), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1022), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n506), .A2(new_n979), .A3(new_n507), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n981), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1021), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n813), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n983), .B1(new_n1032), .B2(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n504), .A2(KEYINPUT113), .A3(new_n979), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT113), .B1(new_n504), .B2(new_n979), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1037), .B1(G2090), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G303), .A2(G8), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1045), .B(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(G8), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1021), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1028), .A2(G1976), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(G8), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1026), .A2(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1049), .A2(new_n1050), .A3(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1028), .A2(G1976), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1049), .A2(new_n1050), .A3(new_n1056), .A4(G8), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT115), .B1(new_n1060), .B2(new_n1057), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1031), .B1(new_n1048), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1026), .A2(new_n1052), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n1061), .B2(new_n1059), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n506), .A2(new_n1039), .A3(new_n979), .A4(new_n507), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1021), .A2(new_n1039), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1049), .A2(KEYINPUT117), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT117), .B1(new_n1049), .B2(new_n1070), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n738), .B(new_n1069), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1009), .B1(new_n1073), .B2(new_n1037), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1066), .B(new_n1048), .C1(new_n1047), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  INV_X1    g651(.A(G1966), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1013), .A2(KEYINPUT45), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1021), .B1(new_n1032), .B2(new_n981), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G2084), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1038), .A2(new_n1081), .A3(new_n1042), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(G168), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1085));
  AOI21_X1  g660(.A(G168), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n1087));
  OAI211_X1 g662(.A(G8), .B(new_n1083), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1076), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1075), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G2078), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1036), .B2(G2078), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1043), .A2(new_n757), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1097), .A2(G301), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1087), .B1(new_n1083), .B2(G8), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1084), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1098), .B1(new_n1102), .B2(new_n1076), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1064), .B1(new_n1090), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1105));
  INV_X1    g680(.A(G1956), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1036), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  OAI21_X1  g685(.A(G299), .B1(KEYINPUT121), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n990), .B(new_n1021), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1043), .B2(new_n798), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n630), .A3(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1033), .A2(new_n1035), .A3(new_n988), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  NAND2_X1  g698(.A1(new_n1049), .A2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1122), .A2(KEYINPUT122), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT122), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1127), .A2(new_n564), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(new_n1124), .A3(KEYINPUT122), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n564), .A3(new_n1130), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1128), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1114), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1109), .A2(KEYINPUT61), .A3(new_n1113), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n630), .B1(new_n1117), .B2(KEYINPUT60), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT124), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1117), .A2(KEYINPUT60), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1146), .B(new_n630), .C1(new_n1117), .C2(KEYINPUT60), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1145), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1121), .B1(new_n1142), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1075), .A2(new_n1102), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n983), .B(KEYINPUT125), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(new_n1034), .A3(new_n1093), .A4(new_n982), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1153), .B1(new_n1156), .B2(G171), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(G301), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(KEYINPUT126), .A3(new_n1158), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1097), .A2(G301), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1156), .A2(G171), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1153), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1152), .A2(new_n1163), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1104), .B1(new_n1151), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1009), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1048), .A2(KEYINPUT63), .A3(new_n635), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1047), .B1(new_n1044), .B2(G8), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT119), .B1(new_n1063), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1044), .A2(G8), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1047), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n1053), .A4(new_n1062), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1170), .B1(new_n1172), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1178), .A2(KEYINPUT120), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n1180));
  AOI211_X1 g755(.A(new_n1180), .B(new_n1170), .C1(new_n1172), .C2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1073), .A2(new_n1037), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1047), .B1(new_n1182), .B2(G8), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1048), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n1063), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1169), .A2(new_n635), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1179), .A2(new_n1181), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n996), .B1(new_n1168), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n984), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1190), .B1(new_n991), .B2(new_n724), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT46), .B1(new_n984), .B2(new_n988), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n984), .A2(KEYINPUT46), .A3(new_n988), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT47), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n831), .A2(new_n985), .ZN(new_n1196));
  OAI22_X1  g771(.A1(new_n992), .A2(new_n1196), .B1(G2067), .B2(new_n787), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1197), .A2(new_n984), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1190), .A2(G290), .A3(G1986), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT127), .Z(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT48), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n994), .A2(new_n984), .ZN(new_n1202));
  AOI211_X1 g777(.A(new_n1195), .B(new_n1198), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1189), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g779(.A1(G229), .A2(new_n463), .ZN(new_n1206));
  NOR2_X1   g780(.A1(G401), .A2(G227), .ZN(new_n1207));
  NAND4_X1  g781(.A1(new_n911), .A2(new_n974), .A3(new_n1206), .A4(new_n1207), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


