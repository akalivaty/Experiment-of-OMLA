

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U551 ( .A1(n680), .A2(n773), .ZN(n736) );
  OR2_X2 U552 ( .A1(n842), .A2(n695), .ZN(n699) );
  OR2_X1 U553 ( .A1(n804), .A2(n521), .ZN(n818) );
  OR2_X1 U554 ( .A1(n730), .A2(n729), .ZN(n747) );
  XNOR2_X1 U555 ( .A(KEYINPUT12), .B(KEYINPUT72), .ZN(n563) );
  AND2_X1 U556 ( .A1(n771), .A2(n770), .ZN(n519) );
  AND2_X1 U557 ( .A1(n972), .A2(n815), .ZN(n520) );
  OR2_X1 U558 ( .A1(n803), .A2(n520), .ZN(n521) );
  INV_X1 U559 ( .A(KEYINPUT100), .ZN(n766) );
  INV_X1 U560 ( .A(KEYINPUT73), .ZN(n577) );
  XNOR2_X1 U561 ( .A(n564), .B(n563), .ZN(n566) );
  NOR2_X2 U562 ( .A1(G164), .A2(G1384), .ZN(n774) );
  XOR2_X1 U563 ( .A(G543), .B(KEYINPUT0), .Z(n619) );
  NOR2_X1 U564 ( .A1(G651), .A2(G543), .ZN(n641) );
  XNOR2_X1 U565 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n542) );
  AND2_X1 U566 ( .A1(n525), .A2(G2104), .ZN(n891) );
  XNOR2_X1 U567 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U568 ( .A(n584), .B(n583), .Z(n842) );
  NOR2_X1 U569 ( .A1(n549), .A2(n548), .ZN(G160) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XOR2_X2 U571 ( .A(KEYINPUT17), .B(n522), .Z(n890) );
  NAND2_X1 U572 ( .A1(G138), .A2(n890), .ZN(n524) );
  INV_X1 U573 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U574 ( .A1(G102), .A2(n891), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n524), .A2(n523), .ZN(n529) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  NAND2_X1 U577 ( .A1(G114), .A2(n894), .ZN(n527) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n525), .ZN(n895) );
  NAND2_X1 U579 ( .A1(G126), .A2(n895), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n529), .A2(n528), .ZN(G164) );
  NOR2_X2 U582 ( .A1(G651), .A2(n619), .ZN(n642) );
  NAND2_X1 U583 ( .A1(G52), .A2(n642), .ZN(n532) );
  INV_X1 U584 ( .A(G651), .ZN(n534) );
  NOR2_X1 U585 ( .A1(G543), .A2(n534), .ZN(n530) );
  XOR2_X2 U586 ( .A(KEYINPUT1), .B(n530), .Z(n645) );
  NAND2_X1 U587 ( .A1(G64), .A2(n645), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U589 ( .A(KEYINPUT67), .B(n533), .Z(n540) );
  NAND2_X1 U590 ( .A1(G90), .A2(n641), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n534), .A2(n619), .ZN(n535) );
  XNOR2_X2 U592 ( .A(n535), .B(KEYINPUT66), .ZN(n638) );
  NAND2_X1 U593 ( .A1(G77), .A2(n638), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U595 ( .A(KEYINPUT9), .B(n538), .Z(n539) );
  NOR2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U597 ( .A(KEYINPUT68), .B(n541), .Z(G301) );
  INV_X1 U598 ( .A(G301), .ZN(G171) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U600 ( .A(G57), .ZN(G237) );
  NAND2_X1 U601 ( .A1(G101), .A2(n891), .ZN(n543) );
  NAND2_X1 U602 ( .A1(G137), .A2(n890), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G113), .A2(n894), .ZN(n547) );
  NAND2_X1 U605 ( .A1(G125), .A2(n895), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n641), .A2(G89), .ZN(n550) );
  XNOR2_X1 U608 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G76), .A2(n638), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U611 ( .A(n553), .B(KEYINPUT5), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G51), .A2(n642), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G63), .A2(n645), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U617 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(n560) );
  XNOR2_X1 U619 ( .A(KEYINPUT76), .B(n560), .ZN(G286) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U621 ( .A(n561), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U622 ( .A(G223), .B(KEYINPUT71), .ZN(n821) );
  NAND2_X1 U623 ( .A1(n821), .A2(G567), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n562), .Z(G234) );
  NAND2_X1 U625 ( .A1(G81), .A2(n641), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G68), .A2(n638), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT13), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G43), .A2(n642), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n645), .A2(G56), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(n570), .Z(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n987) );
  NAND2_X1 U634 ( .A1(n987), .A2(G860), .ZN(G153) );
  INV_X1 U635 ( .A(G868), .ZN(n661) );
  NOR2_X1 U636 ( .A1(G301), .A2(n661), .ZN(n586) );
  XNOR2_X1 U637 ( .A(KEYINPUT15), .B(KEYINPUT74), .ZN(n584) );
  INV_X1 U638 ( .A(KEYINPUT75), .ZN(n582) );
  NAND2_X1 U639 ( .A1(G92), .A2(n641), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G66), .A2(n645), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n642), .A2(G54), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G79), .A2(n638), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(n579) );
  NOR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  INV_X1 U648 ( .A(n842), .ZN(n981) );
  NOR2_X1 U649 ( .A1(n981), .A2(G868), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U651 ( .A1(n638), .A2(G78), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT70), .ZN(n594) );
  NAND2_X1 U653 ( .A1(G53), .A2(n642), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G65), .A2(n645), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G91), .A2(n641), .ZN(n590) );
  XNOR2_X1 U657 ( .A(KEYINPUT69), .B(n590), .ZN(n591) );
  NOR2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(G299) );
  NAND2_X1 U660 ( .A1(G868), .A2(G286), .ZN(n596) );
  NAND2_X1 U661 ( .A1(G299), .A2(n661), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(G297) );
  INV_X1 U663 ( .A(G860), .ZN(n611) );
  NAND2_X1 U664 ( .A1(n611), .A2(G559), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n597), .A2(n842), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U667 ( .A1(G868), .A2(n842), .ZN(n599) );
  NOR2_X1 U668 ( .A1(G559), .A2(n599), .ZN(n601) );
  AND2_X1 U669 ( .A1(n661), .A2(n987), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U671 ( .A1(G123), .A2(n895), .ZN(n602) );
  XNOR2_X1 U672 ( .A(n602), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n894), .A2(G111), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G135), .A2(n890), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G99), .A2(n891), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n924) );
  XNOR2_X1 U679 ( .A(n924), .B(G2096), .ZN(n609) );
  INV_X1 U680 ( .A(G2100), .ZN(n849) );
  NAND2_X1 U681 ( .A1(n609), .A2(n849), .ZN(G156) );
  NAND2_X1 U682 ( .A1(n842), .A2(G559), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(n987), .ZN(n658) );
  NAND2_X1 U684 ( .A1(n611), .A2(n658), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G93), .A2(n641), .ZN(n613) );
  NAND2_X1 U686 ( .A1(G80), .A2(n638), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G55), .A2(n642), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G67), .A2(n645), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n660) );
  XOR2_X1 U692 ( .A(n618), .B(n660), .Z(G145) );
  NAND2_X1 U693 ( .A1(G49), .A2(n642), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G87), .A2(n619), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n645), .A2(n622), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G651), .A2(G74), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(G288) );
  AND2_X1 U699 ( .A1(G72), .A2(n638), .ZN(n628) );
  NAND2_X1 U700 ( .A1(G85), .A2(n641), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G47), .A2(n642), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n645), .A2(G60), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(G290) );
  NAND2_X1 U706 ( .A1(G88), .A2(n641), .ZN(n632) );
  NAND2_X1 U707 ( .A1(G75), .A2(n638), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U709 ( .A1(G50), .A2(n642), .ZN(n633) );
  XNOR2_X1 U710 ( .A(KEYINPUT79), .B(n633), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n645), .A2(G62), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(G303) );
  NAND2_X1 U714 ( .A1(G73), .A2(n638), .ZN(n640) );
  XNOR2_X1 U715 ( .A(KEYINPUT78), .B(KEYINPUT2), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n650) );
  NAND2_X1 U717 ( .A1(G86), .A2(n641), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G48), .A2(n642), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U720 ( .A1(G61), .A2(n645), .ZN(n646) );
  XNOR2_X1 U721 ( .A(KEYINPUT77), .B(n646), .ZN(n647) );
  NOR2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n650), .A2(n649), .ZN(G305) );
  XNOR2_X1 U724 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n652) );
  XNOR2_X1 U725 ( .A(G288), .B(KEYINPUT19), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n660), .B(n653), .ZN(n655) );
  XOR2_X1 U728 ( .A(G290), .B(G303), .Z(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  INV_X1 U730 ( .A(G299), .ZN(n976) );
  XOR2_X1 U731 ( .A(n656), .B(n976), .Z(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(G305), .ZN(n841) );
  XOR2_X1 U733 ( .A(n841), .B(n658), .Z(n659) );
  NOR2_X1 U734 ( .A1(n661), .A2(n659), .ZN(n663) );
  AND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U736 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U743 ( .A1(G132), .A2(G82), .ZN(n668) );
  XNOR2_X1 U744 ( .A(n668), .B(KEYINPUT82), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n669), .B(KEYINPUT22), .ZN(n670) );
  NOR2_X1 U746 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U747 ( .A1(G96), .A2(n671), .ZN(n826) );
  NAND2_X1 U748 ( .A1(n826), .A2(G2106), .ZN(n675) );
  NAND2_X1 U749 ( .A1(G120), .A2(G108), .ZN(n672) );
  NOR2_X1 U750 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G69), .A2(n673), .ZN(n827) );
  NAND2_X1 U752 ( .A1(n827), .A2(G567), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n918) );
  NAND2_X1 U754 ( .A1(G661), .A2(G483), .ZN(n676) );
  XOR2_X1 U755 ( .A(KEYINPUT83), .B(n676), .Z(n677) );
  NOR2_X1 U756 ( .A1(n918), .A2(n677), .ZN(n824) );
  NAND2_X1 U757 ( .A1(n824), .A2(G36), .ZN(n678) );
  XNOR2_X1 U758 ( .A(KEYINPUT84), .B(n678), .ZN(G176) );
  INV_X1 U759 ( .A(G303), .ZN(G166) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n969) );
  INV_X1 U761 ( .A(n774), .ZN(n680) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n773) );
  NAND2_X1 U763 ( .A1(G8), .A2(n736), .ZN(n768) );
  NOR2_X1 U764 ( .A1(G288), .A2(G1976), .ZN(n681) );
  XNOR2_X1 U765 ( .A(n681), .B(KEYINPUT97), .ZN(n751) );
  NOR2_X1 U766 ( .A1(n768), .A2(n751), .ZN(n682) );
  NAND2_X1 U767 ( .A1(KEYINPUT33), .A2(n682), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n969), .A2(n683), .ZN(n758) );
  NAND2_X1 U769 ( .A1(G1341), .A2(n736), .ZN(n688) );
  INV_X1 U770 ( .A(G1996), .ZN(n684) );
  NOR2_X1 U771 ( .A1(n773), .A2(n684), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n774), .A2(n685), .ZN(n686) );
  XNOR2_X1 U773 ( .A(n686), .B(KEYINPUT26), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U775 ( .A(n689), .B(KEYINPUT93), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n690), .A2(n987), .ZN(n692) );
  INV_X1 U777 ( .A(KEYINPUT64), .ZN(n691) );
  XNOR2_X1 U778 ( .A(n692), .B(n691), .ZN(n695) );
  INV_X1 U779 ( .A(n736), .ZN(n715) );
  NOR2_X1 U780 ( .A1(n715), .A2(G1348), .ZN(n694) );
  NOR2_X1 U781 ( .A1(G2067), .A2(n736), .ZN(n693) );
  NOR2_X1 U782 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n842), .A2(n695), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U786 ( .A(n700), .B(KEYINPUT94), .ZN(n707) );
  NAND2_X1 U787 ( .A1(G1956), .A2(n736), .ZN(n701) );
  XNOR2_X1 U788 ( .A(KEYINPUT91), .B(n701), .ZN(n705) );
  XOR2_X1 U789 ( .A(KEYINPUT27), .B(KEYINPUT90), .Z(n703) );
  NAND2_X1 U790 ( .A1(n715), .A2(G2072), .ZN(n702) );
  XOR2_X1 U791 ( .A(n703), .B(n702), .Z(n704) );
  NOR2_X1 U792 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U793 ( .A1(n708), .A2(n976), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n707), .A2(n706), .ZN(n712) );
  NOR2_X1 U795 ( .A1(n708), .A2(n976), .ZN(n710) );
  XOR2_X1 U796 ( .A(KEYINPUT92), .B(KEYINPUT28), .Z(n709) );
  XNOR2_X1 U797 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U799 ( .A(KEYINPUT29), .B(KEYINPUT95), .ZN(n713) );
  XNOR2_X1 U800 ( .A(n714), .B(n713), .ZN(n733) );
  OR2_X1 U801 ( .A1(n715), .A2(G1961), .ZN(n717) );
  XNOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .ZN(n949) );
  NAND2_X1 U803 ( .A1(n715), .A2(n949), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n717), .A2(n716), .ZN(n721) );
  NAND2_X1 U805 ( .A1(n721), .A2(G171), .ZN(n731) );
  NAND2_X1 U806 ( .A1(n733), .A2(n731), .ZN(n725) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n768), .ZN(n727) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n736), .ZN(n726) );
  NOR2_X1 U809 ( .A1(n727), .A2(n726), .ZN(n718) );
  NAND2_X1 U810 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U811 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U812 ( .A1(G168), .A2(n720), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n721), .A2(G171), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U815 ( .A(KEYINPUT31), .B(n724), .Z(n734) );
  AND2_X1 U816 ( .A1(n725), .A2(n734), .ZN(n730) );
  AND2_X1 U817 ( .A1(G8), .A2(n726), .ZN(n728) );
  OR2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U819 ( .A1(n731), .A2(G286), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n743) );
  INV_X1 U821 ( .A(G286), .ZN(n735) );
  OR2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n741) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n768), .ZN(n738) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n739), .A2(G303), .ZN(n740) );
  AND2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U828 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n744), .A2(G8), .ZN(n745) );
  XNOR2_X1 U830 ( .A(n745), .B(KEYINPUT32), .ZN(n746) );
  NAND2_X1 U831 ( .A1(n747), .A2(n746), .ZN(n749) );
  INV_X1 U832 ( .A(KEYINPUT96), .ZN(n748) );
  XNOR2_X1 U833 ( .A(n749), .B(n748), .ZN(n765) );
  OR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NAND2_X1 U835 ( .A1(n751), .A2(n750), .ZN(n973) );
  NOR2_X1 U836 ( .A1(n765), .A2(n973), .ZN(n755) );
  NAND2_X1 U837 ( .A1(G288), .A2(G1976), .ZN(n752) );
  XNOR2_X1 U838 ( .A(n752), .B(KEYINPUT98), .ZN(n975) );
  INV_X1 U839 ( .A(n975), .ZN(n753) );
  OR2_X1 U840 ( .A1(n753), .A2(n768), .ZN(n754) );
  NOR2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U842 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U843 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U844 ( .A(n759), .B(KEYINPUT99), .ZN(n772) );
  NOR2_X1 U845 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XOR2_X1 U846 ( .A(n760), .B(KEYINPUT24), .Z(n761) );
  NOR2_X1 U847 ( .A1(n768), .A2(n761), .ZN(n762) );
  XNOR2_X1 U848 ( .A(n762), .B(KEYINPUT89), .ZN(n771) );
  NAND2_X1 U849 ( .A1(G166), .A2(G8), .ZN(n763) );
  NOR2_X1 U850 ( .A1(G2090), .A2(n763), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n767) );
  XNOR2_X1 U852 ( .A(n767), .B(n766), .ZN(n769) );
  NAND2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n770) );
  AND2_X1 U854 ( .A1(n772), .A2(n519), .ZN(n804) );
  NOR2_X1 U855 ( .A1(n774), .A2(n773), .ZN(n815) );
  NAND2_X1 U856 ( .A1(G140), .A2(n890), .ZN(n776) );
  NAND2_X1 U857 ( .A1(G104), .A2(n891), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n777), .ZN(n782) );
  NAND2_X1 U860 ( .A1(G116), .A2(n894), .ZN(n779) );
  NAND2_X1 U861 ( .A1(G128), .A2(n895), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U863 ( .A(KEYINPUT35), .B(n780), .Z(n781) );
  NOR2_X1 U864 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U865 ( .A(KEYINPUT36), .B(n783), .ZN(n908) );
  XNOR2_X1 U866 ( .A(G2067), .B(KEYINPUT37), .ZN(n813) );
  NOR2_X1 U867 ( .A1(n908), .A2(n813), .ZN(n930) );
  NAND2_X1 U868 ( .A1(n815), .A2(n930), .ZN(n811) );
  NAND2_X1 U869 ( .A1(n890), .A2(G141), .ZN(n784) );
  XNOR2_X1 U870 ( .A(KEYINPUT88), .B(n784), .ZN(n792) );
  NAND2_X1 U871 ( .A1(G117), .A2(n894), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G129), .A2(n895), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n891), .A2(G105), .ZN(n787) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U877 ( .A(KEYINPUT87), .B(n790), .Z(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n903) );
  AND2_X1 U879 ( .A1(n903), .A2(G1996), .ZN(n801) );
  XOR2_X1 U880 ( .A(KEYINPUT86), .B(G1991), .Z(n946) );
  NAND2_X1 U881 ( .A1(n894), .A2(G107), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G131), .A2(n890), .ZN(n793) );
  XOR2_X1 U883 ( .A(KEYINPUT85), .B(n793), .Z(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G95), .A2(n891), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G119), .A2(n895), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n902) );
  NOR2_X1 U889 ( .A1(n946), .A2(n902), .ZN(n800) );
  NOR2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n927) );
  INV_X1 U891 ( .A(n927), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n802), .A2(n815), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n811), .A2(n805), .ZN(n803) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n972) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n903), .ZN(n934) );
  INV_X1 U896 ( .A(n805), .ZN(n808) );
  AND2_X1 U897 ( .A1(n946), .A2(n902), .ZN(n925) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U899 ( .A1(n925), .A2(n806), .ZN(n807) );
  NOR2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U901 ( .A1(n934), .A2(n809), .ZN(n810) );
  XNOR2_X1 U902 ( .A(KEYINPUT39), .B(n810), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n908), .A2(n813), .ZN(n932) );
  NAND2_X1 U905 ( .A1(n814), .A2(n932), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n820) );
  XOR2_X1 U908 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n819) );
  XNOR2_X1 U909 ( .A(n820), .B(n819), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U912 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n823) );
  XNOR2_X1 U914 ( .A(KEYINPUT106), .B(n823), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(n824), .ZN(G188) );
  XOR2_X1 U916 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U918 ( .A(G132), .ZN(G219) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G82), .ZN(G220) );
  NOR2_X1 U921 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U923 ( .A(G1341), .B(G1348), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n828), .B(G2427), .ZN(n838) );
  XOR2_X1 U925 ( .A(G2446), .B(G2430), .Z(n830) );
  XNOR2_X1 U926 ( .A(G2454), .B(G2451), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT102), .B(G2435), .Z(n832) );
  XNOR2_X1 U929 ( .A(KEYINPUT103), .B(G2438), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U931 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U932 ( .A(KEYINPUT104), .B(G2443), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n839), .A2(G14), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n840), .B(KEYINPUT105), .ZN(G401) );
  XNOR2_X1 U937 ( .A(G286), .B(n841), .ZN(n844) );
  XOR2_X1 U938 ( .A(n842), .B(n987), .Z(n843) );
  XNOR2_X1 U939 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U940 ( .A(n845), .B(G171), .Z(n846) );
  NOR2_X1 U941 ( .A1(G37), .A2(n846), .ZN(G397) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2090), .Z(n848) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(n850) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n852) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U947 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U949 ( .A(G2678), .B(KEYINPUT107), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U951 ( .A(n856), .B(n855), .Z(G227) );
  XOR2_X1 U952 ( .A(G2474), .B(G1981), .Z(n858) );
  XNOR2_X1 U953 ( .A(G1966), .B(G1961), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U955 ( .A(n859), .B(KEYINPUT108), .Z(n861) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U958 ( .A(G1976), .B(G1971), .Z(n863) );
  XNOR2_X1 U959 ( .A(G1986), .B(G1956), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U961 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U962 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G136), .A2(n890), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n868), .B(KEYINPUT110), .ZN(n874) );
  NAND2_X1 U966 ( .A1(G100), .A2(n891), .ZN(n869) );
  XOR2_X1 U967 ( .A(KEYINPUT112), .B(n869), .Z(n872) );
  NAND2_X1 U968 ( .A1(n895), .A2(G124), .ZN(n870) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n870), .Z(n871) );
  NOR2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n877) );
  NAND2_X1 U972 ( .A1(G112), .A2(n894), .ZN(n875) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n875), .ZN(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G142), .A2(n890), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G106), .A2(n891), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n880), .B(KEYINPUT45), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G118), .A2(n894), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G130), .A2(n895), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(KEYINPUT113), .B(n883), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n886), .B(n924), .ZN(n887) );
  XNOR2_X1 U985 ( .A(G160), .B(n887), .ZN(n907) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n889) );
  XNOR2_X1 U987 ( .A(G164), .B(G162), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n901) );
  NAND2_X1 U989 ( .A1(G139), .A2(n890), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G103), .A2(n891), .ZN(n892) );
  NAND2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U992 ( .A1(G115), .A2(n894), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G127), .A2(n895), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n919) );
  XOR2_X1 U997 ( .A(n901), .B(n919), .Z(n905) );
  XOR2_X1 U998 ( .A(n903), .B(n902), .Z(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1001 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n910), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(KEYINPUT114), .B(n911), .ZN(G395) );
  NOR2_X1 U1004 ( .A1(G401), .A2(n918), .ZN(n915) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n913), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(n916), .A2(G395), .ZN(n917) );
  XOR2_X1 U1010 ( .A(n917), .B(KEYINPUT115), .Z(G308) );
  INV_X1 U1011 ( .A(G308), .ZN(G225) );
  INV_X1 U1012 ( .A(n918), .ZN(G319) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1015 ( .A(G164), .B(G2078), .ZN(n922) );
  XOR2_X1 U1016 ( .A(G2072), .B(n919), .Z(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT117), .B(n920), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(n923), .B(KEYINPUT50), .ZN(n941) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1021 ( .A1(n927), .A2(n926), .ZN(n929) );
  XOR2_X1 U1022 ( .A(G160), .B(G2084), .Z(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n939) );
  INV_X1 U1024 ( .A(n930), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n937) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1028 ( .A(n935), .B(KEYINPUT51), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1031 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n942), .ZN(n944) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1035 ( .A1(n945), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n961) );
  XNOR2_X1 U1037 ( .A(n946), .B(G25), .ZN(n947) );
  NAND2_X1 U1038 ( .A1(n947), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(n948), .B(KEYINPUT118), .ZN(n958) );
  XNOR2_X1 U1040 ( .A(n949), .B(G27), .ZN(n951) );
  XOR2_X1 U1041 ( .A(G1996), .B(G32), .Z(n950) );
  NAND2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n952), .ZN(n956) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n959), .ZN(n960) );
  NOR2_X1 U1050 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n962) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n962), .ZN(n963) );
  NAND2_X1 U1053 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1054 ( .A(KEYINPUT55), .B(n965), .Z(n967) );
  INV_X1 U1055 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n968), .ZN(n1023) );
  INV_X1 U1058 ( .A(G16), .ZN(n1019) );
  XOR2_X1 U1059 ( .A(n1019), .B(KEYINPUT56), .Z(n993) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n971), .B(KEYINPUT57), .ZN(n991) );
  NOR2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n980) );
  NAND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1066 ( .A(G1956), .B(n976), .Z(n977) );
  NOR2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n985) );
  XOR2_X1 U1069 ( .A(G301), .B(G1961), .Z(n983) );
  XOR2_X1 U1070 ( .A(n981), .B(G1348), .Z(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1073 ( .A(KEYINPUT120), .B(n986), .Z(n989) );
  XOR2_X1 U1074 ( .A(n987), .B(G1341), .Z(n988) );
  NOR2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1077 ( .A1(n993), .A2(n992), .ZN(n1021) );
  XNOR2_X1 U1078 ( .A(KEYINPUT123), .B(G1966), .ZN(n994) );
  XNOR2_X1 U1079 ( .A(n994), .B(G21), .ZN(n1014) );
  XOR2_X1 U1080 ( .A(G1956), .B(G20), .Z(n997) );
  XNOR2_X1 U1081 ( .A(G19), .B(KEYINPUT121), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n995), .B(G1341), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G6), .B(G1981), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(KEYINPUT122), .B(n1000), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1001), .B(G4), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(n1004), .B(KEYINPUT60), .ZN(n1012) );
  XNOR2_X1 U1091 ( .A(G1986), .B(G24), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(G1971), .B(KEYINPUT124), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G22), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(G5), .B(G1961), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1105 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1106 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1107 ( .A(n1026), .B(KEYINPUT62), .ZN(n1027) );
  XNOR2_X1 U1108 ( .A(KEYINPUT125), .B(n1027), .ZN(G311) );
  XOR2_X1 U1109 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

