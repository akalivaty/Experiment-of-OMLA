//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(KEYINPUT3), .A3(G107), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT79), .A2(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT79), .A2(G104), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G107), .A3(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(G107), .B1(new_n192), .B2(new_n193), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n191), .B(new_n194), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT4), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G101), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G116), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G113), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G113), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n208), .ZN(new_n210));
  XNOR2_X1  g024(.A(G116), .B(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n212), .A3(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n212), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n199), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n191), .B1(new_n195), .B2(new_n196), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n194), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT80), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G107), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT79), .A2(G104), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT79), .A2(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n190), .B1(new_n225), .B2(KEYINPUT3), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n223), .A2(new_n224), .ZN(new_n228));
  AOI21_X1  g042(.A(G101), .B1(new_n228), .B2(G107), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n198), .B1(new_n197), .B2(G101), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n217), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n189), .A2(G107), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n219), .B1(new_n225), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n211), .A2(KEYINPUT5), .ZN(new_n236));
  OAI21_X1  g050(.A(G113), .B1(new_n201), .B2(KEYINPUT5), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n212), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI211_X1 g052(.A(new_n235), .B(new_n238), .C1(new_n221), .C2(new_n230), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n188), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n235), .B1(new_n221), .B2(new_n230), .ZN(new_n241));
  INV_X1    g055(.A(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n227), .B1(new_n226), .B2(new_n229), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n232), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n243), .B(new_n187), .C1(new_n247), .C2(new_n217), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n248), .A3(KEYINPUT6), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT64), .A2(G146), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(G143), .A3(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n256), .A2(G146), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT64), .B(G146), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(new_n256), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT0), .B(G128), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G125), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  INV_X1    g079(.A(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n254), .A2(new_n257), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n254), .B2(KEYINPUT1), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n265), .B(new_n268), .C1(new_n269), .C2(new_n261), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G224), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n273), .B(KEYINPUT82), .Z(new_n274));
  XNOR2_X1  g088(.A(new_n271), .B(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(new_n188), .C1(new_n233), .C2(new_n239), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n249), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n187), .B(KEYINPUT8), .Z(new_n279));
  INV_X1    g093(.A(new_n235), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n244), .B2(new_n245), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n238), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n282), .B2(new_n243), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n270), .A4(new_n273), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT83), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n279), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n241), .A2(new_n242), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(new_n239), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT83), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n285), .A2(new_n286), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(new_n294), .A3(new_n248), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n278), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n278), .A2(new_n295), .A3(new_n296), .A4(new_n298), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G113), .B(G122), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(new_n189), .ZN(new_n304));
  XNOR2_X1  g118(.A(G125), .B(G140), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n252), .A3(new_n253), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n251), .B2(new_n305), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n272), .A3(G214), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n256), .ZN(new_n310));
  NOR2_X1   g124(.A1(G237), .A2(G953), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(G143), .A3(G214), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT18), .ZN(new_n314));
  INV_X1    g128(.A(G131), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n310), .A2(new_n312), .B1(KEYINPUT18), .B2(G131), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n307), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n305), .B2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n265), .A2(G140), .ZN(new_n323));
  AND4_X1   g137(.A1(new_n319), .A2(new_n322), .A3(new_n323), .A4(KEYINPUT16), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT74), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT16), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n321), .A4(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n326), .A3(G146), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT16), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n322), .A2(new_n323), .A3(new_n319), .A4(KEYINPUT16), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n331), .A2(new_n334), .A3(G146), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT75), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n331), .A2(new_n334), .A3(new_n335), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n251), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n332), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n312), .ZN(new_n341));
  AOI21_X1  g155(.A(G143), .B1(new_n311), .B2(G214), .ZN(new_n342));
  OAI21_X1  g156(.A(G131), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT17), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n310), .A2(new_n315), .A3(new_n312), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n313), .A2(KEYINPUT17), .A3(G131), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n304), .B(new_n318), .C1(new_n340), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n345), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n305), .B(KEYINPUT19), .Z(new_n351));
  OAI211_X1 g165(.A(new_n336), .B(new_n350), .C1(new_n351), .C2(new_n260), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n318), .ZN(new_n353));
  INV_X1    g167(.A(new_n304), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G475), .A2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT20), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n360), .A3(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n349), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n346), .A2(new_n347), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(new_n332), .A3(new_n339), .A4(new_n337), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n304), .B1(new_n365), .B2(new_n318), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT84), .B(new_n296), .C1(new_n363), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G475), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n318), .B1(new_n340), .B2(new_n348), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n354), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n370), .B2(new_n349), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(KEYINPUT84), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n362), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n256), .A2(KEYINPUT13), .A3(G128), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n266), .A2(G143), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n266), .A2(G143), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT13), .ZN(new_n379));
  OAI221_X1 g193(.A(G134), .B1(new_n374), .B2(new_n375), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n256), .A2(G128), .ZN(new_n381));
  INV_X1    g195(.A(G134), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G122), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G116), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n202), .A2(G122), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G107), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n386), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n222), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n380), .A2(new_n383), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n256), .A2(G128), .ZN(new_n391));
  OAI21_X1  g205(.A(G134), .B1(new_n378), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n383), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(KEYINPUT86), .A3(new_n383), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n222), .B1(new_n385), .B2(KEYINPUT14), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n388), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n397), .A2(new_n388), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n395), .A2(new_n396), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT9), .B(G234), .ZN(new_n401));
  INV_X1    g215(.A(G217), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n401), .A2(new_n402), .A3(G953), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n390), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n390), .B2(new_n400), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n405), .A2(new_n406), .A3(G902), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT15), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n407), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n373), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(G234), .A2(G237), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n413), .A2(G952), .A3(new_n272), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT87), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n413), .A2(G902), .A3(G953), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G214), .B1(G237), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n302), .A2(new_n412), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n272), .A2(G227), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n427));
  AND2_X1   g241(.A1(KEYINPUT64), .A2(G146), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT64), .A2(G146), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n256), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n259), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n262), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT66), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT66), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n258), .B(new_n434), .C1(new_n261), .C2(new_n262), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n433), .A2(new_n199), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n246), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n254), .A2(new_n257), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n266), .B1(new_n431), .B2(KEYINPUT1), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n268), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n280), .B(new_n440), .C1(new_n244), .C2(new_n245), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n268), .B1(new_n269), .B2(new_n261), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n444), .A2(KEYINPUT10), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n241), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n437), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT11), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n382), .B2(G137), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n382), .A2(G137), .ZN(new_n450));
  INV_X1    g264(.A(G137), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT11), .A3(G134), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G131), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n452), .A3(new_n315), .A4(new_n450), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n456), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n436), .A2(new_n246), .B1(new_n241), .B2(new_n445), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(new_n443), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n426), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n441), .B1(new_n241), .B2(new_n444), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n456), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT12), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n458), .A3(new_n443), .ZN(new_n465));
  INV_X1    g279(.A(new_n426), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n462), .A2(new_n467), .A3(new_n456), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G469), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n296), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n296), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n426), .ZN(new_n476));
  INV_X1    g290(.A(new_n460), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n465), .A3(new_n466), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(G469), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n472), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G221), .B1(new_n401), .B2(G902), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n423), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n402), .B1(G234), .B2(new_n296), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT77), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT22), .B(G137), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n266), .A2(G119), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n200), .A2(G128), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT24), .B(G110), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT71), .B1(new_n200), .B2(G128), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT23), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT71), .B(new_n496), .C1(new_n200), .C2(G128), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n490), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G110), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT72), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n501), .A3(G110), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n493), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n340), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G110), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n495), .A2(new_n505), .A3(new_n490), .A4(new_n497), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n491), .A2(new_n492), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n336), .A2(new_n508), .A3(new_n306), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT76), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n512));
  AOI211_X1 g326(.A(new_n512), .B(new_n509), .C1(new_n340), .C2(new_n503), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n488), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n509), .B1(new_n340), .B2(new_n503), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n515), .A2(new_n488), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT25), .B1(new_n517), .B2(new_n296), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n519));
  AOI211_X1 g333(.A(new_n519), .B(G902), .C1(new_n514), .C2(new_n516), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n484), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT78), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT78), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(new_n484), .C1(new_n518), .C2(new_n520), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n484), .A2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n433), .A2(new_n456), .A3(new_n435), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n216), .A2(new_n213), .ZN(new_n529));
  INV_X1    g343(.A(new_n450), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n382), .A2(G137), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n532), .A2(new_n455), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n444), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT28), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n311), .A2(G210), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT27), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n545), .A2(KEYINPUT29), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT69), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n528), .A2(new_n534), .ZN(new_n548));
  INV_X1    g362(.A(new_n529), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n535), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n547), .B1(new_n551), .B2(KEYINPUT28), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n529), .B1(new_n528), .B2(new_n534), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n547), .B(KEYINPUT28), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n541), .B(new_n546), .C1(new_n552), .C2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT28), .B1(new_n553), .B2(new_n554), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT69), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n555), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n562), .A2(KEYINPUT70), .A3(new_n541), .A4(new_n546), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT30), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n444), .A2(new_n533), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n458), .A2(new_n263), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n528), .A2(KEYINPUT30), .A3(new_n534), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n549), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n535), .ZN(new_n570));
  INV_X1    g384(.A(new_n545), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT29), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n458), .A2(new_n263), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n529), .B1(new_n573), .B2(new_n534), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT28), .B1(new_n553), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n540), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n545), .B(KEYINPUT67), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n538), .A4(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(G902), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n559), .A2(new_n563), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G472), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n569), .A2(new_n535), .A3(new_n545), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT31), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n569), .A2(KEYINPUT31), .A3(new_n535), .A4(new_n545), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n576), .A3(new_n538), .ZN(new_n586));
  INV_X1    g400(.A(new_n577), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n584), .A2(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(G472), .A2(G902), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT32), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n584), .A2(new_n585), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n586), .A2(new_n587), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT32), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n589), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n581), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n483), .A2(new_n527), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NOR2_X1   g414(.A1(new_n588), .A2(G902), .ZN(new_n601));
  INV_X1    g415(.A(G472), .ZN(new_n602));
  OAI22_X1  g416(.A1(new_n601), .A2(new_n602), .B1(new_n588), .B2(new_n590), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n482), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n527), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n419), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT92), .B(G478), .ZN(new_n608));
  OR3_X1    g422(.A1(new_n407), .A2(KEYINPUT93), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT93), .B1(new_n407), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT90), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n390), .A2(new_n400), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n403), .B1(new_n613), .B2(KEYINPUT91), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT90), .B1(new_n403), .B2(KEYINPUT91), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n390), .B2(new_n400), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT33), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n408), .A2(G902), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT33), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT89), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR4_X1   g435(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT89), .A4(KEYINPUT33), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n617), .B(new_n618), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n611), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n373), .A2(new_n607), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n300), .A2(KEYINPUT88), .A3(new_n301), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT88), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n297), .A2(new_n627), .A3(new_n299), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n625), .A2(new_n626), .A3(new_n420), .A4(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT94), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n628), .A2(new_n420), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n632), .A2(KEYINPUT94), .A3(new_n626), .A4(new_n625), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n606), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND3_X1  g451(.A1(new_n626), .A2(new_n420), .A3(new_n628), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n411), .B(new_n362), .C1(new_n372), .C2(new_n368), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n638), .A2(new_n419), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n606), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR2_X1   g457(.A1(new_n423), .A2(new_n603), .ZN(new_n644));
  INV_X1    g458(.A(new_n481), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n461), .B2(new_n469), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n473), .B1(new_n646), .B2(new_n471), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n645), .B1(new_n647), .B2(new_n479), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n511), .A2(new_n513), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n488), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n525), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n522), .A2(new_n524), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n644), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  AND2_X1   g470(.A1(new_n653), .A2(new_n648), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n414), .B1(new_n418), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n639), .A2(new_n659), .ZN(new_n660));
  AOI22_X1  g474(.A1(G472), .A2(new_n580), .B1(new_n591), .B2(new_n596), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n638), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XOR2_X1   g478(.A(new_n659), .B(KEYINPUT39), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n648), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT40), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n302), .B(KEYINPUT38), .ZN(new_n668));
  INV_X1    g482(.A(new_n551), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n582), .B1(new_n669), .B2(new_n577), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n602), .B1(new_n670), .B2(new_n296), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n597), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n373), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n410), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n668), .A2(new_n420), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n667), .A2(new_n653), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT95), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  NAND2_X1  g493(.A1(new_n373), .A2(new_n624), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n659), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n657), .A2(new_n662), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  NAND3_X1  g497(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n646), .A2(new_n471), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n481), .A3(new_n472), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n684), .A2(new_n661), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n634), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n640), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NOR2_X1   g506(.A1(new_n638), .A2(new_n686), .ZN(new_n693));
  INV_X1    g507(.A(new_n412), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n581), .B2(new_n597), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(new_n607), .A3(new_n653), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND2_X1  g511(.A1(new_n684), .A2(KEYINPUT96), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT96), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n522), .A2(new_n699), .A3(new_n524), .A4(new_n526), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n638), .A2(new_n686), .A3(new_n419), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n601), .A2(new_n602), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n562), .A2(new_n541), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n592), .B1(new_n704), .B2(new_n577), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n703), .B1(new_n589), .B2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n701), .A2(new_n675), .A3(new_n702), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  AND3_X1   g522(.A1(new_n706), .A2(new_n653), .A3(new_n681), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n693), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  AOI21_X1  g525(.A(new_n661), .B1(new_n698), .B2(new_n700), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n475), .A2(KEYINPUT97), .A3(new_n426), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT97), .B1(new_n475), .B2(new_n426), .ZN(new_n714));
  OAI211_X1 g528(.A(G469), .B(new_n478), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n645), .B1(new_n715), .B2(new_n647), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n300), .A2(new_n301), .A3(new_n420), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT98), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n716), .A2(KEYINPUT98), .A3(new_n718), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n712), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n598), .A2(new_n524), .A3(new_n522), .A4(new_n526), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n721), .B2(new_n722), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT99), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n681), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n684), .A2(new_n661), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n716), .A2(KEYINPUT98), .A3(new_n718), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT98), .B1(new_n716), .B2(new_n718), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n730), .B(new_n681), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT42), .B1(new_n733), .B2(KEYINPUT99), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n725), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n315), .ZN(G33));
  OAI211_X1 g550(.A(new_n730), .B(new_n660), .C1(new_n731), .C2(new_n732), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT100), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n723), .A2(new_n739), .A3(new_n730), .A4(new_n660), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  AOI21_X1  g556(.A(KEYINPUT45), .B1(new_n476), .B2(new_n478), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n471), .ZN(new_n744));
  OAI211_X1 g558(.A(KEYINPUT45), .B(new_n478), .C1(new_n713), .C2(new_n714), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n474), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n472), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT101), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n749), .A2(KEYINPUT101), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n645), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n665), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT102), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(KEYINPUT102), .A3(new_n665), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n674), .A2(new_n624), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT103), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT43), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT104), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n653), .A2(new_n603), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(KEYINPUT44), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT44), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n717), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n759), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT105), .B(G137), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G39));
  NAND2_X1  g584(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n754), .A2(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n661), .A2(new_n684), .A3(new_n681), .A4(new_n718), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n774));
  OAI211_X1 g588(.A(new_n772), .B(new_n773), .C1(new_n754), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  INV_X1    g590(.A(new_n685), .ZN(new_n777));
  INV_X1    g591(.A(new_n472), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT49), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n760), .A2(new_n421), .A3(new_n645), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n780), .A2(KEYINPUT49), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n783), .A2(new_n784), .A3(new_n668), .A4(new_n673), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n701), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n657), .B(new_n662), .C1(new_n660), .C2(new_n681), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n710), .ZN(new_n790));
  INV_X1    g604(.A(new_n638), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n673), .A3(new_n675), .A4(new_n716), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n659), .B(KEYINPUT108), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n522), .A2(new_n524), .A3(new_n652), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n788), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(new_n797), .ZN(new_n800));
  INV_X1    g614(.A(new_n792), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT52), .A3(new_n710), .A4(new_n789), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n661), .A2(new_n694), .A3(new_n659), .A4(new_n717), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n723), .A2(new_n709), .B1(new_n657), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n739), .B1(new_n727), .B2(new_n660), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n680), .A2(new_n639), .ZN(new_n811));
  INV_X1    g625(.A(new_n422), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n300), .B2(new_n301), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n527), .A2(new_n604), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n696), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n599), .A2(new_n654), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n687), .B1(new_n634), .B2(new_n640), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n707), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n810), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n734), .A2(new_n729), .ZN(new_n821));
  INV_X1    g635(.A(new_n725), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT107), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n688), .A2(new_n691), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n696), .A2(new_n599), .A3(new_n654), .A4(new_n815), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n741), .A3(new_n707), .A4(new_n807), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT107), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n828), .A2(new_n829), .A3(new_n735), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n805), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g645(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n832));
  OAI21_X1  g646(.A(new_n787), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n829), .B1(new_n828), .B2(new_n735), .ZN(new_n834));
  INV_X1    g648(.A(new_n819), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n723), .A2(new_n709), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n806), .A2(new_n657), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n740), .B2(new_n738), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n823), .A2(new_n835), .A3(new_n839), .A4(KEYINPUT107), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n804), .B1(new_n834), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n832), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(KEYINPUT112), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n802), .A2(new_n710), .A3(new_n789), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT110), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT52), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n804), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n824), .B2(new_n830), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n833), .A2(new_n843), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(KEYINPUT54), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n828), .A2(new_n850), .A3(new_n735), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n855), .B(new_n856), .C1(new_n841), .C2(new_n842), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n414), .A2(new_n701), .A3(new_n706), .A4(new_n762), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n668), .A2(new_n420), .A3(new_n686), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n859), .A2(KEYINPUT50), .A3(new_n860), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n414), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n686), .A2(new_n866), .A3(new_n717), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n762), .A2(new_n653), .A3(new_n706), .A4(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT113), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n597), .A2(new_n867), .A3(new_n527), .A4(new_n672), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n674), .A2(new_n870), .A3(new_n611), .A4(new_n623), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n865), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n772), .B1(new_n754), .B2(new_n774), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n779), .A2(new_n645), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n859), .A2(new_n718), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n872), .B(KEYINPUT51), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n712), .A2(new_n762), .A3(new_n867), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT114), .Z(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n859), .A2(new_n693), .ZN(new_n884));
  INV_X1    g698(.A(new_n680), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n870), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n884), .A2(G952), .A3(new_n272), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n882), .B2(KEYINPUT48), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT115), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n883), .A2(new_n888), .A3(KEYINPUT115), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n879), .B(new_n880), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n853), .A2(new_n858), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n786), .B1(new_n892), .B2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n272), .A2(G952), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n249), .A2(new_n277), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT116), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n275), .B(KEYINPUT55), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n831), .A2(new_n832), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n296), .B1(new_n900), .B2(new_n855), .ZN(new_n901));
  AOI211_X1 g715(.A(KEYINPUT56), .B(new_n899), .C1(new_n901), .C2(G210), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n855), .B1(new_n841), .B2(new_n842), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(G210), .A3(G902), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT56), .B1(new_n904), .B2(KEYINPUT117), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(KEYINPUT117), .B2(new_n904), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n895), .B(new_n902), .C1(new_n899), .C2(new_n906), .ZN(G51));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  AOI211_X1 g722(.A(new_n296), .B(new_n746), .C1(new_n900), .C2(new_n855), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n473), .B(KEYINPUT118), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT57), .Z(new_n911));
  AOI21_X1  g725(.A(new_n856), .B1(new_n900), .B2(new_n855), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n858), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n909), .B1(new_n913), .B2(new_n470), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n908), .B1(new_n914), .B2(new_n895), .ZN(new_n915));
  INV_X1    g729(.A(new_n895), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n857), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n918), .A2(new_n911), .B1(new_n461), .B2(new_n469), .ZN(new_n919));
  OAI211_X1 g733(.A(KEYINPUT119), .B(new_n916), .C1(new_n919), .C2(new_n909), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n915), .A2(new_n920), .ZN(G54));
  NAND2_X1  g735(.A1(KEYINPUT58), .A2(G475), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT120), .Z(new_n923));
  AND3_X1   g737(.A1(new_n901), .A2(new_n356), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n356), .B1(new_n901), .B2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n895), .ZN(G60));
  OR2_X1    g740(.A1(new_n621), .A2(new_n622), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT59), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n918), .A2(new_n617), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n916), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n853), .B2(new_n858), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n927), .A2(new_n617), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT60), .Z(new_n936));
  AOI21_X1  g750(.A(new_n517), .B1(new_n903), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n895), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT61), .B1(new_n938), .B2(KEYINPUT121), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n903), .A2(new_n651), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G66));
  AOI21_X1  g756(.A(new_n272), .B1(new_n416), .B2(G224), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n819), .B(KEYINPUT122), .Z(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n272), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n897), .B1(G898), .B2(new_n272), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(G69));
  XOR2_X1   g762(.A(new_n790), .B(KEYINPUT125), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n678), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n775), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n718), .B1(new_n811), .B2(KEYINPUT126), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n666), .B(new_n954), .C1(KEYINPUT126), .C2(new_n811), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n730), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n768), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n272), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n567), .A2(new_n568), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT123), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n351), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT124), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n712), .A2(new_n791), .A3(new_n675), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n757), .B2(new_n758), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n949), .A2(new_n741), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n768), .A2(new_n823), .A3(new_n775), .A4(new_n967), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n966), .A2(new_n968), .A3(G953), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n963), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n963), .B(new_n975), .C1(new_n969), .C2(new_n971), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(G72));
  NOR2_X1   g791(.A1(new_n570), .A2(new_n545), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n966), .A2(new_n968), .A3(new_n945), .ZN(new_n979));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n978), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n952), .A2(new_n768), .A3(new_n956), .A4(new_n944), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n981), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n571), .B1(new_n569), .B2(new_n535), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n983), .A2(new_n987), .A3(new_n916), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n978), .A2(new_n982), .A3(new_n986), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n852), .B2(new_n989), .ZN(G57));
endmodule


