//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1381, new_n1382, new_n1383;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n203), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n210), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n214), .B(new_n225), .C1(new_n226), .C2(new_n220), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT0), .ZN(new_n228));
  INV_X1    g0028(.A(G50), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n227), .A2(KEYINPUT0), .ZN(new_n235));
  NAND4_X1  g0035(.A1(new_n223), .A2(new_n228), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n222), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT65), .Z(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n202), .ZN(new_n248));
  XOR2_X1   g0048(.A(KEYINPUT66), .B(G50), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G97), .B(G107), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G232), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G226), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT67), .B(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n255), .B1(new_n257), .B2(new_n258), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g0064(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  AOI21_X1  g0070(.A(G1), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n268), .A2(G274), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n263), .A2(new_n271), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(G238), .B2(new_n274), .ZN(new_n275));
  AND3_X1   g0075(.A1(new_n264), .A2(new_n265), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n265), .B1(new_n264), .B2(new_n275), .ZN(new_n277));
  OAI21_X1  g0077(.A(G169), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT14), .ZN(new_n279));
  INV_X1    g0079(.A(new_n276), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n264), .A2(KEYINPUT75), .A3(new_n275), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT13), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT75), .B1(new_n264), .B2(new_n275), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n280), .B(G179), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n285), .B(G169), .C1(new_n276), .C2(new_n277), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n279), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT68), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n231), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT69), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT69), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n289), .A2(new_n291), .A3(new_n294), .A4(new_n231), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G20), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n298), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G20), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n229), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT76), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT11), .ZN(new_n305));
  INV_X1    g0105(.A(G1), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G13), .A3(G20), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT70), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n306), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n311), .A2(KEYINPUT12), .A3(G68), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT12), .B1(new_n311), .B2(G68), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n309), .A2(new_n310), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n292), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n203), .B1(new_n306), .B2(G20), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n312), .A2(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n305), .A2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n304), .A2(KEYINPUT11), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n287), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n280), .B(G190), .C1(new_n282), .C2(new_n283), .ZN(new_n322));
  OAI21_X1  g0122(.A(G200), .B1(new_n276), .B2(new_n277), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n322), .A2(new_n318), .A3(new_n319), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n306), .B1(G41), .B2(G45), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n268), .A2(G232), .A3(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n272), .A2(new_n327), .A3(KEYINPUT78), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT78), .B1(new_n272), .B2(new_n327), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n260), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT77), .B1(new_n297), .B2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT77), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n331), .A2(new_n337), .B1(new_n297), .B2(new_n213), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n263), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n330), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(G169), .B1(new_n330), .B2(new_n339), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT79), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT79), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n330), .A2(new_n339), .A3(new_n340), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n330), .A2(new_n339), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(G169), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(G20), .B1(G159), .B2(new_n300), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n337), .A2(new_n350), .A3(new_n232), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G68), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n337), .B2(new_n232), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT16), .B(new_n349), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n349), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n256), .B2(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n334), .A2(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n336), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n203), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n354), .B(new_n292), .C1(new_n361), .C2(KEYINPUT16), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n296), .A2(new_n314), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT8), .B(G58), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n306), .B2(G20), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n363), .A2(new_n365), .B1(new_n314), .B2(new_n364), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n343), .A2(new_n347), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT18), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n343), .A2(new_n347), .A3(new_n367), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n367), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n346), .A2(G190), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n330), .A2(new_n339), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G200), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n372), .A2(KEYINPUT17), .A3(new_n373), .A4(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n373), .A2(new_n366), .A3(new_n362), .A4(new_n375), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT17), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n369), .A2(new_n371), .A3(new_n376), .A4(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n325), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n274), .A2(G226), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n272), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n256), .A2(G223), .A3(G1698), .ZN(new_n384));
  INV_X1    g0184(.A(G222), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n384), .B1(new_n217), .B2(new_n256), .C1(new_n261), .C2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n263), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(G179), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n306), .A2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n363), .A2(G50), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n232), .B1(new_n206), .B2(new_n229), .ZN(new_n392));
  INV_X1    g0192(.A(new_n298), .ZN(new_n393));
  INV_X1    g0193(.A(G150), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n364), .A2(new_n393), .B1(new_n394), .B2(new_n301), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n296), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n314), .A2(new_n229), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G169), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n389), .B(new_n399), .C1(new_n400), .C2(new_n388), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n388), .A2(KEYINPUT72), .A3(G200), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT72), .B1(new_n388), .B2(G200), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT10), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT9), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n398), .A2(new_n406), .B1(G190), .B2(new_n387), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(KEYINPUT9), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n404), .A2(new_n405), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n402), .A2(new_n403), .B1(new_n406), .B2(new_n398), .ZN(new_n410));
  INV_X1    g0210(.A(new_n407), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT10), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n401), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT67), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n414), .B1(new_n219), .B2(new_n256), .C1(new_n257), .C2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT71), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n268), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n420), .B2(new_n419), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n273), .B1(G244), .B2(new_n274), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n400), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n315), .A2(G77), .A3(new_n390), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n364), .A2(new_n301), .B1(new_n232), .B2(new_n217), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT15), .B(G87), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n393), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n292), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n426), .B(new_n430), .C1(G77), .C2(new_n311), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n422), .A2(new_n423), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n340), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n431), .B1(new_n433), .B2(G190), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n424), .A2(G200), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT73), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n413), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n413), .B2(new_n439), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n381), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT23), .B1(new_n232), .B2(G107), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT23), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n219), .A3(G20), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT84), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G116), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G20), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n232), .A2(KEYINPUT83), .A3(G33), .A4(G116), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n448), .A2(new_n449), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n445), .A4(new_n447), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT84), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  AND4_X1   g0258(.A1(new_n232), .A2(new_n332), .A3(new_n335), .A4(new_n336), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n213), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n256), .A2(new_n232), .A3(G87), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n459), .A2(new_n461), .B1(new_n462), .B2(new_n460), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n457), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n458), .B1(new_n457), .B2(new_n463), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n292), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n309), .A2(new_n219), .A3(new_n310), .ZN(new_n467));
  XOR2_X1   g0267(.A(new_n467), .B(KEYINPUT25), .Z(new_n468));
  NAND2_X1  g0268(.A1(new_n306), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n293), .A2(new_n311), .A3(new_n295), .A4(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n219), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n270), .A2(G1), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G264), .A3(new_n268), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT5), .B(G41), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(new_n268), .A3(G274), .A4(new_n474), .ZN(new_n480));
  INV_X1    g0280(.A(G294), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n297), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n415), .A2(new_n417), .A3(G250), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G257), .A2(G1698), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n332), .A2(new_n335), .A3(new_n336), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n478), .B(new_n480), .C1(new_n487), .C2(new_n268), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT85), .B1(new_n488), .B2(G169), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(KEYINPUT85), .A3(G169), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n260), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n491), .A2(new_n337), .B1(new_n297), .B2(new_n481), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n263), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(G179), .A3(new_n478), .A4(new_n480), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n473), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G200), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT87), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT87), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n488), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT86), .B1(new_n488), .B2(G190), .ZN(new_n502));
  INV_X1    g0302(.A(new_n478), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n492), .B2(new_n263), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT86), .ZN(new_n505));
  INV_X1    g0305(.A(G190), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n480), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n499), .A2(new_n501), .A3(new_n502), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n457), .A2(new_n463), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT24), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n457), .A2(new_n463), .A3(new_n458), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n471), .B1(new_n512), .B2(new_n292), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT88), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n496), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n496), .B2(new_n514), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n477), .A2(G270), .A3(new_n268), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n519), .A2(new_n480), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n220), .A2(new_n258), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n418), .B2(new_n226), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(new_n486), .B1(G303), .B2(new_n358), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n520), .B1(new_n524), .B2(new_n268), .ZN(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n314), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n266), .B1(new_n528), .B2(new_n290), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n526), .B1(new_n306), .B2(G33), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n311), .A2(new_n289), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(G20), .B1(G33), .B2(G283), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n297), .A2(G97), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n532), .A2(new_n533), .B1(G20), .B2(new_n526), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n292), .A2(KEYINPUT20), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT20), .B1(new_n292), .B2(new_n534), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n527), .B(new_n531), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n525), .A2(new_n537), .A3(G169), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT21), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n523), .A2(new_n486), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n358), .A2(G303), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n268), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n519), .A2(new_n480), .ZN(new_n544));
  OAI21_X1  g0344(.A(G200), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n537), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n521), .B1(new_n260), .B2(G257), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n542), .B1(new_n547), .B2(new_n337), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n263), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(G190), .A3(new_n520), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n544), .B1(new_n548), .B2(new_n263), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(new_n537), .A3(G179), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n525), .A2(new_n537), .A3(KEYINPUT21), .A4(G169), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n540), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n306), .A2(G45), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G250), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n263), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n268), .A2(G274), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n560), .B2(new_n474), .ZN(new_n561));
  INV_X1    g0361(.A(new_n451), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n218), .A2(new_n258), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n418), .B2(new_n212), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n562), .B1(new_n565), .B2(new_n486), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n561), .B(new_n340), .C1(new_n566), .C2(new_n268), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n559), .A2(new_n556), .B1(new_n263), .B2(new_n557), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n563), .B1(new_n260), .B2(G238), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n451), .B1(new_n569), .B2(new_n337), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n568), .B1(new_n570), .B2(new_n263), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n571), .B2(G169), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n309), .A2(new_n310), .A3(new_n428), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n297), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n334), .A2(G33), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n577), .A2(new_n232), .A3(G68), .A4(new_n332), .ZN(new_n578));
  OR2_X1    g0378(.A1(KEYINPUT82), .A2(G87), .ZN(new_n579));
  INV_X1    g0379(.A(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(KEYINPUT82), .A2(G87), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n219), .A4(new_n581), .ZN(new_n582));
  OR2_X1    g0382(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n583));
  NAND2_X1  g0383(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n255), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n582), .B1(new_n585), .B2(G20), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n232), .A2(G33), .A3(G97), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n587), .A2(new_n583), .A3(new_n584), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n578), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n574), .B1(new_n590), .B2(new_n292), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n428), .B2(new_n470), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n294), .B1(new_n529), .B2(new_n289), .ZN(new_n593));
  INV_X1    g0393(.A(new_n295), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n595), .A2(G87), .A3(new_n311), .A4(new_n469), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n561), .B(new_n506), .C1(new_n566), .C2(new_n268), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n571), .B2(G200), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n573), .A2(new_n592), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n477), .A2(G257), .A3(new_n268), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n480), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT80), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT80), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n601), .A2(new_n604), .A3(new_n480), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT4), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n218), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n256), .A2(new_n260), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G33), .A2(G283), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n336), .A2(new_n357), .A3(G250), .A4(G1698), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n260), .A2(G244), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n607), .B1(new_n613), .B2(new_n337), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n268), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n400), .B1(new_n606), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n595), .A2(G97), .A3(new_n311), .A4(new_n469), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT6), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n618), .A2(new_n580), .A3(G107), .ZN(new_n619));
  XNOR2_X1  g0419(.A(G97), .B(G107), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n621), .A2(new_n232), .B1(new_n217), .B2(new_n301), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n219), .B1(new_n356), .B2(new_n359), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n292), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n314), .A2(new_n580), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n617), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n418), .A2(new_n218), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT4), .B1(new_n627), .B2(new_n486), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n263), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(new_n340), .A3(new_n603), .A4(new_n605), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n616), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(G200), .B1(new_n606), .B2(new_n615), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n620), .A2(new_n618), .ZN(new_n634));
  INV_X1    g0434(.A(new_n619), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n636), .A2(G20), .B1(G77), .B2(new_n300), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n356), .A2(new_n359), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G107), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(new_n292), .B1(new_n580), .B2(new_n314), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n630), .A2(G190), .A3(new_n603), .A4(new_n605), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n633), .A2(new_n641), .A3(new_n642), .A4(new_n617), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n555), .A2(new_n600), .A3(new_n632), .A4(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n444), .A2(new_n518), .A3(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n401), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n369), .A2(new_n371), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n324), .A2(new_n434), .A3(new_n432), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n321), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n376), .A2(new_n379), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n647), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n409), .A2(new_n412), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n646), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n470), .A2(new_n428), .ZN(new_n657));
  INV_X1    g0457(.A(new_n292), .ZN(new_n658));
  AND2_X1   g0458(.A1(G33), .A2(G97), .ZN(new_n659));
  AND2_X1   g0459(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g0460(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n232), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n588), .B1(new_n663), .B2(new_n582), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n664), .B2(new_n578), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n657), .A2(new_n665), .A3(new_n574), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n572), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n616), .A2(new_n626), .A3(new_n631), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n561), .B1(new_n566), .B2(new_n268), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n400), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n590), .A2(new_n292), .ZN(new_n671));
  INV_X1    g0471(.A(new_n574), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n567), .B(new_n670), .C1(new_n673), .C2(new_n657), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n599), .A2(new_n591), .A3(new_n596), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n668), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n667), .B1(new_n676), .B2(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n591), .A2(new_n596), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n669), .A2(new_n497), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n598), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT89), .B1(new_n680), .B2(new_n667), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT89), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n675), .A2(new_n674), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n681), .A2(new_n682), .A3(new_n668), .A4(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n643), .A2(new_n632), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n554), .A2(new_n553), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n400), .B1(new_n549), .B2(new_n520), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT21), .B1(new_n689), .B2(new_n537), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT90), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT90), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n540), .A2(new_n692), .A3(new_n553), .A4(new_n554), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n687), .B1(new_n694), .B2(new_n496), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n675), .A2(new_n674), .A3(new_n683), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n683), .B1(new_n675), .B2(new_n674), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n514), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n686), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n656), .B1(new_n444), .B2(new_n701), .ZN(G369));
  NAND3_X1  g0502(.A1(new_n306), .A2(new_n232), .A3(G13), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G213), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G343), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n513), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n518), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n495), .ZN(new_n712));
  INV_X1    g0512(.A(new_n489), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n712), .A2(new_n713), .B1(new_n466), .B2(new_n472), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n714), .B2(new_n708), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n555), .B1(new_n546), .B2(new_n709), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n537), .A2(new_n708), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n694), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n688), .A2(new_n690), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n708), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n501), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n500), .B1(new_n488), .B2(new_n497), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n507), .A2(new_n502), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n473), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT88), .B1(new_n728), .B2(new_n714), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n496), .A2(new_n514), .A3(new_n515), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n723), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n496), .A2(new_n708), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n720), .A2(new_n733), .ZN(G399));
  NOR2_X1   g0534(.A1(new_n225), .A2(G41), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n230), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n582), .A2(G116), .ZN(new_n737));
  OAI21_X1  g0537(.A(G1), .B1(new_n225), .B2(G41), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT28), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n681), .A2(new_n668), .A3(new_n684), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT26), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n680), .A2(new_n632), .A3(new_n667), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n667), .B1(new_n743), .B2(new_n682), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n681), .A2(new_n514), .A3(new_n684), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT93), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n687), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n495), .A2(new_n489), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n721), .B1(new_n748), .B2(new_n513), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n643), .A2(new_n632), .A3(KEYINPUT93), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n742), .B(new_n744), .C1(new_n745), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT94), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n752), .A2(new_n753), .A3(new_n709), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n752), .B2(new_n709), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT29), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n708), .B1(new_n686), .B2(new_n699), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(KEYINPUT29), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT30), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n504), .A2(new_n552), .A3(new_n571), .A4(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n630), .A2(new_n603), .A3(new_n605), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT91), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g0565(.A(KEYINPUT91), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n606), .A2(new_n615), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n525), .A2(new_n340), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n478), .B1(new_n487), .B2(new_n268), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n669), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n767), .A2(new_n768), .A3(new_n770), .A4(KEYINPUT30), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n552), .A2(G179), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n772), .A2(new_n762), .A3(new_n488), .A4(new_n669), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n765), .A2(new_n766), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n708), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT31), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT92), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n771), .A2(new_n773), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n763), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n777), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(KEYINPUT31), .B1(new_n774), .B2(new_n708), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n776), .B(new_n709), .C1(new_n779), .C2(new_n763), .ZN(new_n784));
  OAI21_X1  g0584(.A(KEYINPUT92), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n644), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n786), .B(new_n709), .C1(new_n516), .C2(new_n517), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n782), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n756), .A2(new_n759), .B1(G330), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n740), .B1(new_n789), .B2(G1), .ZN(G364));
  AND2_X1   g0590(.A1(new_n232), .A2(G13), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n306), .B1(new_n791), .B2(G45), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n735), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n225), .A2(new_n358), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G355), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G116), .B2(new_n224), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n250), .A2(G45), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n486), .A2(new_n225), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n270), .B2(new_n230), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n797), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n231), .B1(G20), .B2(new_n400), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n794), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n232), .A2(new_n340), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G200), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n506), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n229), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G179), .A2(G200), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(G20), .A3(new_n506), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G159), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT32), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n579), .A2(new_n581), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n232), .A2(new_n506), .A3(new_n497), .A4(G179), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n814), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n811), .A2(G190), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n232), .B1(new_n815), .B2(G190), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n823), .A2(G68), .B1(G97), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT96), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n810), .A2(G190), .A3(new_n497), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G190), .A2(G200), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n810), .A2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n828), .A2(new_n202), .B1(new_n830), .B2(new_n217), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT95), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n232), .A2(new_n497), .A3(G179), .A4(G190), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n256), .B1(new_n834), .B2(new_n219), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(KEYINPUT95), .B2(new_n831), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n822), .A2(new_n827), .A3(new_n832), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G322), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n828), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n358), .B1(new_n830), .B2(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(G329), .C2(new_n817), .ZN(new_n842));
  XNOR2_X1  g0642(.A(KEYINPUT97), .B(G326), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n813), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(KEYINPUT33), .B(G317), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n823), .A2(new_n845), .B1(G294), .B2(new_n825), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n821), .A2(G303), .B1(new_n833), .B2(G283), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n842), .A2(new_n844), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n837), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n809), .B1(new_n849), .B2(new_n806), .ZN(new_n850));
  INV_X1    g0650(.A(new_n805), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n718), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n794), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n719), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n718), .A2(G330), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT98), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G396));
  NAND2_X1  g0658(.A1(new_n431), .A2(new_n708), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT100), .Z(new_n860));
  AOI22_X1  g0660(.A1(new_n438), .A2(new_n860), .B1(new_n432), .B2(new_n434), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n432), .A2(new_n434), .A3(new_n709), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n757), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n788), .A2(G330), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n794), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n806), .ZN(new_n870));
  INV_X1    g0670(.A(new_n828), .ZN(new_n871));
  INV_X1    g0671(.A(new_n830), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n871), .A2(G143), .B1(new_n872), .B2(G159), .ZN(new_n873));
  INV_X1    g0673(.A(G137), .ZN(new_n874));
  INV_X1    g0674(.A(new_n823), .ZN(new_n875));
  OAI221_X1 g0675(.A(new_n873), .B1(new_n813), .B2(new_n874), .C1(new_n394), .C2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT34), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(G132), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n486), .B1(new_n879), .B2(new_n816), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n834), .A2(new_n203), .B1(new_n202), .B2(new_n824), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n880), .B(new_n881), .C1(G50), .C2(new_n821), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(G303), .ZN(new_n885));
  INV_X1    g0685(.A(new_n821), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n813), .A2(new_n885), .B1(new_n219), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(G87), .B2(new_n833), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n256), .B1(new_n871), .B2(G294), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n872), .A2(G116), .B1(new_n817), .B2(G311), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n823), .A2(G283), .B1(G97), .B2(new_n825), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n870), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n806), .A2(new_n803), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n853), .B(new_n893), .C1(new_n217), .C2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT99), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n804), .B2(new_n864), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT101), .Z(new_n898));
  NOR2_X1   g0698(.A1(new_n869), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(G384));
  NOR2_X1   g0700(.A1(new_n321), .A2(new_n708), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n354), .A2(new_n296), .ZN(new_n903));
  INV_X1    g0703(.A(new_n353), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(G68), .A3(new_n351), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT16), .B1(new_n905), .B2(new_n349), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n366), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n706), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n380), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n367), .A2(new_n908), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n368), .A2(new_n912), .A3(new_n377), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n343), .A2(new_n347), .A3(new_n907), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n915), .A2(new_n377), .A3(new_n909), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n916), .B2(new_n912), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n911), .A2(new_n917), .A3(KEYINPUT38), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n911), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n913), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n368), .A2(new_n377), .A3(new_n913), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n380), .A2(new_n921), .B1(new_n923), .B2(new_n914), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT103), .B1(new_n924), .B2(KEYINPUT38), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n902), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n911), .A2(new_n917), .A3(KEYINPUT38), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(KEYINPUT38), .B2(new_n924), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n928), .A2(KEYINPUT103), .A3(KEYINPUT39), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n901), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n700), .A2(new_n709), .A3(new_n864), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n862), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n320), .A2(new_n708), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n321), .A2(new_n324), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n287), .A2(new_n320), .A3(new_n708), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n932), .A2(KEYINPUT102), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT102), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n863), .B1(new_n757), .B2(new_n864), .ZN(new_n939));
  INV_X1    g0739(.A(new_n936), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n920), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n647), .A2(new_n706), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n930), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n381), .ZN(new_n946));
  INV_X1    g0746(.A(new_n443), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n947), .B2(new_n441), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n756), .A2(new_n948), .A3(new_n759), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT104), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n756), .A2(new_n948), .A3(KEYINPUT104), .A4(new_n759), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n655), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n945), .B(new_n953), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n863), .B(new_n861), .C1(new_n934), .C2(new_n935), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n774), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n783), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT105), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n957), .A2(new_n958), .A3(new_n787), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n957), .B2(new_n787), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n928), .B(new_n955), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT40), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n936), .A2(new_n864), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n708), .B(new_n644), .C1(new_n729), .C2(new_n730), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n774), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n777), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT105), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n957), .A2(new_n958), .A3(new_n787), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n911), .A2(new_n917), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT38), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT40), .B1(new_n972), .B2(new_n927), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n962), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n975), .B(new_n948), .C1(new_n959), .C2(new_n960), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n961), .A2(KEYINPUT40), .B1(new_n969), .B2(new_n973), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n959), .A2(new_n960), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n444), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(G330), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n954), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(KEYINPUT106), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(KEYINPUT106), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n954), .A2(new_n980), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n791), .A2(new_n306), .ZN(new_n985));
  NOR4_X1   g0785(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n636), .A2(KEYINPUT35), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n636), .A2(KEYINPUT35), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n987), .A2(G116), .A3(new_n233), .A4(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT36), .Z(new_n990));
  OAI211_X1 g0790(.A(new_n230), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n229), .A2(G68), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n306), .B(G13), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n986), .A2(new_n990), .A3(new_n993), .ZN(G367));
  NAND2_X1  g0794(.A1(new_n626), .A2(new_n708), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n747), .A2(new_n750), .A3(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(new_n496), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n708), .B1(new_n997), .B2(new_n632), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT42), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n668), .A2(new_n708), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n999), .B1(new_n731), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT107), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT107), .B1(new_n998), .B2(new_n1002), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1001), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n722), .B1(new_n516), .B2(new_n517), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT42), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1005), .A2(new_n1006), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n678), .A2(new_n708), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n674), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n698), .B2(new_n1012), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT43), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1011), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1009), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1019), .A2(new_n1015), .A3(new_n1014), .A4(new_n1006), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n715), .A2(new_n719), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n1001), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n1018), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1023), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n735), .B(KEYINPUT41), .Z(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT108), .B1(new_n733), .B2(new_n1001), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n732), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1008), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT108), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n1007), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1028), .A2(KEYINPUT44), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1008), .A2(new_n1001), .A3(new_n1029), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT45), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT44), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1021), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT44), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1032), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1031), .B1(new_n1030), .B2(new_n1007), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1043), .A2(new_n720), .A3(new_n1036), .A4(new_n1033), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n723), .B1(new_n496), .B2(new_n709), .C1(new_n518), .C2(new_n710), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n1008), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n719), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1039), .A2(new_n789), .A3(new_n1044), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1027), .B1(new_n1049), .B2(new_n789), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1026), .B1(new_n1050), .B2(new_n793), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1014), .A2(new_n805), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n875), .A2(new_n481), .B1(new_n824), .B2(new_n219), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G97), .B2(new_n833), .ZN(new_n1054));
  INV_X1    g0854(.A(G283), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n828), .A2(new_n885), .B1(new_n830), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G317), .B2(new_n817), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n486), .B1(new_n812), .B2(G311), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n821), .A2(G116), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT46), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1054), .A2(new_n1057), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n834), .A2(new_n217), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G143), .B2(new_n812), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n256), .B1(new_n828), .B2(new_n394), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G50), .B2(new_n872), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n823), .A2(G159), .B1(G68), .B2(new_n825), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n821), .A2(G58), .B1(new_n817), .B2(G137), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT109), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1061), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT47), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n806), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n807), .B1(new_n224), .B2(new_n428), .C1(new_n800), .C2(new_n245), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1052), .A2(new_n794), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1051), .A2(new_n1074), .ZN(G387));
  OR2_X1    g0875(.A1(new_n242), .A2(new_n270), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1076), .A2(new_n799), .B1(new_n737), .B2(new_n795), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n364), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n229), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n270), .B1(new_n203), .B2(new_n217), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1080), .A2(new_n737), .A3(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1077), .A2(new_n1082), .B1(G107), .B2(new_n224), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n853), .B1(new_n1083), .B2(new_n807), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n824), .A2(new_n428), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n812), .B2(G159), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n886), .A2(new_n217), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1078), .B2(new_n823), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n828), .A2(new_n229), .B1(new_n830), .B2(new_n203), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G150), .B2(new_n817), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n337), .B1(G97), .B2(new_n833), .ZN(new_n1091));
  AND4_X1   g0891(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n886), .A2(new_n481), .B1(new_n1055), .B2(new_n824), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n871), .A2(G317), .B1(new_n872), .B2(G303), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n813), .B2(new_n838), .C1(new_n840), .C2(new_n875), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT48), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT49), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT111), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n337), .B1(new_n843), .B2(new_n816), .C1(new_n834), .C2(new_n526), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1099), .B2(KEYINPUT111), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1092), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1084), .B1(new_n1103), .B2(new_n870), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n715), .B2(new_n805), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1048), .A2(new_n793), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT110), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1048), .A2(KEYINPUT110), .A3(new_n793), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1048), .A2(new_n789), .A3(KEYINPUT112), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT112), .B1(new_n1048), .B2(new_n789), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1048), .A2(new_n789), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1112), .A2(new_n735), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1110), .B1(new_n1111), .B2(new_n1114), .ZN(G393));
  NAND3_X1  g0915(.A1(new_n1039), .A2(new_n793), .A3(new_n1044), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n807), .B1(new_n580), .B2(new_n224), .C1(new_n800), .C2(new_n253), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n794), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n875), .A2(new_n885), .B1(new_n824), .B2(new_n526), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n358), .B1(new_n816), .B2(new_n838), .C1(new_n830), .C2(new_n481), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n886), .A2(new_n1055), .B1(new_n834), .B2(new_n219), .ZN(new_n1121));
  OR3_X1    g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G317), .A2(new_n812), .B1(new_n871), .B2(G311), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G150), .A2(new_n812), .B1(new_n871), .B2(G159), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT51), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n823), .A2(G50), .B1(G77), .B2(new_n825), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n872), .A2(new_n1078), .B1(new_n817), .B2(G143), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n821), .A2(G68), .B1(new_n833), .B2(G87), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1128), .A2(new_n486), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1122), .A2(new_n1125), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1118), .B1(new_n1132), .B2(new_n806), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1001), .B2(new_n851), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1049), .A2(new_n735), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1039), .A2(new_n1044), .B1(new_n789), .B2(new_n1048), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1116), .B(new_n1134), .C1(new_n1135), .C2(new_n1136), .ZN(G390));
  OAI21_X1  g0937(.A(new_n744), .B1(new_n751), .B2(new_n745), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n742), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n709), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT94), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n752), .A2(new_n753), .A3(new_n709), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n862), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n438), .A2(new_n860), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n435), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1145), .A3(new_n936), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n928), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(new_n901), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n939), .A2(new_n940), .B1(new_n321), .B2(new_n708), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n925), .A2(new_n927), .A3(new_n972), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(KEYINPUT39), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1147), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1150), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n788), .A2(G330), .A3(new_n864), .A4(new_n936), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1149), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1151), .A2(KEYINPUT39), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1158), .A2(new_n1150), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1159));
  INV_X1    g0959(.A(G330), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n967), .B2(new_n968), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n955), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1157), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1158), .A2(new_n803), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n894), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n794), .B1(new_n1078), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n821), .A2(G150), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT53), .Z(new_n1169));
  INV_X1    g0969(.A(G125), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n828), .A2(new_n879), .B1(new_n1170), .B2(new_n816), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT54), .B(G143), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n256), .B1(new_n830), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n823), .A2(G137), .B1(G159), .B2(new_n825), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n812), .A2(G128), .B1(G50), .B2(new_n833), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1169), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n875), .A2(new_n219), .B1(new_n203), .B2(new_n834), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n813), .A2(new_n1055), .B1(new_n213), .B2(new_n886), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n358), .B1(new_n816), .B2(new_n481), .C1(new_n830), .C2(new_n580), .ZN(new_n1180));
  OR3_X1    g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n828), .A2(new_n526), .B1(new_n824), .B2(new_n217), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT115), .Z(new_n1183));
  OAI21_X1  g0983(.A(new_n1177), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1167), .B1(new_n1184), .B2(new_n806), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1164), .A2(new_n793), .B1(new_n1165), .B2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n754), .A2(new_n755), .A3(new_n863), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1156), .B1(new_n1187), .B2(new_n861), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n936), .B1(new_n1161), .B2(new_n864), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n788), .A2(G330), .A3(new_n864), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1161), .A2(new_n955), .B1(new_n1190), .B2(new_n940), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1188), .A2(new_n1189), .B1(new_n1191), .B2(new_n939), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n951), .A2(new_n952), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1161), .A2(new_n948), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n656), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1163), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n735), .B1(new_n1195), .B2(new_n1163), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(KEYINPUT114), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT114), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1194), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n655), .B(new_n1200), .C1(new_n951), .C2(new_n952), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1149), .A2(new_n1155), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n955), .A3(new_n1161), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1203), .A3(new_n1157), .A4(new_n1192), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1199), .B1(new_n1204), .B2(new_n735), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1186), .B1(new_n1198), .B2(new_n1205), .ZN(G378));
  NAND3_X1  g1006(.A1(new_n930), .A2(new_n943), .A3(new_n944), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n398), .B(new_n908), .C1(new_n654), .C2(new_n401), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n413), .B1(new_n399), .B2(new_n706), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n975), .B2(G330), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n977), .A2(new_n1160), .A3(new_n1213), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1207), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1213), .B1(new_n977), .B2(new_n1160), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n975), .A2(G330), .A3(new_n1214), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n945), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1213), .A2(new_n803), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n794), .B1(G50), .B2(new_n1166), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n875), .A2(new_n879), .B1(new_n813), .B2(new_n1170), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n871), .A2(G128), .B1(new_n872), .B2(G137), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n886), .B2(new_n1172), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G150), .C2(new_n825), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT116), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(G124), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(G124), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n817), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n297), .A3(new_n269), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G159), .B2(new_n833), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1229), .A2(new_n1230), .A3(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n871), .A2(G107), .B1(G283), .B2(new_n817), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n428), .B2(new_n830), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1087), .B(new_n1239), .C1(G68), .C2(new_n825), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n813), .A2(new_n526), .B1(new_n202), .B2(new_n834), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G97), .B2(new_n823), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1240), .A2(new_n269), .A3(new_n337), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT58), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G50), .B1(new_n297), .B2(new_n269), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n486), .B2(G41), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1237), .A2(new_n1245), .A3(new_n1246), .A4(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1223), .B1(new_n1249), .B2(new_n806), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1221), .A2(new_n793), .B1(new_n1222), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n758), .B1(new_n1252), .B2(KEYINPUT29), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT104), .B1(new_n1253), .B2(new_n948), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n952), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n656), .B(new_n1194), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT117), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT117), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n953), .A2(new_n1258), .A3(new_n1194), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1195), .A2(new_n1163), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT57), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT118), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1217), .A2(new_n1220), .A3(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n945), .A2(KEYINPUT118), .A3(new_n1219), .A4(new_n1218), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n735), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1257), .B(new_n1259), .C1(new_n1163), .C2(new_n1195), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT57), .B1(new_n1268), .B2(new_n1221), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1251), .B1(new_n1267), .B2(new_n1269), .ZN(G375));
  AOI21_X1  g1070(.A(new_n853), .B1(new_n203), .B2(new_n894), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G116), .A2(new_n823), .B1(new_n812), .B2(G294), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n580), .B2(new_n886), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n256), .B1(new_n817), .B2(G303), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n1274), .B1(new_n219), .B2(new_n830), .C1(new_n1055), .C2(new_n828), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1273), .A2(new_n1275), .A3(new_n1062), .A4(new_n1085), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n812), .A2(G132), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1277), .B1(new_n874), .B2(new_n828), .C1(new_n875), .C2(new_n1172), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(KEYINPUT119), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n824), .A2(new_n229), .ZN(new_n1280));
  INV_X1    g1080(.A(G128), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n830), .A2(new_n394), .B1(new_n816), .B2(new_n1281), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1280), .B(new_n1282), .C1(G159), .C2(new_n821), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n486), .B1(new_n834), .B2(new_n202), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT120), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1283), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1276), .B1(new_n1279), .B2(new_n1288), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n1271), .B1(new_n870), .B2(new_n1289), .C1(new_n936), .C2(new_n804), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1192), .B2(new_n793), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1027), .B1(new_n1201), .B2(new_n1192), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1192), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1256), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1293), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(G381));
  XOR2_X1   g1098(.A(G375), .B(KEYINPUT121), .Z(new_n1299));
  INV_X1    g1099(.A(G378), .ZN(new_n1300));
  OR4_X1    g1100(.A1(G396), .A2(G390), .A3(G393), .A4(G384), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1301), .A2(G387), .A3(G381), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1299), .A2(new_n1300), .A3(new_n1302), .ZN(G407));
  NAND2_X1  g1103(.A1(new_n707), .A2(G213), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1299), .A2(new_n1300), .A3(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G407), .A2(new_n1306), .A3(G213), .ZN(G409));
  OAI211_X1 g1107(.A(G378), .B(new_n1251), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1222), .A2(new_n1250), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1264), .A2(new_n793), .A3(new_n1265), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1268), .A2(new_n1221), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1309), .B(new_n1310), .C1(new_n1311), .C2(new_n1027), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1205), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1204), .A2(new_n1199), .A3(new_n735), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1196), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1312), .A2(new_n1315), .A3(new_n1186), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1308), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1195), .A2(KEYINPUT60), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1318), .A2(new_n1296), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1256), .A2(new_n1295), .A3(KEYINPUT60), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n735), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1292), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n899), .ZN(new_n1323));
  OAI211_X1 g1123(.A(G384), .B(new_n1292), .C1(new_n1319), .C2(new_n1321), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1317), .A2(new_n1304), .A3(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT122), .ZN(new_n1330));
  INV_X1    g1130(.A(G390), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1330), .B1(G387), .B2(new_n1331), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(G393), .B(G396), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1051), .A2(new_n1074), .A3(G390), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(G390), .B1(new_n1051), .B2(new_n1074), .ZN(new_n1336));
  OAI22_X1  g1136(.A1(new_n1332), .A2(new_n1333), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1336), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(G393), .B(new_n857), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1330), .A4(new_n1334), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1337), .A2(new_n1338), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(KEYINPUT123), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT123), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1337), .A2(new_n1344), .A3(new_n1341), .A4(new_n1338), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1317), .A2(new_n1304), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1305), .A2(G2897), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1323), .A2(new_n1324), .A3(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1347), .A2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1329), .A2(new_n1346), .A3(new_n1352), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1323), .A2(KEYINPUT63), .A3(new_n1324), .ZN(new_n1354));
  AND4_X1   g1154(.A1(KEYINPUT124), .A2(new_n1317), .A3(new_n1304), .A4(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1305), .B1(new_n1308), .B2(new_n1316), .ZN(new_n1356));
  AOI21_X1  g1156(.A(KEYINPUT124), .B1(new_n1356), .B2(new_n1354), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1355), .A2(new_n1357), .ZN(new_n1358));
  OAI21_X1  g1158(.A(KEYINPUT125), .B1(new_n1353), .B2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1356), .A2(new_n1354), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT124), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1356), .A2(KEYINPUT124), .A3(new_n1354), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT125), .ZN(new_n1365));
  AOI22_X1  g1165(.A1(new_n1343), .A2(new_n1345), .B1(new_n1347), .B2(new_n1351), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1364), .A2(new_n1365), .A3(new_n1329), .A4(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1359), .A2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1337), .A2(new_n1341), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1327), .A2(KEYINPUT126), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT62), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1372), .A2(new_n1338), .A3(new_n1352), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1369), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1368), .A2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1376), .A2(KEYINPUT127), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT127), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1368), .A2(new_n1375), .A3(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1377), .A2(new_n1379), .ZN(G405));
  NAND2_X1  g1180(.A1(G375), .A2(new_n1300), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1381), .A2(new_n1308), .ZN(new_n1382));
  XNOR2_X1  g1182(.A(new_n1382), .B(new_n1326), .ZN(new_n1383));
  XNOR2_X1  g1183(.A(new_n1383), .B(new_n1369), .ZN(G402));
endmodule


