//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT87), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT86), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT85), .B(G224), .Z(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT7), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT64), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT64), .A2(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n197), .B1(new_n200), .B2(G143), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n196), .A2(G143), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n200), .B2(G143), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(new_n208), .B2(new_n202), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n196), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT64), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(G143), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n207), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n213), .A2(new_n206), .A3(new_n214), .A4(new_n202), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n205), .B1(new_n209), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G125), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(new_n214), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n213), .A2(new_n223), .A3(new_n214), .A4(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G125), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n200), .B2(G143), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n201), .B1(new_n228), .B2(new_n219), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  AOI211_X1 g044(.A(new_n190), .B(new_n195), .C1(new_n218), .C2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n213), .A2(new_n214), .A3(new_n202), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n233), .A2(new_n215), .B1(new_n201), .B2(new_n204), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n230), .B1(new_n226), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT86), .B1(new_n235), .B2(new_n194), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G104), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G107), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(G107), .ZN(new_n241));
  OAI21_X1  g055(.A(G101), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT3), .B1(new_n238), .B2(G107), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n244));
  INV_X1    g058(.A(G107), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G104), .ZN(new_n246));
  INV_X1    g060(.A(G101), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n243), .A2(new_n246), .A3(new_n247), .A4(new_n239), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT68), .A2(G119), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT68), .A2(G119), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(G116), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(G113), .B1(new_n252), .B2(KEYINPUT5), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n250), .A2(KEYINPUT69), .A3(G116), .A4(new_n251), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT68), .A2(G119), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT68), .A2(G119), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT69), .B1(new_n257), .B2(G119), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n254), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n253), .B1(new_n261), .B2(KEYINPUT5), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT2), .B(G113), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n252), .A2(new_n259), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n254), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n249), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n249), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n264), .B2(new_n254), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n268), .B(new_n269), .C1(new_n271), .C2(new_n253), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G110), .B(G122), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT8), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n218), .A2(KEYINPUT7), .A3(new_n193), .A4(new_n230), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n189), .B1(new_n237), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n243), .A2(new_n246), .A3(new_n239), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G101), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(G101), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT4), .A3(new_n248), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n264), .A2(new_n263), .A3(new_n254), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n282), .B(new_n284), .C1(new_n285), .C2(new_n265), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT82), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n284), .A2(new_n282), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT82), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n264), .A2(new_n263), .A3(new_n254), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n268), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n287), .A2(new_n292), .A3(new_n272), .A4(new_n274), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n233), .A2(new_n215), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n226), .B1(new_n295), .B2(new_n205), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n194), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n190), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n235), .A2(KEYINPUT86), .A3(new_n194), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n300), .A2(KEYINPUT87), .A3(new_n277), .A4(new_n276), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n279), .A2(new_n293), .A3(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n274), .B(KEYINPUT83), .Z(new_n303));
  OAI21_X1  g117(.A(new_n272), .B1(new_n286), .B2(KEYINPUT82), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n289), .B1(new_n288), .B2(new_n291), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n293), .A3(KEYINPUT6), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT84), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n306), .A2(KEYINPUT6), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n306), .A2(new_n293), .A3(KEYINPUT84), .A4(KEYINPUT6), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n235), .B(new_n192), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n309), .A2(new_n310), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n302), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G210), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n302), .A2(new_n313), .A3(new_n314), .A4(new_n316), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n188), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT9), .B(G234), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT77), .ZN(new_n322));
  OAI21_X1  g136(.A(G221), .B1(new_n322), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(G469), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G140), .ZN(new_n325));
  INV_X1    g139(.A(G953), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(G227), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n325), .B(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n223), .B1(new_n208), .B2(new_n220), .ZN(new_n329));
  INV_X1    g143(.A(new_n224), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n219), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n208), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n213), .A2(new_n214), .ZN(new_n335));
  INV_X1    g149(.A(new_n333), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT78), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n269), .B1(new_n331), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n225), .A2(new_n249), .A3(new_n229), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G134), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(G137), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT11), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT11), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n342), .B2(G137), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(G137), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(G131), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT12), .B1(new_n341), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT12), .ZN(new_n351));
  INV_X1    g165(.A(new_n349), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n351), .B(new_n352), .C1(new_n339), .C2(new_n340), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n229), .B1(new_n329), .B2(new_n330), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n225), .A2(KEYINPUT70), .A3(new_n229), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n249), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n339), .A2(new_n359), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n288), .A2(new_n234), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n352), .A4(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n328), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n328), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(KEYINPUT79), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n339), .A2(new_n359), .B1(new_n288), .B2(new_n234), .ZN(new_n370));
  AOI211_X1 g184(.A(new_n369), .B(new_n352), .C1(new_n370), .C2(new_n361), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT80), .B1(new_n372), .B2(new_n349), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n368), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT79), .B1(new_n364), .B2(new_n367), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n366), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT78), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT78), .B1(new_n335), .B2(new_n336), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n249), .B1(new_n381), .B2(new_n225), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n363), .B1(new_n382), .B2(KEYINPUT10), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n225), .A2(KEYINPUT70), .A3(new_n229), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT70), .B1(new_n225), .B2(new_n229), .ZN(new_n385));
  INV_X1    g199(.A(new_n360), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n349), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n369), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n372), .A2(KEYINPUT80), .A3(new_n349), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n375), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n368), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT81), .A3(new_n366), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n324), .B1(new_n378), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n367), .B1(new_n391), .B2(new_n364), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n364), .A2(new_n367), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n354), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n324), .B(new_n314), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n324), .A2(new_n314), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n320), .B(new_n323), .C1(new_n395), .C2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(G475), .A2(G902), .ZN(new_n405));
  XNOR2_X1  g219(.A(G125), .B(G140), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n200), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n196), .B2(new_n406), .ZN(new_n408));
  INV_X1    g222(.A(G237), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n326), .A3(G214), .ZN(new_n410));
  INV_X1    g224(.A(G143), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n409), .A2(new_n326), .A3(G143), .A4(G214), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT89), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n416));
  INV_X1    g230(.A(G131), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR4_X1   g233(.A1(new_n414), .A2(KEYINPUT89), .A3(new_n416), .A4(new_n417), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n408), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G113), .B(G122), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n238), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n414), .A2(G131), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n417), .A3(new_n413), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n406), .A2(KEYINPUT16), .ZN(new_n428));
  OR3_X1    g242(.A1(new_n226), .A2(KEYINPUT16), .A3(G140), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(G146), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n196), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n414), .A2(KEYINPUT17), .A3(G131), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n427), .A2(new_n430), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n421), .A2(new_n423), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n406), .B(KEYINPUT19), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n200), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n424), .A2(new_n426), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n430), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n423), .B1(new_n421), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n405), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n445), .B(new_n405), .C1(new_n435), .C2(new_n440), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n423), .B1(new_n421), .B2(new_n434), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n314), .B1(new_n435), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G475), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G952), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  NAND2_X1  g267(.A1(G234), .A2(G237), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(G902), .A3(G953), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(G898), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(G119), .A2(G128), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n250), .A2(new_n251), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(G128), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT24), .B(G110), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(KEYINPUT23), .ZN(new_n467));
  AOI21_X1  g281(.A(G128), .B1(new_n250), .B2(new_n251), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n468), .A2(KEYINPUT23), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT74), .B(G110), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n407), .A3(new_n430), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(G110), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n432), .A2(new_n430), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n464), .A2(new_n465), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT75), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT75), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT22), .B(G137), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n326), .A2(G221), .A3(G234), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n484), .B(KEYINPUT76), .Z(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n473), .A2(new_n477), .A3(new_n484), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G217), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(G234), .B2(new_n314), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n486), .A2(new_n487), .A3(new_n314), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n496), .B2(new_n490), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n499));
  INV_X1    g313(.A(new_n347), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(new_n343), .ZN(new_n501));
  MUX2_X1   g315(.A(new_n501), .B(new_n348), .S(new_n417), .Z(new_n502));
  NAND2_X1  g316(.A1(new_n355), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n349), .B1(new_n234), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n295), .A2(new_n504), .A3(new_n205), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n291), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n357), .A2(new_n358), .A3(new_n502), .ZN(new_n509));
  INV_X1    g323(.A(new_n291), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n234), .A2(new_n349), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n512), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n409), .A2(new_n326), .A3(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n499), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n520), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n512), .A2(new_n515), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n514), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n508), .B2(new_n512), .ZN(new_n526));
  OAI211_X1 g340(.A(KEYINPUT73), .B(new_n522), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n507), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n509), .A2(KEYINPUT30), .A3(new_n511), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n291), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n512), .A2(new_n534), .A3(new_n520), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n512), .B2(new_n520), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n537), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n539), .A2(KEYINPUT31), .A3(new_n533), .A4(new_n535), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n528), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G472), .A2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT32), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n509), .A2(new_n511), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n291), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n515), .B1(new_n548), .B2(new_n512), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n524), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n522), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(G902), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n513), .A2(new_n514), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n520), .A3(new_n523), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n533), .A2(new_n512), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n522), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n557), .A3(new_n551), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n542), .A2(new_n546), .B1(new_n559), .B2(G472), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n521), .A2(new_n527), .B1(new_n538), .B2(new_n540), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n545), .B1(new_n561), .B2(new_n544), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n498), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G122), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G116), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n257), .A2(G122), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n245), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n411), .B2(G128), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n219), .A2(KEYINPUT91), .A3(G143), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n411), .A2(G128), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n342), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G134), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n569), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n257), .A2(G122), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n579), .B(new_n566), .C1(new_n580), .C2(KEYINPUT14), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n564), .A2(G116), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT14), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n582), .B1(new_n583), .B2(new_n565), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT94), .B1(new_n566), .B2(KEYINPUT14), .ZN(new_n585));
  OAI211_X1 g399(.A(G107), .B(new_n581), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n566), .B1(new_n580), .B2(KEYINPUT14), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n591), .A2(KEYINPUT95), .A3(G107), .A4(new_n581), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n578), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n322), .A2(new_n489), .A3(G953), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT13), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n574), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n411), .A2(KEYINPUT13), .A3(G128), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n573), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI22_X1  g413(.A1(KEYINPUT92), .A2(new_n575), .B1(new_n599), .B2(G134), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n245), .B1(new_n565), .B2(new_n566), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(KEYINPUT90), .A3(new_n567), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n604));
  INV_X1    g418(.A(new_n567), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n604), .B1(new_n605), .B2(new_n601), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n600), .B(new_n607), .C1(KEYINPUT92), .C2(new_n575), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n594), .A2(new_n595), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n595), .B1(new_n594), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n314), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT96), .ZN(new_n612));
  INV_X1    g426(.A(G478), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(KEYINPUT15), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(new_n314), .C1(new_n609), .C2(new_n610), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n614), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n314), .B(new_n618), .C1(new_n609), .C2(new_n610), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n404), .A2(new_n461), .A3(new_n563), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  OAI21_X1  g440(.A(G472), .B1(new_n561), .B2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n542), .A2(new_n543), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n323), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n393), .A2(KEYINPUT81), .A3(new_n366), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT81), .B1(new_n393), .B2(new_n366), .ZN(new_n632));
  OAI21_X1  g446(.A(G469), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n364), .B1(new_n371), .B2(new_n373), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n328), .ZN(new_n635));
  INV_X1    g449(.A(new_n398), .ZN(new_n636));
  AOI21_X1  g450(.A(G902), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n400), .B1(new_n637), .B2(new_n324), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n630), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n629), .A2(new_n639), .A3(new_n497), .ZN(new_n640));
  INV_X1    g454(.A(new_n293), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n278), .B1(new_n298), .B2(new_n299), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(KEYINPUT87), .ZN(new_n643));
  AOI21_X1  g457(.A(G902), .B1(new_n643), .B2(new_n279), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n316), .B1(new_n644), .B2(new_n313), .ZN(new_n645));
  INV_X1    g459(.A(new_n319), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n187), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n612), .A2(new_n613), .A3(new_n616), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT98), .B(KEYINPUT33), .Z(new_n649));
  OR3_X1    g463(.A1(new_n609), .A2(new_n610), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n609), .B2(new_n610), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n650), .A2(G478), .A3(new_n314), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n451), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n647), .A2(new_n460), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n640), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT34), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  INV_X1    g474(.A(new_n460), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n318), .A2(new_n319), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n441), .A2(new_n443), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n444), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n441), .A2(KEYINPUT99), .A3(new_n443), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n450), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n624), .A2(new_n667), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n661), .A2(new_n662), .A3(new_n187), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n640), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT100), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT35), .B(G107), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NAND2_X1  g488(.A1(new_n496), .A2(new_n490), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n479), .A2(new_n481), .ZN(new_n676));
  OR3_X1    g490(.A1(new_n676), .A2(KEYINPUT36), .A3(new_n485), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n676), .B1(KEYINPUT36), .B2(new_n485), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n491), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n628), .A2(new_n627), .A3(new_n681), .A4(new_n624), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n404), .A2(new_n461), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT101), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT37), .B(G110), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  NAND2_X1  g500(.A1(new_n542), .A2(new_n546), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n559), .A2(G472), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n562), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n496), .A2(new_n490), .B1(new_n491), .B2(new_n679), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n456), .B1(new_n458), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n450), .B(new_n693), .C1(new_n665), .C2(new_n666), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n690), .A2(new_n624), .A3(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n639), .A2(new_n689), .A3(new_n695), .A4(new_n320), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  NAND2_X1  g511(.A1(new_n623), .A2(new_n451), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n681), .A2(new_n188), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n318), .B2(new_n319), .ZN(new_n701));
  INV_X1    g515(.A(new_n700), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n662), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n699), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n539), .A2(new_n533), .A3(new_n535), .ZN(new_n705));
  INV_X1    g519(.A(new_n512), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n522), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(G472), .B1(new_n709), .B2(G902), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n562), .A2(new_n687), .A3(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT103), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT103), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n704), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(new_n692), .B(KEYINPUT39), .Z(new_n715));
  NAND2_X1  g529(.A1(new_n639), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n639), .A2(KEYINPUT104), .A3(new_n715), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n714), .B1(new_n720), .B2(KEYINPUT40), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT40), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n718), .B2(new_n719), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n411), .ZN(G45));
  INV_X1    g539(.A(new_n655), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n693), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n690), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n639), .A2(new_n320), .A3(new_n689), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AOI21_X1  g544(.A(new_n398), .B1(new_n634), .B2(new_n328), .ZN(new_n731));
  OAI21_X1  g545(.A(G469), .B1(new_n731), .B2(G902), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n323), .A3(new_n399), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n656), .A2(new_n563), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND3_X1  g551(.A1(new_n563), .A2(new_n669), .A3(new_n734), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  NOR2_X1   g553(.A1(new_n647), .A2(new_n733), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n690), .A2(new_n623), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n461), .A3(new_n689), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NAND2_X1  g557(.A1(new_n698), .A2(KEYINPUT106), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n623), .A2(new_n745), .A3(new_n451), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT107), .B1(new_n647), .B2(new_n747), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n444), .A2(new_n446), .B1(G475), .B2(new_n449), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n619), .B(KEYINPUT97), .ZN(new_n750));
  AOI211_X1 g564(.A(KEYINPUT106), .B(new_n749), .C1(new_n750), .C2(new_n617), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n745), .B1(new_n623), .B2(new_n451), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n320), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT28), .B1(new_n706), .B2(new_n707), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n520), .B1(new_n757), .B2(new_n523), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n541), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n543), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n758), .B1(new_n538), .B2(new_n540), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n763), .B2(new_n544), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n627), .A2(new_n761), .A3(new_n497), .A4(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n732), .A2(new_n661), .A3(new_n399), .A4(new_n323), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n756), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT108), .B(G122), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G24));
  AND3_X1   g584(.A1(new_n627), .A2(new_n761), .A3(new_n764), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n740), .A3(new_n728), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  NAND2_X1  g587(.A1(new_n562), .A2(new_n687), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n774), .A2(new_n775), .B1(G472), .B2(new_n559), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n562), .A2(new_n687), .A3(KEYINPUT111), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n498), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n630), .A2(new_n188), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n318), .A2(new_n319), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n366), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n374), .B2(new_n375), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT109), .A4(new_n368), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n324), .B(new_n781), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT110), .B1(new_n785), .B2(new_n402), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(G469), .A3(new_n366), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n638), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n727), .B(new_n780), .C1(new_n786), .C2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n778), .A2(KEYINPUT42), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT42), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n786), .A2(new_n790), .ZN(new_n794));
  INV_X1    g608(.A(new_n780), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n563), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n793), .B1(new_n796), .B2(new_n727), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(KEYINPUT112), .B(G131), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G33));
  NOR2_X1   g614(.A1(new_n624), .A2(new_n694), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n794), .A2(new_n563), .A3(new_n801), .A4(new_n795), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  NOR2_X1   g617(.A1(new_n662), .A2(new_n188), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n451), .B1(new_n648), .B2(new_n653), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n805), .A2(KEYINPUT114), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n806), .B1(new_n805), .B2(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n629), .A2(new_n809), .A3(new_n690), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n804), .B1(new_n810), .B2(KEYINPUT44), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(KEYINPUT44), .B2(new_n810), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n787), .A2(KEYINPUT45), .A3(new_n366), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT45), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n378), .A2(new_n817), .A3(new_n394), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(G469), .ZN(new_n819));
  OAI211_X1 g633(.A(KEYINPUT46), .B(new_n401), .C1(new_n816), .C2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT46), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n819), .B1(new_n814), .B2(new_n815), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n400), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n399), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n812), .A2(new_n824), .A3(new_n323), .A4(new_n715), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G137), .ZN(G39));
  INV_X1    g640(.A(new_n804), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n827), .A2(new_n689), .A3(new_n497), .A4(new_n727), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(KEYINPUT47), .A3(new_n323), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT47), .B1(new_n824), .B2(new_n323), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g646(.A(KEYINPUT115), .B(G140), .Z(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(G42));
  NAND2_X1  g648(.A1(new_n452), .A2(new_n326), .ZN(new_n835));
  INV_X1    g649(.A(new_n831), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n732), .A2(new_n399), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n323), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n829), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT120), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n836), .A2(new_n842), .A3(new_n829), .A4(new_n839), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n765), .A2(new_n809), .A3(new_n455), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n827), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n841), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n703), .A2(new_n701), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n850), .A2(new_n187), .A3(new_n733), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n848), .B1(new_n851), .B2(new_n844), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT50), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n809), .A2(new_n455), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n627), .A2(new_n681), .A3(new_n761), .A4(new_n764), .ZN(new_n855));
  INV_X1    g669(.A(new_n837), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n795), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n712), .A2(new_n713), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n498), .A2(new_n837), .A3(new_n780), .A4(new_n455), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n654), .A2(new_n451), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n853), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n852), .A2(KEYINPUT50), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n847), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(new_n726), .A3(new_n859), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n844), .A2(new_n740), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n453), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(KEYINPUT121), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n778), .A2(new_n856), .A3(new_n795), .A4(new_n854), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT48), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n862), .A2(new_n864), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n830), .A2(new_n831), .A3(new_n838), .ZN(new_n876));
  INV_X1    g690(.A(new_n846), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n874), .B1(new_n878), .B2(new_n863), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n866), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n681), .A2(new_n630), .A3(new_n692), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n785), .A2(new_n402), .A3(KEYINPUT110), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n789), .B1(new_n638), .B2(new_n788), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n711), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n320), .A2(new_n753), .A3(new_n754), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n754), .B1(new_n320), .B2(new_n753), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n696), .A2(new_n772), .A3(new_n729), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n882), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n756), .A2(new_n711), .A3(new_n794), .A4(new_n883), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n404), .B(new_n689), .C1(new_n695), .C2(new_n728), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT52), .A4(new_n772), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n897), .B(new_n882), .C1(new_n890), .C2(new_n891), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n893), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n625), .A2(new_n768), .A3(new_n683), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n655), .B1(new_n624), .B2(new_n451), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n320), .A2(new_n661), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(new_n629), .A3(new_n639), .A4(new_n497), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n735), .A2(new_n903), .A3(new_n738), .A4(new_n742), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n727), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n794), .A2(new_n855), .A3(new_n906), .A4(new_n795), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n694), .B1(new_n633), .B2(new_n638), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n689), .A3(new_n741), .A4(new_n795), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n802), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AND4_X1   g725(.A1(KEYINPUT53), .A2(new_n905), .A3(new_n798), .A4(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT52), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n890), .B2(new_n891), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n896), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n910), .B1(new_n792), .B2(new_n797), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n905), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n899), .A2(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n916), .A2(new_n905), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT53), .B1(new_n922), .B2(new_n899), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n917), .A2(new_n918), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n921), .B1(new_n925), .B2(new_n920), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n835), .B1(new_n880), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n497), .A2(new_n779), .A3(new_n805), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(KEYINPUT49), .B2(new_n837), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT116), .Z(new_n930));
  INV_X1    g744(.A(KEYINPUT49), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n850), .B1(new_n931), .B2(new_n856), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n858), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n927), .A2(new_n933), .ZN(G75));
  NOR2_X1   g748(.A1(new_n919), .A2(new_n314), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(G210), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n312), .ZN(new_n939));
  XOR2_X1   g753(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n936), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n936), .B2(new_n937), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n326), .A2(G952), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(G51));
  XNOR2_X1  g759(.A(new_n919), .B(KEYINPUT54), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n400), .B(KEYINPUT57), .Z(new_n947));
  OAI22_X1  g761(.A1(new_n946), .A2(new_n947), .B1(new_n396), .B2(new_n398), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n935), .A2(new_n822), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(G54));
  OR2_X1    g764(.A1(new_n435), .A2(new_n440), .ZN(new_n951));
  NAND2_X1  g765(.A1(KEYINPUT58), .A2(G475), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT123), .Z(new_n953));
  AND3_X1   g767(.A1(new_n935), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n935), .B2(new_n953), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n944), .ZN(G60));
  INV_X1    g770(.A(new_n944), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n650), .A2(new_n652), .ZN(new_n958));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT59), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n957), .B1(new_n946), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n958), .B1(new_n926), .B2(new_n960), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT60), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT53), .B1(new_n922), .B2(new_n915), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n905), .A2(new_n798), .A3(KEYINPUT53), .A4(new_n911), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n898), .A2(new_n896), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n893), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n944), .B1(new_n972), .B2(new_n488), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n912), .A2(new_n899), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n917), .A2(new_n918), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n966), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n974), .B1(new_n977), .B2(new_n679), .ZN(new_n978));
  INV_X1    g792(.A(new_n679), .ZN(new_n979));
  NOR4_X1   g793(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n979), .A4(new_n966), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n973), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n973), .B(KEYINPUT61), .C1(new_n978), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(G66));
  OAI21_X1  g799(.A(G953), .B1(new_n191), .B2(new_n459), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n905), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n938), .B1(G898), .B2(new_n326), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  NAND2_X1  g803(.A1(new_n531), .A2(new_n532), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(new_n436), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(G900), .B2(G953), .ZN(new_n992));
  INV_X1    g806(.A(new_n891), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n993), .A2(new_n802), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n825), .A2(new_n798), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n778), .A2(new_n756), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n824), .A2(new_n323), .A3(new_n996), .A4(new_n715), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n995), .A2(new_n832), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n992), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n993), .B1(new_n721), .B2(new_n723), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n563), .A2(new_n804), .A3(new_n901), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n720), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1006), .B(new_n993), .C1(new_n721), .C2(new_n723), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1003), .A2(new_n1005), .A3(new_n825), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n828), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n836), .B2(new_n829), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n326), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n991), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1001), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n326), .B1(G227), .B2(G900), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT126), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1013), .B(new_n1015), .ZN(G72));
  AOI21_X1  g830(.A(new_n522), .B1(new_n533), .B2(new_n512), .ZN(new_n1017));
  INV_X1    g831(.A(new_n905), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1008), .A2(new_n1010), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT63), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1017), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n999), .A2(new_n998), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n825), .A2(new_n798), .A3(new_n994), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1023), .A2(new_n1010), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1021), .B1(new_n1025), .B2(new_n905), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n533), .A2(new_n512), .A3(new_n522), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n957), .B(new_n1022), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1029));
  INV_X1    g843(.A(new_n925), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1021), .B1(new_n705), .B2(new_n557), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1029), .B(new_n1031), .C1(new_n923), .C2(new_n924), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1028), .A2(new_n1035), .ZN(G57));
endmodule


