//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT82), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n192), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n198), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G107), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n205), .A2(KEYINPUT3), .A3(G104), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT3), .B1(new_n205), .B2(G104), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n202), .B(new_n204), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT83), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n205), .B2(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G104), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n203), .A2(KEYINPUT83), .A3(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n201), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n214), .A2(new_n208), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n196), .A2(G146), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n194), .B2(G143), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n198), .B1(new_n221), .B2(new_n199), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n215), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n224), .B(new_n225), .C1(new_n226), .C2(G137), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT11), .A3(G134), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(G137), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(G134), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n224), .B1(new_n232), .B2(new_n225), .ZN(new_n233));
  OAI21_X1  g047(.A(G131), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n229), .A2(new_n230), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n226), .A2(G137), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(new_n236), .B2(KEYINPUT11), .ZN(new_n237));
  INV_X1    g051(.A(G131), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .A4(new_n227), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n223), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT12), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G101), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT0), .A4(G128), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n221), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT69), .B(new_n246), .C1(new_n221), .C2(new_n247), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n243), .A2(new_n252), .A3(G101), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n245), .A2(new_n250), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n222), .A2(KEYINPUT70), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(new_n198), .C1(new_n221), .C2(new_n199), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n255), .A2(new_n216), .A3(KEYINPUT10), .A4(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n240), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT10), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n215), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n254), .A2(new_n258), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n223), .A2(new_n263), .A3(new_n240), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n242), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT84), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n242), .A2(new_n262), .A3(KEYINPUT84), .A4(new_n264), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n191), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n191), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n254), .A2(new_n258), .A3(new_n261), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n240), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n272), .B2(new_n262), .ZN(new_n273));
  OAI21_X1  g087(.A(G469), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n262), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n270), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n242), .A2(new_n262), .A3(new_n191), .A4(new_n264), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT85), .ZN(new_n278));
  INV_X1    g092(.A(new_n198), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n219), .A2(new_n220), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n195), .ZN(new_n281));
  INV_X1    g095(.A(new_n199), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n214), .A2(new_n208), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI221_X4 g099(.A(KEYINPUT12), .B1(new_n239), .B2(new_n234), .C1(new_n285), .C2(new_n215), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n263), .B1(new_n223), .B2(new_n240), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n191), .A4(new_n262), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n276), .A2(new_n278), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n274), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT101), .ZN(new_n301));
  OAI21_X1  g115(.A(G214), .B1(G237), .B2(G902), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n302), .B(KEYINPUT86), .Z(new_n303));
  NAND2_X1  g117(.A1(new_n248), .A2(G125), .ZN(new_n304));
  INV_X1    g118(.A(G125), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n305), .B(new_n198), .C1(new_n221), .C2(new_n199), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n187), .A2(G224), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(KEYINPUT89), .A2(KEYINPUT6), .ZN(new_n311));
  INV_X1    g125(.A(G116), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G119), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G116), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT2), .B(G113), .Z(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n214), .A2(new_n318), .A3(new_n208), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT5), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT87), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT5), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT68), .B1(new_n313), .B2(new_n315), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n314), .A2(G116), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n312), .A2(G119), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n324), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n313), .A2(new_n321), .A3(new_n323), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT88), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n313), .A2(new_n321), .A3(new_n323), .A4(KEYINPUT88), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(G113), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n319), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT2), .B(G113), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n325), .A2(new_n337), .A3(new_n329), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n318), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n245), .A2(new_n339), .A3(new_n253), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n336), .A2(new_n340), .A3(new_n342), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n311), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n342), .B1(new_n336), .B2(new_n340), .ZN(new_n347));
  INV_X1    g161(.A(new_n311), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n310), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n304), .A2(KEYINPUT7), .A3(new_n308), .A4(new_n306), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n304), .A2(new_n306), .B1(KEYINPUT7), .B2(new_n308), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT91), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n355), .A2(new_n333), .A3(G113), .A4(new_n334), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n319), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n318), .B1(new_n335), .B2(new_n330), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n357), .A2(new_n358), .B1(new_n359), .B2(new_n284), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n319), .A2(KEYINPUT90), .A3(new_n356), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n342), .B(KEYINPUT8), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n352), .B(new_n354), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G210), .B1(G237), .B2(G902), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n350), .A2(new_n293), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n366), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n336), .A2(new_n340), .A3(new_n342), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n348), .B1(new_n369), .B2(new_n347), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n344), .A2(new_n311), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n309), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n247), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n281), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n305), .B1(new_n374), .B2(new_n246), .ZN(new_n375));
  INV_X1    g189(.A(new_n306), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT7), .ZN(new_n377));
  INV_X1    g191(.A(new_n308), .ZN(new_n378));
  OAI22_X1  g192(.A1(new_n375), .A2(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT91), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n353), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n380), .A2(new_n345), .A3(new_n382), .A4(new_n351), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n364), .B1(new_n360), .B2(new_n361), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n293), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n368), .B1(new_n372), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n303), .B1(new_n367), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G478), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(KEYINPUT15), .ZN(new_n389));
  INV_X1    g203(.A(G122), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT14), .B1(new_n390), .B2(G116), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(G116), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT97), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n312), .A2(G122), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n394), .A2(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT97), .ZN(new_n397));
  OAI21_X1  g211(.A(G107), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n390), .A2(G116), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n394), .A3(KEYINPUT96), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT96), .B1(new_n399), .B2(new_n394), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n205), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G128), .B(G143), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n226), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n398), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT13), .B1(new_n192), .B2(G143), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(new_n226), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(new_n404), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n401), .A2(new_n205), .A3(new_n402), .ZN(new_n410));
  INV_X1    g224(.A(new_n402), .ZN(new_n411));
  AOI21_X1  g225(.A(G107), .B1(new_n411), .B2(new_n400), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G217), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n298), .A2(new_n414), .A3(G953), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n406), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT98), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n406), .A2(new_n413), .A3(new_n418), .A4(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n406), .A2(new_n413), .ZN(new_n420));
  INV_X1    g234(.A(new_n415), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n417), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n293), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT99), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n389), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(G234), .A2(G237), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n427), .A2(G952), .A3(new_n187), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(G902), .A3(G953), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n429), .B(KEYINPUT100), .Z(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(G898), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n389), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n423), .A2(KEYINPUT99), .A3(new_n293), .A4(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n426), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n196), .ZN(new_n438));
  NOR2_X1   g252(.A1(G237), .A2(G953), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(G214), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G237), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n187), .A3(G214), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT92), .A2(G143), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G131), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT17), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n443), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n438), .A2(G214), .A3(new_n439), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n238), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT94), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n448), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT17), .A3(G131), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT16), .ZN(new_n454));
  INV_X1    g268(.A(G140), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(G125), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(G125), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n305), .A2(G140), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n456), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n194), .ZN(new_n461));
  OAI211_X1 g275(.A(G146), .B(new_n456), .C1(new_n459), .C2(new_n454), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n453), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n445), .A2(new_n464), .A3(new_n446), .A4(new_n449), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G113), .B(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n203), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT18), .A2(G131), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n447), .A2(new_n448), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT93), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT78), .B1(new_n459), .B2(G146), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT78), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n457), .A2(new_n458), .A3(new_n473), .A4(new_n194), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n459), .A2(G146), .ZN(new_n476));
  INV_X1    g290(.A(new_n469), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n452), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n466), .A2(new_n468), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT95), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n466), .A2(new_n479), .A3(new_n482), .A4(new_n468), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n445), .A2(new_n449), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n459), .B(KEYINPUT19), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n485), .B(new_n462), .C1(G146), .C2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n468), .B1(new_n479), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n491));
  NOR2_X1   g305(.A1(G475), .A2(G902), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n488), .B1(new_n481), .B2(new_n483), .ZN(new_n494));
  INV_X1    g308(.A(new_n492), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT20), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n468), .B1(new_n466), .B2(new_n479), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n481), .B2(new_n483), .ZN(new_n499));
  OAI21_X1  g313(.A(G475), .B1(new_n499), .B2(G902), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n436), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n300), .A2(new_n301), .A3(new_n387), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n297), .A2(new_n387), .A3(new_n299), .ZN(new_n503));
  INV_X1    g317(.A(new_n498), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n484), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n293), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n493), .A2(new_n496), .B1(new_n506), .B2(G475), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n436), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT101), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n314), .A2(G128), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n192), .A2(G119), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT75), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT75), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT24), .B(G110), .Z(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n514), .A2(KEYINPUT76), .A3(new_n516), .A4(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT77), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n314), .B2(G128), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT23), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT23), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n512), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n511), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n461), .A2(new_n462), .B1(G110), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n528), .A2(G110), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n517), .B1(new_n514), .B2(new_n516), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n462), .B(new_n475), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT79), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT22), .B(G137), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n530), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n530), .B2(new_n533), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT25), .A3(new_n293), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n530), .A2(new_n533), .ZN(new_n542));
  INV_X1    g356(.A(new_n537), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n530), .A2(new_n533), .A3(new_n537), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n293), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n414), .B1(G234), .B2(new_n293), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n552));
  INV_X1    g366(.A(new_n540), .ZN(new_n553));
  INV_X1    g367(.A(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n293), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT80), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n554), .B1(new_n541), .B2(new_n548), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT81), .B1(new_n560), .B2(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n232), .A2(new_n230), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G131), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n255), .A2(new_n239), .A3(new_n564), .A4(new_n257), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n240), .A2(new_n250), .A3(new_n251), .ZN(new_n566));
  INV_X1    g380(.A(new_n339), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n439), .A2(G210), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT27), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT26), .B(G101), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT30), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT65), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n248), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT65), .B(new_n246), .C1(new_n221), .C2(new_n247), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n240), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT67), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n222), .A2(new_n239), .A3(new_n564), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n240), .A2(new_n576), .A3(KEYINPUT67), .A4(new_n577), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT30), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n574), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n573), .B1(new_n585), .B2(new_n339), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n582), .A2(new_n581), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n239), .A2(new_n234), .B1(new_n248), .B2(new_n575), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT67), .B1(new_n591), .B2(new_n577), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n584), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n574), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n339), .ZN(new_n595));
  INV_X1    g409(.A(new_n573), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n588), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT72), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT31), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n595), .B2(new_n596), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n589), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n572), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT28), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n339), .B1(new_n590), .B2(new_n592), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n604), .B2(new_n568), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n565), .A2(new_n566), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT73), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n339), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT73), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT28), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n602), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT74), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT74), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(new_n602), .C1(new_n605), .C2(new_n610), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n601), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(G472), .A2(G902), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT32), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n606), .A2(new_n339), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n603), .B1(new_n621), .B2(new_n568), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n610), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT29), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n602), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n568), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n585), .B2(new_n339), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n624), .B1(new_n628), .B2(new_n572), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n605), .A2(new_n610), .A3(new_n602), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n616), .A2(new_n620), .B1(G472), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n597), .B(KEYINPUT72), .C1(new_n586), .C2(new_n599), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n633), .A2(new_n589), .B1(new_n612), .B2(new_n614), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n619), .B1(new_n634), .B2(new_n618), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n562), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n510), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  AOI21_X1  g452(.A(G902), .B1(new_n601), .B2(new_n615), .ZN(new_n639));
  INV_X1    g453(.A(G472), .ZN(new_n640));
  OAI22_X1  g454(.A1(new_n639), .A2(new_n640), .B1(new_n618), .B2(new_n634), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n297), .A2(new_n561), .A3(new_n559), .A4(new_n299), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n422), .A2(KEYINPUT33), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n416), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n416), .A2(new_n645), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT102), .B(KEYINPUT33), .Z(new_n649));
  AOI22_X1  g463(.A1(new_n647), .A2(new_n648), .B1(new_n423), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n388), .A2(G902), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n650), .A2(new_n651), .B1(new_n388), .B2(new_n424), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n497), .B2(new_n500), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n303), .B(new_n432), .C1(new_n367), .C2(new_n386), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n643), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n496), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g474(.A(KEYINPUT104), .B(KEYINPUT20), .C1(new_n494), .C2(new_n495), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n495), .B1(new_n484), .B2(new_n489), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n662), .B1(new_n663), .B2(new_n491), .ZN(new_n664));
  NOR4_X1   g478(.A1(new_n494), .A2(KEYINPUT105), .A3(KEYINPUT20), .A4(new_n495), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n660), .B(new_n661), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n426), .A2(new_n435), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(new_n500), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n666), .A2(new_n654), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n643), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  INV_X1    g486(.A(new_n641), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n543), .A2(KEYINPUT36), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(new_n542), .Z(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n556), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n560), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n673), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT106), .B1(new_n641), .B2(new_n678), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n510), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT107), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n428), .B1(new_n430), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n666), .A2(new_n668), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n666), .A2(KEYINPUT108), .A3(new_n668), .A4(new_n688), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n297), .A2(new_n679), .A3(new_n387), .A4(new_n299), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n631), .A2(G472), .ZN(new_n696));
  INV_X1    g510(.A(new_n620), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n696), .B1(new_n634), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT32), .B1(new_n616), .B2(new_n617), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n695), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n192), .ZN(G30));
  XOR2_X1   g516(.A(new_n687), .B(KEYINPUT39), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n300), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT111), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n494), .A2(KEYINPUT20), .A3(new_n495), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n500), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n667), .ZN(new_n711));
  INV_X1    g525(.A(new_n628), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n572), .ZN(new_n713));
  INV_X1    g527(.A(new_n621), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n627), .ZN(new_n715));
  AOI21_X1  g529(.A(G902), .B1(new_n715), .B2(new_n602), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n640), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n616), .B2(new_n620), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n711), .B1(new_n718), .B2(new_n635), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n367), .A2(new_n386), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT109), .B(KEYINPUT38), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT110), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n303), .A3(new_n679), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n706), .A2(new_n707), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n196), .ZN(G45));
  NOR3_X1   g541(.A1(new_n507), .A2(new_n652), .A3(new_n687), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n695), .B(new_n728), .C1(new_n698), .C2(new_n699), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT112), .B(G146), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G48));
  NAND2_X1  g545(.A1(new_n291), .A2(new_n293), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n299), .A3(new_n294), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n562), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n655), .B(new_n735), .C1(new_n698), .C2(new_n699), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  OAI211_X1 g552(.A(new_n669), .B(new_n735), .C1(new_n699), .C2(new_n698), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  INV_X1    g554(.A(new_n303), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n720), .A2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n734), .A2(new_n742), .A3(new_n678), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n743), .B(new_n501), .C1(new_n698), .C2(new_n699), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  NAND3_X1  g559(.A1(new_n710), .A2(new_n387), .A3(new_n667), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n733), .A2(new_n299), .A3(new_n294), .A4(new_n433), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n560), .A2(new_n557), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n602), .B1(new_n610), .B2(new_n622), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n601), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n617), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT113), .B(G472), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n634), .B2(G902), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n748), .A2(new_n749), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  AND4_X1   g570(.A1(new_n387), .A2(new_n733), .A3(new_n299), .A4(new_n294), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n728), .A3(new_n679), .ZN(new_n758));
  INV_X1    g572(.A(new_n753), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n752), .B1(new_n639), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n305), .ZN(G27));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  INV_X1    g577(.A(new_n749), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n632), .B2(new_n635), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n274), .A2(KEYINPUT114), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n767), .B(G469), .C1(new_n269), .C2(new_n273), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n766), .A2(new_n294), .A3(new_n296), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n299), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n720), .A2(new_n303), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n728), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n763), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n632), .A2(new_n635), .ZN(new_n775));
  INV_X1    g589(.A(new_n653), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(KEYINPUT42), .A3(new_n687), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n552), .B1(new_n551), .B2(new_n558), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n560), .A2(KEYINPUT81), .A3(new_n557), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n769), .A2(new_n780), .A3(new_n771), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n775), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT115), .B1(new_n774), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n749), .B1(new_n698), .B2(new_n699), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT42), .B1(new_n784), .B2(new_n772), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n775), .A2(new_n777), .A3(new_n781), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n238), .ZN(G33));
  NAND4_X1  g604(.A1(new_n775), .A2(new_n781), .A3(new_n691), .A4(new_n692), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  OR3_X1    g606(.A1(new_n269), .A2(KEYINPUT45), .A3(new_n273), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT45), .B1(new_n269), .B2(new_n273), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(G469), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n296), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n296), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n294), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(new_n299), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n703), .ZN(new_n802));
  INV_X1    g616(.A(new_n652), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n507), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT116), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT43), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n641), .A3(new_n679), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n367), .A2(new_n386), .A3(new_n741), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n806), .A2(KEYINPUT44), .A3(new_n641), .A4(new_n679), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n802), .A2(new_n809), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G137), .ZN(G39));
  XNOR2_X1  g628(.A(new_n801), .B(KEYINPUT47), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n728), .A2(new_n562), .A3(new_n811), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n775), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NAND4_X1  g633(.A1(new_n723), .A2(new_n749), .A3(new_n741), .A4(new_n299), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n804), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n718), .A2(new_n635), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n733), .A2(new_n294), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT49), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n667), .B(new_n500), .C1(new_n708), .C2(new_n709), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n654), .B1(new_n828), .B2(new_n653), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n641), .A2(new_n829), .A3(new_n642), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n510), .B2(new_n636), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(new_n682), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n297), .A2(new_n679), .A3(new_n299), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n500), .A2(new_n435), .A3(new_n426), .A4(new_n688), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n810), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n666), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n666), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n775), .A2(new_n833), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n618), .B1(new_n601), .B2(new_n750), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n616), .A2(new_n293), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n842), .B2(new_n753), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n769), .A2(new_n771), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n679), .A4(new_n728), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n791), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n739), .A2(new_n736), .A3(new_n744), .A4(new_n755), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n832), .A2(new_n848), .A3(new_n783), .A4(new_n788), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n691), .A2(new_n692), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n694), .B1(new_n632), .B2(new_n635), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n761), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n560), .A2(new_n677), .A3(new_n770), .A4(new_n687), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n769), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n742), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n769), .A2(KEYINPUT118), .A3(new_n854), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n719), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n852), .A2(new_n853), .A3(new_n729), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n843), .A2(new_n728), .A3(new_n743), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n729), .C1(new_n693), .C2(new_n700), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n857), .A2(new_n719), .A3(new_n858), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT52), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n826), .B1(new_n849), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n791), .A2(new_n840), .A3(new_n845), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n736), .A2(new_n739), .A3(new_n744), .A4(new_n755), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n682), .A4(new_n831), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n789), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n860), .A2(new_n864), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT54), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n774), .A2(new_n782), .A3(new_n826), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n871), .A2(new_n832), .A3(new_n848), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n866), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n806), .A2(new_n428), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n734), .A2(new_n810), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT120), .Z(new_n885));
  AND2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n679), .A3(new_n843), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n780), .A3(new_n428), .A4(new_n822), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n888), .A2(new_n710), .A3(new_n803), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n749), .A2(new_n806), .A3(new_n428), .A4(new_n843), .ZN(new_n890));
  AND4_X1   g704(.A1(new_n303), .A2(new_n723), .A3(new_n299), .A4(new_n823), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n890), .A2(KEYINPUT50), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT50), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n887), .B(new_n889), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n811), .ZN(new_n895));
  INV_X1    g709(.A(new_n815), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n823), .A2(new_n770), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n881), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(KEYINPUT121), .B(KEYINPUT48), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n883), .A2(new_n765), .A3(new_n885), .A4(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(G952), .A3(new_n187), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n890), .A2(new_n757), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n776), .B2(new_n888), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n886), .A2(new_n765), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(KEYINPUT48), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n902), .B(new_n904), .C1(new_n905), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n874), .B1(new_n873), .B2(KEYINPUT54), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n894), .A2(new_n898), .A3(new_n881), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n880), .A2(new_n909), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n825), .B1(new_n912), .B2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n187), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n293), .B1(new_n866), .B2(new_n877), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n346), .A2(new_n349), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n309), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n350), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n918), .B2(new_n923), .ZN(G51));
  AOI211_X1 g739(.A(new_n293), .B(new_n795), .C1(new_n866), .C2(new_n877), .ZN(new_n926));
  INV_X1    g740(.A(new_n291), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n870), .B2(new_n871), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n832), .A2(new_n848), .A3(new_n876), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n865), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT54), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n879), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n295), .B(KEYINPUT57), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n926), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n933), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n931), .B2(new_n879), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT122), .B1(new_n938), .B2(new_n927), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n915), .B1(new_n936), .B2(new_n939), .ZN(G54));
  NAND3_X1  g754(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n941), .A2(new_n494), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n494), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n915), .ZN(G60));
  NAND2_X1  g758(.A1(G478), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT59), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n932), .A2(new_n650), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n916), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n880), .B2(new_n910), .ZN(new_n950));
  INV_X1    g764(.A(new_n650), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n928), .B2(new_n930), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n915), .B1(new_n956), .B2(new_n553), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT61), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n676), .B2(new_n956), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI221_X1 g775(.A(new_n957), .B1(new_n958), .B2(KEYINPUT61), .C1(new_n676), .C2(new_n956), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G66));
  INV_X1    g777(.A(new_n431), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n187), .B1(new_n964), .B2(G224), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n832), .A2(new_n868), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n187), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n919), .B1(G898), .B2(new_n187), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n967), .B(new_n968), .Z(G69));
  OR3_X1    g783(.A1(new_n726), .A2(KEYINPUT62), .A3(new_n862), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT62), .B1(new_n726), .B2(new_n862), .ZN(new_n971));
  INV_X1    g785(.A(new_n636), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n811), .B1(new_n828), .B2(new_n653), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n705), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n813), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n970), .A2(new_n818), .A3(new_n971), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n187), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n585), .B(new_n486), .ZN(new_n978));
  XNOR2_X1  g792(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n978), .B(new_n979), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n983));
  NAND2_X1  g797(.A1(G900), .A2(G953), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n784), .A2(new_n746), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n802), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n813), .A2(new_n986), .A3(new_n791), .ZN(new_n987));
  INV_X1    g801(.A(new_n789), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n862), .B1(new_n815), .B2(new_n817), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n980), .B(new_n984), .C1(new_n990), .C2(G953), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n982), .A2(new_n983), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n982), .A2(new_n991), .A3(new_n983), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n976), .B2(new_n966), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n572), .A3(new_n712), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n628), .A2(new_n572), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n873), .B(new_n999), .C1(new_n586), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n712), .A2(new_n572), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n966), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1006), .B1(new_n1008), .B2(new_n999), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT127), .ZN(new_n1010));
  OR3_X1    g824(.A1(new_n1009), .A2(new_n1010), .A3(new_n915), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1010), .B1(new_n1009), .B2(new_n915), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1004), .B1(new_n1011), .B2(new_n1012), .ZN(G57));
endmodule


