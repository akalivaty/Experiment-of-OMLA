//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1192, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT65), .Z(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n203), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT66), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n203), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND3_X1  g0015(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n217), .B2(new_n218), .C1(new_n210), .C2(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n212), .A2(new_n219), .ZN(G361));
  XNOR2_X1  g0020(.A(G238), .B(G244), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(G232), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT2), .B(G226), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(G264), .B(G270), .Z(new_n225));
  XNOR2_X1  g0025(.A(G250), .B(G257), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n224), .B(new_n227), .ZN(G358));
  XOR2_X1   g0028(.A(G68), .B(G77), .Z(new_n229));
  XOR2_X1   g0029(.A(G50), .B(G58), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G87), .B(G97), .Z(new_n232));
  XOR2_X1   g0032(.A(G107), .B(G116), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G351));
  XNOR2_X1  g0035(.A(KEYINPUT67), .B(G1), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n236), .A2(G13), .A3(G20), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(KEYINPUT69), .ZN(new_n239));
  INV_X1    g0039(.A(G33), .ZN(new_n240));
  OAI21_X1  g0040(.A(new_n239), .B1(new_n203), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(G1), .A2(G13), .ZN(new_n242));
  NAND4_X1  g0042(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n236), .A2(G20), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(G50), .A3(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n240), .A2(G20), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT70), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G150), .ZN(new_n253));
  NOR3_X1   g0053(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n254));
  INV_X1    g0054(.A(G20), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n244), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n238), .A2(new_n258), .ZN(new_n259));
  AND3_X1   g0059(.A1(new_n247), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G169), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(new_n265), .A3(G274), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT67), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G1), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(G1), .B(G13), .C1(new_n240), .C2(new_n262), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G226), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n240), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n279), .A2(G223), .B1(new_n282), .B2(G77), .ZN(new_n283));
  INV_X1    g0083(.A(G222), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n275), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n286), .B(new_n287), .C1(new_n280), .C2(new_n281), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n283), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n271), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n274), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n260), .B1(new_n261), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(G179), .B2(new_n292), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G20), .A2(G77), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n252), .A2(KEYINPUT71), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n252), .A2(KEYINPUT71), .ZN(new_n297));
  OR3_X1    g0097(.A1(new_n296), .A2(new_n250), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT15), .B(G87), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n255), .A2(G33), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n295), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n244), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n245), .A2(G77), .A3(new_n246), .ZN(new_n304));
  INV_X1    g0104(.A(G77), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n238), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(G238), .B1(new_n280), .B2(new_n281), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(G1698), .B1(new_n282), .B2(G107), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT3), .B(G33), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(G232), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n271), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  INV_X1    g0118(.A(G244), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n266), .B1(new_n272), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n261), .B1(new_n316), .B2(new_n320), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n307), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n317), .A2(G190), .A3(new_n321), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n302), .A2(new_n244), .B1(new_n305), .B2(new_n238), .ZN(new_n326));
  OAI21_X1  g0126(.A(G200), .B1(new_n316), .B2(new_n320), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n304), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n260), .A2(KEYINPUT9), .B1(new_n292), .B2(G200), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT10), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n247), .A2(new_n257), .A3(new_n259), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT9), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n332), .A2(new_n333), .B1(new_n291), .B2(G190), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n330), .B2(new_n334), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n294), .B(new_n329), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n314), .A2(new_n338), .A3(G20), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n282), .B2(new_n255), .ZN(new_n340));
  OAI21_X1  g0140(.A(G68), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(G58), .B(G68), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(G20), .B1(G159), .B2(new_n252), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n341), .A2(KEYINPUT16), .A3(new_n343), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n244), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n244), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n250), .B1(G20), .B2(new_n236), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n238), .A2(new_n250), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n266), .ZN(new_n353));
  INV_X1    g0153(.A(new_n272), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(G232), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n279), .A2(G226), .ZN(new_n356));
  INV_X1    g0156(.A(G87), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n240), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G223), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n288), .A2(KEYINPUT75), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT75), .B1(new_n288), .B2(new_n359), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n355), .B1(new_n362), .B2(new_n271), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n261), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n318), .B(new_n355), .C1(new_n362), .C2(new_n271), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n352), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT18), .ZN(new_n367));
  INV_X1    g0167(.A(new_n351), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n349), .B1(new_n344), .B2(new_n345), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n347), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n363), .A2(G200), .ZN(new_n371));
  OAI211_X1 g0171(.A(G190), .B(new_n355), .C1(new_n362), .C2(new_n271), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n352), .A2(new_n376), .A3(new_n364), .A4(new_n365), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT17), .A4(new_n372), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n367), .A2(new_n375), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n337), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT74), .ZN(new_n381));
  INV_X1    g0181(.A(G68), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n249), .B2(new_n305), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n244), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT11), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n238), .A2(KEYINPUT12), .A3(new_n382), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT12), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n237), .B2(G68), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n245), .A2(G68), .A3(new_n246), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n385), .B2(new_n386), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT14), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n288), .A2(new_n273), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G232), .A2(G1698), .ZN(new_n399));
  INV_X1    g0199(.A(G97), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n282), .A2(new_n399), .B1(new_n240), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n290), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n270), .A2(G238), .A3(new_n271), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n403), .A2(new_n266), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT13), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n399), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n314), .A2(new_n407), .B1(G33), .B2(G97), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n313), .A2(new_n314), .A3(G226), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n271), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n403), .A2(new_n266), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT13), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n261), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n405), .B1(new_n402), .B2(new_n404), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT13), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n397), .A2(new_n413), .B1(new_n416), .B2(G179), .ZN(new_n417));
  OAI21_X1  g0217(.A(G169), .B1(new_n414), .B2(new_n415), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n396), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n397), .B(G169), .C1(new_n414), .C2(new_n415), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n406), .A2(new_n412), .A3(G179), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n406), .A2(new_n412), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n397), .B1(new_n424), .B2(G169), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n423), .A2(KEYINPUT73), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n395), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G190), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n394), .B1(new_n428), .B2(new_n424), .ZN(new_n429));
  INV_X1    g0229(.A(G200), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n416), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n381), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT73), .B1(new_n423), .B2(new_n425), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n419), .A2(new_n396), .A3(new_n422), .A4(new_n421), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n394), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n437), .A2(new_n432), .A3(KEYINPUT74), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n380), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT76), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n380), .B(KEYINPUT76), .C1(new_n434), .C2(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AND4_X1   g0244(.A1(G45), .A2(new_n267), .A3(new_n269), .A4(G274), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(KEYINPUT80), .A3(new_n271), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n271), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n267), .A2(new_n269), .A3(G45), .A4(G274), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n236), .A2(G45), .ZN(new_n453));
  INV_X1    g0253(.A(new_n446), .ZN(new_n454));
  OAI211_X1 g0254(.A(G264), .B(new_n271), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(G257), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G294), .ZN(new_n457));
  INV_X1    g0257(.A(G250), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n288), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n290), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n452), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n430), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n452), .A2(new_n460), .A3(new_n428), .A4(new_n455), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(KEYINPUT86), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT85), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT25), .ZN(new_n466));
  AOI21_X1  g0266(.A(G107), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n238), .A2(new_n467), .B1(KEYINPUT85), .B2(KEYINPUT25), .ZN(new_n468));
  NOR4_X1   g0268(.A1(new_n237), .A2(new_n465), .A3(new_n466), .A4(G107), .ZN(new_n469));
  INV_X1    g0269(.A(G107), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n236), .A2(G33), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n349), .A2(new_n237), .A3(new_n471), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n468), .A2(new_n469), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT23), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n255), .B2(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n470), .A2(KEYINPUT23), .A3(G20), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n475), .A2(new_n476), .B1(new_n248), .B2(G116), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n255), .B(G87), .C1(new_n280), .C2(new_n281), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n478), .A2(KEYINPUT22), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(KEYINPUT22), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT24), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n473), .B1(new_n485), .B2(new_n244), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n464), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n461), .A2(G179), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n461), .A2(new_n261), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n349), .B1(new_n482), .B2(new_n484), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n473), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT72), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n299), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n245), .A2(new_n495), .A3(new_n471), .ZN(new_n496));
  NAND3_X1  g0296(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n255), .ZN(new_n498));
  NOR4_X1   g0298(.A1(KEYINPUT82), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  NOR2_X1   g0300(.A1(G87), .A2(G97), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(new_n470), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT83), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT19), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n504), .B(new_n505), .C1(new_n301), .C2(new_n400), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n314), .A2(new_n255), .A3(G68), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n301), .B2(new_n400), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT83), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n503), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n244), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n300), .A2(new_n238), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n496), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n286), .A2(new_n287), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n308), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n290), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n458), .B1(new_n236), .B2(G45), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n271), .B1(new_n519), .B2(new_n445), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n318), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT81), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n518), .A2(new_n520), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n261), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n518), .A2(KEYINPUT81), .A3(new_n520), .A4(new_n318), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n513), .A2(new_n523), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(G200), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n349), .A2(new_n237), .A3(new_n471), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G87), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n510), .A2(new_n244), .B1(new_n238), .B2(new_n300), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n518), .A2(G190), .A3(new_n520), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n528), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n493), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(G107), .B1(new_n339), .B2(new_n340), .ZN(new_n536));
  XNOR2_X1  g0336(.A(G97), .B(G107), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT77), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n400), .A2(KEYINPUT6), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n540), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n541), .A2(G20), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n252), .A2(G77), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n536), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n244), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n237), .A2(G97), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n529), .B2(G97), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g0350(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n288), .B2(new_n319), .ZN(new_n552));
  INV_X1    g0352(.A(G283), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n240), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n279), .B2(G250), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT4), .A4(G244), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT79), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n552), .A2(new_n555), .A3(KEYINPUT79), .A4(new_n556), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n290), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G257), .B(new_n271), .C1(new_n453), .C2(new_n454), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n452), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(G190), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n271), .B1(new_n557), .B2(new_n558), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n566), .B2(new_n560), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n550), .B(new_n565), .C1(new_n430), .C2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n561), .A2(new_n318), .A3(new_n564), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n547), .A2(new_n549), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(G169), .C2(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n529), .A2(G116), .ZN(new_n574));
  INV_X1    g0374(.A(G116), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n238), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n554), .ZN(new_n577));
  AOI21_X1  g0377(.A(G20), .B1(new_n240), .B2(G97), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n577), .A2(new_n578), .B1(G20), .B2(new_n575), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n579), .A2(new_n244), .A3(KEYINPUT20), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT20), .B1(new_n579), .B2(new_n244), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n574), .B(new_n576), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n313), .A2(new_n314), .A3(G257), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n314), .A2(G264), .A3(G1698), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n282), .A2(G303), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n290), .ZN(new_n588));
  OAI211_X1 g0388(.A(G270), .B(new_n271), .C1(new_n453), .C2(new_n454), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n452), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G200), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n583), .B(new_n591), .C1(new_n428), .C2(new_n590), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n452), .A2(new_n588), .A3(G179), .A4(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(G169), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n582), .ZN(new_n597));
  XNOR2_X1  g0397(.A(KEYINPUT84), .B(KEYINPUT21), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n583), .B2(new_n594), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n592), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n535), .A2(new_n573), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n444), .A2(new_n601), .ZN(G372));
  OR2_X1    g0402(.A1(new_n335), .A2(new_n336), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n375), .A2(new_n378), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n432), .A2(new_n324), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n427), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n367), .A2(new_n377), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n603), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n294), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT26), .B1(new_n571), .B2(new_n534), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT87), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n525), .A2(new_n613), .A3(new_n521), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n525), .B2(new_n521), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n513), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n571), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n568), .A2(new_n488), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n597), .A2(new_n599), .A3(new_n492), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n533), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n612), .B(new_n616), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n611), .B1(new_n444), .B2(new_n624), .ZN(G369));
  INV_X1    g0425(.A(KEYINPUT27), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n255), .A2(G13), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n236), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT88), .ZN(new_n629));
  INV_X1    g0429(.A(G213), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n626), .B1(new_n236), .B2(new_n627), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT89), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n631), .A2(G343), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n582), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n600), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n597), .A2(new_n599), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n635), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G330), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT90), .ZN(new_n640));
  INV_X1    g0440(.A(new_n634), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n488), .B(new_n492), .C1(new_n486), .C2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n492), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n634), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n597), .A2(new_n599), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n641), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n649), .A2(new_n493), .B1(new_n492), .B2(new_n634), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT91), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n647), .A2(new_n651), .ZN(G399));
  OR3_X1    g0452(.A1(new_n499), .A2(new_n502), .A3(G116), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n213), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(G1), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n218), .B2(new_n657), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT29), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n623), .A2(new_n661), .A3(new_n641), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT92), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n572), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n616), .A2(new_n488), .A3(new_n533), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n568), .A2(new_n571), .A3(KEYINPUT92), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n664), .A2(new_n619), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT93), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n616), .A2(new_n488), .A3(new_n533), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n637), .B2(new_n492), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT93), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n664), .A4(new_n666), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n621), .B1(new_n571), .B2(new_n534), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n533), .A2(KEYINPUT26), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n561), .A2(new_n564), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n261), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n674), .A2(new_n570), .A3(new_n569), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n616), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n668), .A2(new_n672), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n641), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n662), .B1(new_n682), .B2(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n460), .A2(new_n455), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n593), .A2(new_n684), .A3(new_n524), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n567), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(KEYINPUT30), .A3(new_n567), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n461), .A2(new_n318), .A3(new_n524), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n675), .A3(new_n590), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n634), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n695), .B(new_n696), .C1(new_n601), .C2(new_n634), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n683), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n660), .B1(new_n700), .B2(G1), .ZN(G364));
  AOI21_X1  g0501(.A(new_n265), .B1(new_n627), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n656), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n640), .B(new_n705), .C1(G330), .C2(new_n638), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n314), .A2(new_n213), .ZN(new_n707));
  INV_X1    g0507(.A(G355), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(G116), .B2(new_n213), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n231), .A2(G45), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n655), .A2(new_n314), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n218), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n263), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n709), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G13), .A2(G33), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n242), .B1(G20), .B2(new_n261), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n704), .B1(new_n715), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n255), .A2(new_n318), .A3(new_n430), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT94), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G190), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n318), .A2(new_n430), .A3(KEYINPUT95), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT95), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G179), .B2(G200), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n428), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n255), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n725), .A2(G68), .B1(G97), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n724), .A2(new_n428), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n255), .A2(G190), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n726), .B2(new_n728), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G159), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n732), .B1(new_n258), .B2(new_n734), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n255), .A2(new_n318), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G190), .A3(new_n430), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G58), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n736), .A2(new_n318), .A3(G200), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n282), .B1(new_n748), .B2(G77), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n255), .A2(G179), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n750), .A2(new_n428), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n752), .A2(G87), .B1(new_n754), .B2(G107), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n743), .A2(new_n747), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(KEYINPUT33), .B(G317), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G326), .A2(new_n733), .B1(new_n725), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G294), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(new_n730), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n752), .A2(G303), .B1(new_n754), .B2(G283), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n314), .B1(new_n746), .B2(G322), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n737), .A2(G329), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n748), .A2(G311), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n742), .A2(new_n756), .B1(new_n760), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n722), .B1(new_n766), .B2(new_n719), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n718), .B(KEYINPUT97), .Z(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n638), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n706), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(G396));
  NAND2_X1  g0571(.A1(new_n634), .A2(new_n307), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n328), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n324), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n324), .A2(new_n634), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT101), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT101), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n774), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n624), .B2(new_n634), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n618), .A2(new_n619), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n622), .B1(new_n784), .B2(new_n571), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n612), .A2(new_n616), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n641), .B(new_n781), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n704), .B1(new_n788), .B2(new_n698), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n698), .B2(new_n788), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n719), .A2(new_n716), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n704), .B1(new_n792), .B2(G77), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n357), .A2(new_n753), .B1(new_n751), .B2(new_n470), .ZN(new_n794));
  INV_X1    g0594(.A(new_n748), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n282), .B1(new_n759), .B2(new_n745), .C1(new_n795), .C2(new_n575), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(G311), .C2(new_n737), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n733), .A2(G303), .B1(G97), .B2(new_n731), .ZN(new_n798));
  INV_X1    g0598(.A(new_n725), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n798), .C1(new_n553), .C2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n748), .A2(G159), .B1(new_n746), .B2(G143), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  INV_X1    g0603(.A(G150), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(new_n734), .B2(new_n803), .C1(new_n804), .C2(new_n799), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n258), .A2(new_n751), .B1(new_n753), .B2(new_n382), .ZN(new_n808));
  INV_X1    g0608(.A(G58), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n730), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n282), .B1(new_n737), .B2(G132), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n808), .B(new_n810), .C1(KEYINPUT100), .C2(new_n811), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(KEYINPUT100), .B2(new_n811), .C1(new_n805), .C2(new_n806), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n801), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n793), .B1(new_n814), .B2(new_n719), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n717), .B2(new_n781), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n790), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G384));
  NOR2_X1   g0618(.A1(new_n217), .A2(new_n575), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT35), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n823), .B(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(G77), .B1(new_n809), .B2(new_n382), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n826), .A2(new_n218), .B1(G50), .B2(new_n382), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n236), .A2(G13), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n631), .A2(new_n633), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n607), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT39), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n352), .A2(new_n830), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n366), .A2(new_n373), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n379), .A2(new_n352), .A3(new_n830), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT38), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT38), .B1(new_n835), .B2(new_n836), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n832), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT38), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n379), .A2(new_n352), .A3(new_n830), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n834), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n427), .A2(new_n634), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n831), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n787), .A2(new_n776), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n427), .A2(new_n433), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n394), .A2(new_n641), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n845), .A2(new_n837), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT103), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n683), .B2(new_n444), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n661), .B1(new_n681), .B2(new_n641), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n443), .B(KEYINPUT103), .C1(new_n862), .C2(new_n662), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n610), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n859), .B(new_n864), .Z(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n697), .A2(new_n781), .ZN(new_n867));
  INV_X1    g0667(.A(new_n853), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n852), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n854), .A2(KEYINPUT104), .A3(new_n697), .A4(new_n781), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n857), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT40), .B1(new_n838), .B2(new_n839), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n854), .A2(new_n697), .A3(new_n781), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT105), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n873), .B1(new_n845), .B2(new_n837), .ZN(new_n878));
  INV_X1    g0678(.A(new_n867), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n854), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n874), .A2(new_n882), .A3(G330), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n443), .A2(G330), .A3(new_n697), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT106), .Z(new_n886));
  AOI22_X1  g0686(.A1(new_n877), .A2(new_n881), .B1(new_n872), .B2(new_n873), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n887), .A2(new_n443), .A3(new_n697), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n865), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n236), .B2(new_n627), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n886), .A2(new_n865), .A3(new_n888), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n829), .B1(new_n890), .B2(new_n891), .ZN(G367));
  OAI221_X1 g0692(.A(new_n720), .B1(new_n300), .B2(new_n213), .C1(new_n227), .C2(new_n712), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(new_n704), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n641), .B1(new_n530), .B2(new_n531), .ZN(new_n895));
  INV_X1    g0695(.A(new_n616), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n897), .A2(KEYINPUT107), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n616), .A2(new_n533), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n899), .A2(new_n895), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(KEYINPUT107), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n719), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n799), .A2(new_n739), .B1(new_n258), .B2(new_n795), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n904), .A2(KEYINPUT112), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(KEYINPUT112), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n282), .B1(new_n746), .B2(G150), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n907), .B1(new_n809), .B2(new_n751), .C1(new_n305), .C2(new_n753), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(G137), .B2(new_n737), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n733), .A2(G143), .B1(G68), .B2(new_n731), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n905), .A2(new_n906), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n753), .A2(new_n400), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n282), .B1(new_n795), .B2(new_n553), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(G303), .C2(new_n746), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n737), .A2(G317), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT46), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n752), .A2(G116), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n731), .A2(G107), .ZN(new_n920));
  AOI22_X1  g0720(.A1(G294), .A2(new_n725), .B1(new_n733), .B2(G311), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n914), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n911), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT47), .Z(new_n924));
  OAI221_X1 g0724(.A(new_n894), .B1(new_n902), .B2(new_n768), .C1(new_n903), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n664), .B(new_n666), .C1(new_n550), .C2(new_n641), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n617), .A2(new_n634), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n927), .A2(KEYINPUT108), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT108), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n649), .A2(new_n493), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n617), .B1(new_n932), .B2(new_n643), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n634), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n926), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OR4_X1    g0742(.A1(KEYINPUT43), .A2(new_n936), .A3(new_n902), .A4(new_n939), .ZN(new_n943));
  INV_X1    g0743(.A(new_n647), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n931), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT110), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n942), .A2(new_n943), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(new_n945), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n931), .A2(new_n651), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT44), .Z(new_n952));
  NOR2_X1   g0752(.A1(new_n931), .A2(new_n651), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT45), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n944), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n944), .B1(new_n952), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n646), .A2(new_n649), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n933), .B1(new_n959), .B2(KEYINPUT111), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(KEYINPUT111), .B2(new_n959), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n640), .B(new_n961), .Z(new_n962));
  AOI21_X1  g0762(.A(new_n699), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n656), .B(KEYINPUT41), .Z(new_n964));
  OAI21_X1  g0764(.A(new_n702), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n947), .B2(new_n946), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n925), .B1(new_n950), .B2(new_n966), .ZN(G387));
  INV_X1    g0767(.A(new_n962), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n699), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n699), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n656), .A3(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n645), .A2(new_n768), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n711), .B1(new_n224), .B2(new_n263), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n654), .B2(new_n707), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n250), .A2(G50), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT50), .ZN(new_n977));
  AOI21_X1  g0777(.A(G45), .B1(G68), .B2(G77), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n654), .A3(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n975), .A2(new_n979), .B1(new_n470), .B2(new_n655), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n704), .B1(new_n980), .B2(new_n721), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n752), .A2(G77), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n400), .B2(new_n753), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n314), .B1(new_n258), .B2(new_n745), .C1(new_n795), .C2(new_n382), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(G150), .C2(new_n737), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n733), .A2(G159), .B1(new_n495), .B2(new_n731), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(new_n250), .C2(new_n799), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n737), .A2(G326), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n314), .B1(new_n754), .B2(G116), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n730), .A2(new_n553), .B1(new_n759), .B2(new_n751), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n725), .A2(G311), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n748), .A2(G303), .B1(new_n746), .B2(G317), .ZN(new_n992));
  INV_X1    g0792(.A(G322), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n992), .C1(new_n734), .C2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT48), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n995), .B2(new_n994), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT49), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n988), .B(new_n989), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n987), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n981), .B1(new_n1001), .B2(new_n719), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n962), .A2(new_n703), .B1(new_n973), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n972), .A2(new_n1003), .ZN(G393));
  INV_X1    g0804(.A(new_n958), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n656), .B1(new_n1005), .B2(new_n970), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n970), .B2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n931), .A2(new_n718), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n234), .A2(new_n711), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1009), .B(new_n720), .C1(new_n400), .C2(new_n213), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT113), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1012), .A2(new_n1013), .A3(new_n705), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n738), .A2(new_n993), .B1(new_n553), .B2(new_n751), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT115), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n282), .B1(new_n470), .B2(new_n753), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n1016), .B2(new_n1015), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT116), .Z(new_n1019));
  OAI22_X1  g0819(.A1(new_n795), .A2(new_n759), .B1(new_n730), .B2(new_n575), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n733), .A2(G317), .B1(G311), .B2(new_n746), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT52), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1020), .B(new_n1022), .C1(G303), .C2(new_n725), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n314), .B1(new_n751), .B2(new_n382), .C1(new_n357), .C2(new_n753), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G143), .B2(new_n737), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT114), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n730), .A2(new_n305), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n799), .A2(new_n258), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n795), .A2(new_n250), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n733), .A2(G150), .B1(G159), .B2(new_n746), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT51), .Z(new_n1032));
  AOI22_X1  g0832(.A1(new_n1019), .A2(new_n1023), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1008), .B(new_n1014), .C1(new_n903), .C2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1005), .B2(new_n702), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1007), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(G390));
  NAND4_X1  g0837(.A1(new_n854), .A2(G330), .A3(new_n697), .A4(new_n781), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n681), .A2(new_n641), .A3(new_n781), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n869), .B1(new_n1039), .B2(new_n776), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n849), .B1(new_n845), .B2(new_n837), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(KEYINPUT117), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT117), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n679), .B1(new_n667), .B2(KEYINPUT93), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n634), .B1(new_n1045), .B2(new_n672), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n775), .B1(new_n1046), .B2(new_n781), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1044), .B(new_n1041), .C1(new_n1047), .C2(new_n869), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n849), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n855), .A2(new_n1050), .B1(new_n840), .B2(new_n846), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1038), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1038), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1054), .B(new_n1051), .C1(new_n1043), .C2(new_n1048), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT118), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n863), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n623), .A2(new_n661), .A3(new_n641), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1046), .B2(new_n661), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT103), .B1(new_n1060), .B2(new_n443), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n611), .B(new_n884), .C1(new_n1058), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n851), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n869), .B1(new_n698), .B2(new_n782), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1063), .B1(new_n1038), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1038), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n1047), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1057), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1047), .A2(new_n1038), .A3(new_n1064), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1066), .B2(new_n1063), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n864), .A2(KEYINPUT118), .A3(new_n884), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1072), .A2(KEYINPUT119), .A3(new_n1056), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT119), .B1(new_n1072), .B2(new_n1056), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n656), .B1(new_n1056), .B2(new_n1072), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n792), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n705), .B1(new_n1076), .B2(new_n250), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n752), .A2(G150), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT53), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n733), .A2(G128), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT54), .B(G143), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n748), .A2(new_n1082), .B1(new_n746), .B2(G132), .ZN(new_n1083));
  INV_X1    g0883(.A(G125), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1080), .B(new_n1083), .C1(new_n1084), .C2(new_n738), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1079), .B(new_n1085), .C1(G159), .C2(new_n731), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n314), .B1(new_n753), .B2(new_n258), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n799), .A2(new_n803), .B1(KEYINPUT120), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(KEYINPUT120), .B2(new_n1087), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n382), .A2(new_n753), .B1(new_n751), .B2(new_n357), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n282), .B1(new_n575), .B2(new_n745), .C1(new_n795), .C2(new_n400), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(G294), .C2(new_n737), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n734), .A2(new_n553), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1027), .B(new_n1093), .C1(G107), .C2(new_n725), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1086), .A2(new_n1089), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1077), .B1(new_n903), .B2(new_n1095), .C1(new_n848), .C2(new_n717), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1056), .B2(new_n703), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1075), .A2(new_n1098), .ZN(G378));
  NAND2_X1  g0899(.A1(new_n603), .A2(new_n294), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n830), .A2(new_n332), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT55), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1100), .B(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1104));
  XOR2_X1   g0904(.A(new_n1103), .B(new_n1104), .Z(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n717), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n748), .A2(G137), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n746), .A2(G128), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n752), .A2(new_n1082), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n734), .A2(new_n1084), .B1(new_n730), .B2(new_n804), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G132), .C2(new_n725), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1113), .A2(KEYINPUT59), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(KEYINPUT59), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n240), .B(new_n262), .C1(new_n753), .C2(new_n739), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G124), .B2(new_n737), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n725), .A2(G97), .B1(G68), .B2(new_n731), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n575), .B2(new_n734), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n314), .A2(G41), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G107), .B2(new_n746), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1123), .B(new_n982), .C1(new_n809), .C2(new_n753), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n300), .A2(new_n795), .B1(new_n738), .B2(new_n553), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1120), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT58), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1122), .B(new_n258), .C1(G33), .C2(G41), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1126), .A2(KEYINPUT58), .ZN(new_n1129));
  AND4_X1   g0929(.A1(new_n1118), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n704), .B1(G50), .B2(new_n792), .C1(new_n1130), .C2(new_n903), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1106), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n883), .A2(new_n1105), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1105), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n887), .A2(G330), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n859), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT122), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1134), .A2(new_n1136), .A3(new_n859), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n859), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT122), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1133), .B1(new_n1145), .B2(new_n702), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT57), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1072), .A2(new_n1056), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT119), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1072), .A2(new_n1056), .A3(KEYINPUT119), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1062), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1147), .B1(new_n1152), .B2(new_n1145), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1062), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1147), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n657), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1146), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(G375));
  NAND2_X1  g0959(.A1(new_n869), .A2(new_n716), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n704), .B1(new_n792), .B2(G68), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n752), .A2(G97), .B1(new_n754), .B2(G77), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n314), .B1(new_n748), .B2(G107), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n737), .A2(G303), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n746), .A2(G283), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n725), .A2(G116), .B1(new_n495), .B2(new_n731), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n759), .B2(new_n734), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n733), .A2(G132), .B1(G50), .B2(new_n731), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n799), .B2(new_n1081), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n752), .A2(G159), .B1(new_n754), .B2(G58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n282), .B1(new_n748), .B2(G150), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n737), .A2(G128), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n746), .A2(G137), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1166), .A2(new_n1168), .B1(new_n1170), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1161), .B1(new_n1176), .B2(new_n719), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1070), .A2(new_n703), .B1(new_n1160), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n964), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1178), .B1(new_n1072), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT123), .Z(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(G381));
  OR2_X1    g0984(.A1(G387), .A2(G390), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(G378), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n1158), .A4(new_n1183), .ZN(G407));
  NOR2_X1   g0990(.A1(new_n630), .A2(G343), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1158), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(G407), .A2(G213), .A3(new_n1192), .ZN(G409));
  NOR3_X1   g0993(.A1(new_n1152), .A2(new_n964), .A3(new_n1145), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1141), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n703), .B1(new_n1195), .B2(new_n1143), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1133), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT125), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1189), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1146), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(KEYINPUT124), .A3(G378), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT124), .B1(new_n1158), .B2(G378), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1199), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1191), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1068), .A2(new_n1071), .A3(KEYINPUT60), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1208), .A2(new_n1179), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT60), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n656), .B1(new_n1179), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(G384), .A3(new_n1178), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1178), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n817), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(KEYINPUT126), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1191), .A2(G2897), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT126), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1214), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1216), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1219), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT61), .B1(new_n1207), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1205), .A2(new_n1206), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT63), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(G393), .B(new_n770), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G387), .A2(G390), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1185), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1185), .B2(new_n1234), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1156), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n656), .B1(new_n1152), .B2(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1155), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G378), .B(new_n1201), .C1(new_n1240), .C2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1202), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1191), .B1(new_n1246), .B2(new_n1199), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1228), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1227), .A2(new_n1231), .A3(new_n1238), .A4(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1247), .B2(new_n1225), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT62), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1229), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1247), .A2(KEYINPUT62), .A3(new_n1228), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1251), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT127), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1237), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(KEYINPUT127), .A3(new_n1235), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1249), .B1(new_n1255), .B2(new_n1260), .ZN(G405));
  OAI21_X1  g1061(.A(new_n1246), .B1(G378), .B2(new_n1158), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(new_n1228), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1228), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1238), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(new_n1238), .A3(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(G402));
endmodule


