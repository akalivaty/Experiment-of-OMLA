//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1131, new_n1132, new_n1134;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT66), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT67), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n464), .A2(G136), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(G162));
  NAND2_X1  g056(.A1(new_n476), .A2(G126), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n465), .A2(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n463), .B2(new_n484), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n461), .A2(new_n462), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n465), .A2(G138), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n482), .A2(new_n485), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  NAND2_X1  g067(.A1(G50), .A2(G543), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT5), .A2(G543), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G88), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n504), .B(KEYINPUT70), .C1(new_n500), .C2(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(G166));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT72), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n501), .A2(new_n515), .A3(new_n502), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n514), .A2(new_n516), .A3(G51), .A4(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT71), .B1(new_n494), .B2(new_n495), .ZN(new_n522));
  AND2_X1   g097(.A1(G63), .A2(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT73), .B(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n503), .A2(new_n505), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n517), .A2(new_n524), .A3(new_n528), .A4(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n518), .A2(new_n520), .B1(new_n501), .B2(new_n502), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(new_n529), .B1(new_n527), .B2(new_n526), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n535), .A2(KEYINPUT74), .A3(new_n517), .A4(new_n524), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(G168));
  AND2_X1   g112(.A1(new_n521), .A2(new_n522), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n500), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n534), .A2(G90), .ZN(new_n542));
  INV_X1    g117(.A(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n503), .B2(KEYINPUT72), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(new_n516), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n541), .A2(new_n547), .ZN(G171));
  NAND3_X1  g123(.A1(new_n521), .A2(new_n522), .A3(G56), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n500), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n534), .A2(G81), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n514), .A2(new_n516), .A3(G43), .A4(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT76), .Z(G188));
  NAND3_X1  g137(.A1(new_n503), .A2(new_n505), .A3(G91), .ZN(new_n563));
  INV_X1    g138(.A(G78), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n505), .B2(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n563), .B1(new_n566), .B2(new_n500), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n514), .A2(new_n516), .A3(G53), .A4(G543), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(G299));
  OR2_X1    g147(.A1(new_n541), .A2(new_n547), .ZN(G301));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n533), .A2(new_n574), .A3(new_n536), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n574), .B1(new_n533), .B2(new_n536), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND3_X1  g153(.A1(new_n544), .A2(G49), .A3(new_n516), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n534), .A2(G87), .ZN(new_n580));
  AOI21_X1  g155(.A(G74), .B1(new_n521), .B2(new_n522), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n500), .C2(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n500), .ZN(new_n584));
  NAND2_X1  g159(.A1(G48), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n496), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(new_n503), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n538), .A2(G60), .ZN(new_n590));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n500), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n534), .A2(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n545), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n496), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n514), .A2(new_n516), .A3(G54), .A4(G543), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT10), .B1(new_n534), .B2(G92), .ZN(new_n604));
  AND4_X1   g179(.A1(KEYINPUT10), .A2(new_n503), .A3(new_n505), .A4(G92), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(G868), .B2(new_n607), .ZN(G284));
  OAI21_X1  g183(.A(new_n598), .B1(G868), .B2(new_n607), .ZN(G321));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g185(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n607), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(KEYINPUT78), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(KEYINPUT78), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n616), .B(new_n617), .C1(G868), .C2(new_n555), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g194(.A1(G123), .A2(new_n476), .B1(new_n464), .B2(G135), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n621), .A2(new_n465), .A3(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n465), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT80), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n488), .A2(new_n466), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n627), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n639), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT82), .ZN(G401));
  XNOR2_X1  g224(.A(G2072), .B(G2078), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT17), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT83), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n652), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n657), .B(new_n654), .C1(new_n650), .C2(new_n652), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n650), .A3(new_n652), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n674), .C1(new_n666), .C2(new_n673), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  XOR2_X1   g251(.A(G1981), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(new_n681), .ZN(G229));
  NOR2_X1   g257(.A1(G29), .A2(G35), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G162), .B2(G29), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT29), .B(G2090), .Z(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n687));
  NAND2_X1  g262(.A1(G103), .A2(G2104), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(G2105), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n465), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n690));
  AOI22_X1  g265(.A1(new_n464), .A2(G139), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI22_X1  g266(.A1(new_n488), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n465), .B2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G33), .B(new_n693), .S(G29), .Z(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G2072), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G26), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n464), .A2(G140), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n476), .A2(G128), .ZN(new_n701));
  OR2_X1    g276(.A1(G104), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n697), .ZN(new_n706));
  INV_X1    g281(.A(G2067), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n697), .A2(G32), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT95), .B(KEYINPUT26), .ZN(new_n710));
  AND3_X1   g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n712), .A2(new_n713), .B1(G105), .B2(new_n466), .ZN(new_n714));
  AOI22_X1  g289(.A1(G129), .A2(new_n476), .B1(new_n464), .B2(G141), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(new_n697), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT96), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n695), .A2(new_n708), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n555), .A2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G16), .B2(G19), .ZN(new_n724));
  INV_X1    g299(.A(G1341), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G5), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G171), .B2(new_n727), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n726), .B1(G1961), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n491), .A2(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n697), .A2(G27), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G34), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n697), .B1(new_n736), .B2(G34), .ZN(new_n738));
  OAI22_X1  g313(.A1(new_n472), .A2(new_n697), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n734), .A2(G2078), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  INV_X1    g316(.A(new_n739), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n741), .A2(new_n733), .B1(new_n742), .B2(G2084), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(new_n743), .C1(new_n725), .C2(new_n724), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n686), .A2(new_n722), .A3(new_n730), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n729), .A2(G1961), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT98), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT31), .B(G11), .Z(new_n748));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n697), .B1(new_n749), .B2(G28), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(KEYINPUT97), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(KEYINPUT97), .B1(new_n749), .B2(G28), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n625), .B2(new_n697), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n727), .A2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G168), .B2(new_n727), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n755), .B1(new_n757), .B2(G1966), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n747), .B(new_n758), .C1(G1966), .C2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT99), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n727), .A2(G4), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n607), .B2(new_n727), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT92), .B(G1348), .Z(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT93), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n762), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n727), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT100), .B(G1956), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n745), .A2(new_n760), .A3(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n759), .A2(KEYINPUT99), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n727), .A2(G22), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT91), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n727), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1971), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n727), .A2(G6), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n583), .A2(new_n500), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n503), .B2(new_n587), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n780), .B1(new_n782), .B2(new_n727), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XOR2_X1   g359(.A(new_n783), .B(new_n784), .Z(new_n785));
  MUX2_X1   g360(.A(G23), .B(G288), .S(G16), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT33), .B(G1976), .Z(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n779), .A2(new_n785), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n697), .A2(G25), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT87), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n476), .A2(G119), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT88), .Z(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n797));
  INV_X1    g372(.A(G107), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G2105), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n464), .B2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n794), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT35), .B(G1991), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT89), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n802), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n727), .A2(G24), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n596), .A2(KEYINPUT90), .ZN(new_n807));
  OAI21_X1  g382(.A(G16), .B1(new_n596), .B2(KEYINPUT90), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n805), .B1(G1986), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G1986), .B2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n790), .A2(new_n791), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n792), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT36), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(KEYINPUT36), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n775), .B1(new_n814), .B2(new_n815), .ZN(G311));
  INV_X1    g391(.A(G311), .ZN(G150));
  NAND3_X1  g392(.A1(new_n521), .A2(new_n522), .A3(G67), .ZN(new_n818));
  INV_X1    g393(.A(G80), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n543), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G651), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n534), .A2(G93), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n514), .A2(new_n516), .A3(G55), .A4(G543), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT101), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT101), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n607), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  INV_X1    g405(.A(new_n555), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n555), .B(new_n821), .C1(new_n825), .C2(new_n824), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n830), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n838));
  AOI21_X1  g413(.A(G860), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n835), .A2(new_n836), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT103), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n828), .B1(new_n840), .B2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(KEYINPUT106), .B(G37), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n801), .B(new_n629), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n693), .A2(KEYINPUT104), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n717), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n491), .B(new_n704), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n464), .A2(G142), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n465), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT105), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n476), .A2(new_n855), .A3(G130), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n476), .B2(G130), .ZN(new_n857));
  OAI221_X1 g432(.A(new_n852), .B1(new_n853), .B2(new_n854), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n851), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n850), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n625), .B(new_n472), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n848), .A2(new_n859), .A3(new_n849), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n863), .B1(new_n861), .B2(new_n864), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n844), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT9), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n544), .A2(new_n871), .A3(G53), .A4(new_n516), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n567), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n606), .B1(new_n873), .B2(KEYINPUT107), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT107), .ZN(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(G299), .A2(new_n875), .A3(new_n606), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n869), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n869), .A3(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n834), .B(new_n614), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n877), .A2(KEYINPUT108), .A3(new_n878), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT108), .B1(new_n877), .B2(new_n878), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n889));
  XNOR2_X1  g464(.A(G166), .B(G288), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n596), .B(new_n782), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n884), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n889), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n892), .B1(new_n889), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(G868), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n826), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(G868), .B2(new_n898), .ZN(G295));
  OAI21_X1  g474(.A(new_n897), .B1(G868), .B2(new_n898), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n832), .A2(new_n833), .ZN(new_n903));
  NAND2_X1  g478(.A1(G168), .A2(KEYINPUT77), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n533), .A2(new_n574), .A3(new_n536), .ZN(new_n905));
  AOI21_X1  g480(.A(G301), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(G171), .A2(G168), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(G171), .B1(new_n575), .B2(new_n576), .ZN(new_n909));
  OR2_X1    g484(.A1(G171), .A2(G168), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n834), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n882), .A2(new_n902), .A3(new_n908), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n911), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n877), .A2(new_n869), .A3(new_n878), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n914), .A2(new_n879), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT110), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n877), .A2(new_n878), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n908), .B2(new_n911), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n912), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n892), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  XOR2_X1   g497(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n923));
  INV_X1    g498(.A(new_n917), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n909), .A2(new_n834), .A3(new_n910), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n834), .B1(new_n909), .B2(new_n910), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n927), .B(KEYINPUT110), .C1(new_n915), .C2(new_n913), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(new_n892), .A3(new_n912), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n892), .B1(new_n928), .B2(new_n912), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n880), .A2(KEYINPUT111), .A3(new_n881), .ZN(new_n932));
  OR3_X1    g507(.A1(new_n917), .A2(KEYINPUT111), .A3(KEYINPUT41), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n913), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI22_X1  g509(.A1(new_n925), .A2(new_n926), .B1(new_n885), .B2(new_n886), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n892), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n844), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n901), .B1(new_n930), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n923), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n931), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n921), .A2(new_n922), .A3(new_n929), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(new_n901), .ZN(G397));
  XOR2_X1   g519(.A(KEYINPUT112), .B(G1384), .Z(new_n945));
  AOI21_X1  g520(.A(KEYINPUT45), .B1(new_n491), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  OR3_X1    g525(.A1(new_n950), .A2(G1986), .A3(G290), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(G1986), .A3(G290), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT113), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n801), .B(new_n803), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n704), .B(new_n707), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n717), .A2(G1996), .ZN(new_n957));
  INV_X1    g532(.A(G1996), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n716), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n950), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n491), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n948), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n491), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n741), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT126), .B(KEYINPUT53), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n948), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n491), .A2(new_n973), .A3(new_n965), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1961), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n970), .A2(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n948), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n978), .A2(KEYINPUT53), .A3(new_n741), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT127), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n969), .A4(new_n947), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n969), .A2(new_n978), .A3(KEYINPUT53), .A4(new_n741), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT127), .B1(new_n982), .B2(new_n946), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(G171), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT125), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n491), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n968), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n989), .B2(G2078), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n968), .A2(KEYINPUT125), .A3(new_n741), .A4(new_n988), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(KEYINPUT53), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(G301), .B1(new_n992), .B2(new_n977), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n964), .B1(new_n986), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n533), .A2(G8), .A3(new_n536), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n972), .A2(new_n735), .A3(new_n974), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(G1966), .B1(new_n968), .B2(new_n988), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(G8), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT51), .B1(new_n996), .B2(KEYINPUT124), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1001), .A2(new_n995), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n1001), .B2(new_n995), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n985), .A2(G171), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n992), .A2(G301), .A3(new_n977), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(KEYINPUT54), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n509), .A2(G8), .A3(new_n510), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT55), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n972), .A2(new_n974), .ZN(new_n1011));
  INV_X1    g586(.A(G2090), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n491), .A2(new_n965), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n978), .B(new_n969), .C1(new_n1013), .C2(KEYINPUT45), .ZN(new_n1014));
  INV_X1    g589(.A(G1971), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1011), .A2(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n1013), .B2(new_n978), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(G288), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G288), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(KEYINPUT114), .A3(G1976), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  OAI21_X1  g601(.A(G1981), .B1(new_n781), .B2(KEYINPUT115), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n782), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n584), .B(new_n588), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(KEYINPUT49), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n782), .A2(new_n1027), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1031), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1036), .A3(new_n1019), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1021), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .A4(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1026), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n972), .A2(new_n1012), .A3(new_n974), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1017), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1010), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1018), .A2(new_n1040), .A3(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n994), .A2(new_n1005), .A3(new_n1008), .A4(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1013), .A2(new_n978), .A3(KEYINPUT119), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n966), .B2(new_n948), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT58), .B(G1341), .Z(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(G1996), .B2(new_n1014), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n555), .A2(KEYINPUT121), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(KEYINPUT59), .A3(new_n1054), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT56), .B(G2072), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n1011), .A2(G1956), .B1(new_n1014), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n872), .A2(new_n870), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT57), .B1(new_n1062), .B2(KEYINPUT118), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(new_n873), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT61), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1058), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1014), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1068), .A2(new_n1059), .B1(new_n975), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1064), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1067), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n975), .A2(new_n763), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1076), .B(KEYINPUT60), .C1(new_n1077), .C2(G2067), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(KEYINPUT123), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(KEYINPUT123), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n607), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(KEYINPUT123), .A3(new_n606), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1076), .B1(new_n1077), .B2(G2067), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1075), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1084), .A2(new_n607), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1070), .B1(new_n1089), .B2(new_n1071), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1064), .A2(KEYINPUT120), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1072), .A2(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1047), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1043), .B(new_n1010), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1095), .A2(new_n993), .A3(new_n1040), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1040), .A2(new_n1044), .A3(new_n1043), .ZN(new_n1100));
  NOR2_X1   g675(.A1(G305), .A2(G1981), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT116), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G288), .A2(G1976), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1037), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1019), .B1(new_n1104), .B2(KEYINPUT117), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1106), .B(new_n1102), .C1(new_n1037), .C2(new_n1103), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1100), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1001), .A2(G286), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1018), .A2(new_n1109), .A3(new_n1040), .A4(new_n1045), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1095), .A2(KEYINPUT63), .A3(new_n1040), .A4(new_n1109), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1099), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n963), .B1(new_n1093), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n949), .A2(new_n958), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT46), .Z(new_n1118));
  AOI21_X1  g693(.A(new_n950), .B1(new_n956), .B2(new_n717), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT47), .Z(new_n1121));
  INV_X1    g696(.A(KEYINPUT48), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n962), .B1(new_n1122), .B2(new_n951), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1122), .B2(new_n951), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n796), .A2(new_n800), .A3(new_n803), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n960), .A2(new_n1125), .B1(G2067), .B2(new_n704), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n949), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1121), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1116), .A2(new_n1128), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g704(.A1(G401), .A2(G229), .A3(new_n459), .A4(G227), .ZN(new_n1131));
  NAND2_X1  g705(.A1(new_n1131), .A2(new_n867), .ZN(new_n1132));
  NOR2_X1   g706(.A1(new_n943), .A2(new_n1132), .ZN(G308));
  AND2_X1   g707(.A1(new_n942), .A2(new_n940), .ZN(new_n1134));
  OAI211_X1 g708(.A(new_n867), .B(new_n1131), .C1(new_n1134), .C2(new_n941), .ZN(G225));
endmodule


