

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U323 ( .A(n383), .B(n332), .ZN(n333) );
  BUF_X1 U324 ( .A(n464), .Z(n547) );
  XNOR2_X1 U325 ( .A(n334), .B(n333), .ZN(n390) );
  INV_X1 U326 ( .A(KEYINPUT101), .ZN(n471) );
  INV_X1 U327 ( .A(G92GAT), .ZN(n319) );
  XNOR2_X1 U328 ( .A(n471), .B(KEYINPUT25), .ZN(n472) );
  XNOR2_X1 U329 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U330 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U331 ( .A(n365), .B(n321), .ZN(n323) );
  XNOR2_X1 U332 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n398) );
  INV_X1 U333 ( .A(KEYINPUT55), .ZN(n455) );
  XNOR2_X1 U334 ( .A(n399), .B(n398), .ZN(n544) );
  XNOR2_X1 U335 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U336 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U337 ( .A(n310), .B(n309), .ZN(n312) );
  XNOR2_X1 U338 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U339 ( .A(G43GAT), .ZN(n495) );
  XNOR2_X1 U340 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U341 ( .A(n495), .B(KEYINPUT40), .ZN(n496) );
  XNOR2_X1 U342 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n497), .B(n496), .ZN(G1330GAT) );
  XNOR2_X1 U344 ( .A(G134GAT), .B(G127GAT), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n291), .B(KEYINPUT0), .ZN(n424) );
  XOR2_X1 U346 ( .A(n424), .B(G120GAT), .Z(n296) );
  XOR2_X1 U347 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U348 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U349 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U350 ( .A(KEYINPUT19), .B(n294), .ZN(n414) );
  XOR2_X1 U351 ( .A(G113GAT), .B(n414), .Z(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n310) );
  XOR2_X1 U353 ( .A(KEYINPUT86), .B(KEYINPUT82), .Z(n298) );
  XNOR2_X1 U354 ( .A(KEYINPUT84), .B(G71GAT), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U356 ( .A(G176GAT), .B(KEYINPUT80), .Z(n300) );
  XNOR2_X1 U357 ( .A(KEYINPUT83), .B(KEYINPUT81), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n308) );
  XOR2_X1 U360 ( .A(KEYINPUT20), .B(G15GAT), .Z(n304) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G43GAT), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U363 ( .A(G99GAT), .B(G190GAT), .Z(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n464) );
  INV_X1 U367 ( .A(KEYINPUT69), .ZN(n313) );
  NAND2_X1 U368 ( .A1(n313), .A2(G85GAT), .ZN(n316) );
  INV_X1 U369 ( .A(G85GAT), .ZN(n314) );
  NAND2_X1 U370 ( .A1(n314), .A2(KEYINPUT69), .ZN(n315) );
  NAND2_X1 U371 ( .A1(n316), .A2(n315), .ZN(n318) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G106GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n365) );
  NAND2_X1 U374 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  INV_X1 U375 ( .A(KEYINPUT9), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U377 ( .A(G190GAT), .B(G218GAT), .Z(n408) );
  XNOR2_X1 U378 ( .A(KEYINPUT70), .B(n408), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n334) );
  XOR2_X1 U380 ( .A(G29GAT), .B(KEYINPUT8), .Z(n327) );
  XNOR2_X1 U381 ( .A(G43GAT), .B(G36GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U383 ( .A(G50GAT), .B(KEYINPUT7), .Z(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n383) );
  XOR2_X1 U385 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n331) );
  XNOR2_X1 U386 ( .A(G134GAT), .B(G162GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U388 ( .A(KEYINPUT36), .B(n390), .ZN(n487) );
  XOR2_X1 U389 ( .A(KEYINPUT12), .B(KEYINPUT77), .Z(n336) );
  XNOR2_X1 U390 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n356) );
  XOR2_X1 U392 ( .A(KEYINPUT71), .B(G64GAT), .Z(n338) );
  XNOR2_X1 U393 ( .A(G1GAT), .B(G8GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U395 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n340) );
  XNOR2_X1 U396 ( .A(KEYINPUT72), .B(KEYINPUT15), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U398 ( .A(n342), .B(n341), .Z(n354) );
  XNOR2_X1 U399 ( .A(G22GAT), .B(G15GAT), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n343), .B(KEYINPUT66), .ZN(n374) );
  XOR2_X1 U401 ( .A(n374), .B(KEYINPUT14), .Z(n345) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n352) );
  XOR2_X1 U404 ( .A(G57GAT), .B(G211GAT), .Z(n347) );
  XNOR2_X1 U405 ( .A(G127GAT), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U407 ( .A(G71GAT), .B(KEYINPUT13), .Z(n369) );
  XOR2_X1 U408 ( .A(n348), .B(n369), .Z(n350) );
  XNOR2_X1 U409 ( .A(G183GAT), .B(G155GAT), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n498) );
  INV_X1 U414 ( .A(n498), .ZN(n589) );
  NAND2_X1 U415 ( .A1(n487), .A2(n589), .ZN(n358) );
  XOR2_X1 U416 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n359), .B(KEYINPUT112), .ZN(n388) );
  XOR2_X1 U419 ( .A(G204GAT), .B(G78GAT), .Z(n449) );
  XOR2_X1 U420 ( .A(KEYINPUT31), .B(KEYINPUT68), .Z(n361) );
  NAND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n363) );
  INV_X1 U423 ( .A(KEYINPUT33), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n367) );
  XNOR2_X1 U425 ( .A(G176GAT), .B(G92GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n364), .B(G64GAT), .ZN(n406) );
  XNOR2_X1 U427 ( .A(n365), .B(n406), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n368), .B(KEYINPUT32), .ZN(n371) );
  XOR2_X1 U430 ( .A(G148GAT), .B(n369), .Z(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n449), .B(n372), .ZN(n373) );
  XOR2_X1 U433 ( .A(G120GAT), .B(G57GAT), .Z(n425) );
  XNOR2_X1 U434 ( .A(n373), .B(n425), .ZN(n585) );
  INV_X1 U435 ( .A(n585), .ZN(n490) );
  XOR2_X1 U436 ( .A(n374), .B(KEYINPUT65), .Z(n376) );
  NAND2_X1 U437 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U439 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n378) );
  XNOR2_X1 U440 ( .A(G197GAT), .B(G141GAT), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U442 ( .A(n380), .B(n379), .Z(n382) );
  XOR2_X1 U443 ( .A(G113GAT), .B(G1GAT), .Z(n421) );
  XOR2_X1 U444 ( .A(G169GAT), .B(G8GAT), .Z(n409) );
  XNOR2_X1 U445 ( .A(n421), .B(n409), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U447 ( .A(n384), .B(n383), .Z(n385) );
  XOR2_X1 U448 ( .A(n385), .B(KEYINPUT67), .Z(n571) );
  INV_X1 U449 ( .A(n571), .ZN(n386) );
  AND2_X1 U450 ( .A1(n490), .A2(n386), .ZN(n387) );
  AND2_X1 U451 ( .A1(n388), .A2(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(n389), .B(KEYINPUT113), .Z(n397) );
  INV_X1 U453 ( .A(KEYINPUT41), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n391), .B(n585), .ZN(n522) );
  NAND2_X1 U455 ( .A1(n522), .A2(n385), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n392), .B(KEYINPUT46), .ZN(n393) );
  NAND2_X1 U457 ( .A1(n393), .A2(n498), .ZN(n394) );
  NOR2_X1 U458 ( .A1(n390), .A2(n394), .ZN(n395) );
  XOR2_X1 U459 ( .A(KEYINPUT47), .B(n395), .Z(n396) );
  NOR2_X1 U460 ( .A1(n397), .A2(n396), .ZN(n399) );
  XOR2_X1 U461 ( .A(KEYINPUT96), .B(KEYINPUT71), .Z(n401) );
  XNOR2_X1 U462 ( .A(G36GAT), .B(G204GAT), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n413) );
  XOR2_X1 U464 ( .A(G211GAT), .B(KEYINPUT87), .Z(n403) );
  XNOR2_X1 U465 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n446) );
  XOR2_X1 U467 ( .A(n446), .B(KEYINPUT95), .Z(n405) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U471 ( .A(n409), .B(n408), .Z(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n416) );
  INV_X1 U474 ( .A(n414), .ZN(n415) );
  XOR2_X1 U475 ( .A(n416), .B(n415), .Z(n469) );
  BUF_X1 U476 ( .A(n469), .Z(n537) );
  NOR2_X1 U477 ( .A1(n544), .A2(n537), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n417), .B(KEYINPUT54), .ZN(n441) );
  XOR2_X1 U479 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n419) );
  XNOR2_X1 U480 ( .A(KEYINPUT90), .B(KEYINPUT4), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U482 ( .A(n420), .B(G85GAT), .Z(n423) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n429) );
  XOR2_X1 U485 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U488 ( .A(n429), .B(n428), .Z(n440) );
  XOR2_X1 U489 ( .A(G148GAT), .B(G155GAT), .Z(n431) );
  XNOR2_X1 U490 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U492 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n433) );
  XNOR2_X1 U493 ( .A(G162GAT), .B(KEYINPUT88), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n435), .B(n434), .Z(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n437) );
  XNOR2_X1 U497 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n445), .B(n438), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n476) );
  XNOR2_X1 U501 ( .A(KEYINPUT94), .B(n476), .ZN(n535) );
  NAND2_X1 U502 ( .A1(n441), .A2(n535), .ZN(n580) );
  XOR2_X1 U503 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n443) );
  XNOR2_X1 U504 ( .A(G50GAT), .B(G22GAT), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n454) );
  XOR2_X1 U507 ( .A(KEYINPUT23), .B(n446), .Z(n448) );
  NAND2_X1 U508 ( .A1(G228GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X1 U510 ( .A(n450), .B(n449), .Z(n452) );
  XNOR2_X1 U511 ( .A(G218GAT), .B(G106GAT), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n454), .B(n453), .ZN(n481) );
  NOR2_X1 U514 ( .A1(n580), .A2(n481), .ZN(n458) );
  XNOR2_X1 U515 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n547), .A2(n459), .ZN(n577) );
  NAND2_X1 U517 ( .A1(n577), .A2(n390), .ZN(n463) );
  XOR2_X1 U518 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n461) );
  INV_X1 U519 ( .A(G190GAT), .ZN(n460) );
  XOR2_X1 U520 ( .A(KEYINPUT100), .B(KEYINPUT26), .Z(n466) );
  NAND2_X1 U521 ( .A1(n481), .A2(n464), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U523 ( .A(KEYINPUT99), .B(n467), .ZN(n579) );
  XNOR2_X1 U524 ( .A(KEYINPUT27), .B(KEYINPUT97), .ZN(n468) );
  XOR2_X1 U525 ( .A(n468), .B(n537), .Z(n479) );
  OR2_X1 U526 ( .A1(n579), .A2(n479), .ZN(n475) );
  NOR2_X1 U527 ( .A1(n547), .A2(n469), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n481), .A2(n470), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n475), .A2(n474), .ZN(n477) );
  NAND2_X1 U530 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U531 ( .A(n478), .B(KEYINPUT102), .ZN(n485) );
  NOR2_X1 U532 ( .A1(n479), .A2(n535), .ZN(n480) );
  XOR2_X1 U533 ( .A(KEYINPUT98), .B(n480), .Z(n543) );
  XOR2_X1 U534 ( .A(n481), .B(KEYINPUT28), .Z(n545) );
  INV_X1 U535 ( .A(n545), .ZN(n482) );
  NOR2_X1 U536 ( .A1(n543), .A2(n482), .ZN(n483) );
  NAND2_X1 U537 ( .A1(n483), .A2(n547), .ZN(n484) );
  NAND2_X1 U538 ( .A1(n485), .A2(n484), .ZN(n502) );
  NAND2_X1 U539 ( .A1(n498), .A2(n502), .ZN(n486) );
  XOR2_X1 U540 ( .A(KEYINPUT106), .B(n486), .Z(n488) );
  NAND2_X1 U541 ( .A1(n488), .A2(n487), .ZN(n489) );
  XOR2_X1 U542 ( .A(KEYINPUT37), .B(n489), .Z(n534) );
  NAND2_X1 U543 ( .A1(n571), .A2(n490), .ZN(n504) );
  NOR2_X1 U544 ( .A1(n534), .A2(n504), .ZN(n491) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(n491), .Z(n518) );
  NOR2_X1 U546 ( .A1(n518), .A2(n537), .ZN(n494) );
  INV_X1 U547 ( .A(G36GAT), .ZN(n492) );
  XNOR2_X1 U548 ( .A(n492), .B(KEYINPUT108), .ZN(n493) );
  XNOR2_X1 U549 ( .A(n494), .B(n493), .ZN(G1329GAT) );
  NOR2_X1 U550 ( .A1(n518), .A2(n547), .ZN(n497) );
  NOR2_X1 U551 ( .A1(n390), .A2(n498), .ZN(n500) );
  XNOR2_X1 U552 ( .A(KEYINPUT16), .B(KEYINPUT79), .ZN(n499) );
  XNOR2_X1 U553 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U554 ( .A(KEYINPUT78), .B(n501), .Z(n503) );
  NAND2_X1 U555 ( .A1(n503), .A2(n502), .ZN(n524) );
  OR2_X1 U556 ( .A1(n504), .A2(n524), .ZN(n512) );
  NOR2_X1 U557 ( .A1(n535), .A2(n512), .ZN(n505) );
  XOR2_X1 U558 ( .A(G1GAT), .B(n505), .Z(n506) );
  XNOR2_X1 U559 ( .A(KEYINPUT34), .B(n506), .ZN(G1324GAT) );
  NOR2_X1 U560 ( .A1(n537), .A2(n512), .ZN(n507) );
  XOR2_X1 U561 ( .A(G8GAT), .B(n507), .Z(G1325GAT) );
  NOR2_X1 U562 ( .A1(n512), .A2(n547), .ZN(n511) );
  XOR2_X1 U563 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n509) );
  XNOR2_X1 U564 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n508) );
  XNOR2_X1 U565 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U566 ( .A(n511), .B(n510), .ZN(G1326GAT) );
  NOR2_X1 U567 ( .A1(n545), .A2(n512), .ZN(n513) );
  XOR2_X1 U568 ( .A(G22GAT), .B(n513), .Z(G1327GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n515) );
  XNOR2_X1 U570 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n514) );
  XNOR2_X1 U571 ( .A(n515), .B(n514), .ZN(n517) );
  NOR2_X1 U572 ( .A1(n518), .A2(n535), .ZN(n516) );
  XOR2_X1 U573 ( .A(n517), .B(n516), .Z(G1328GAT) );
  NOR2_X1 U574 ( .A1(n545), .A2(n518), .ZN(n519) );
  XOR2_X1 U575 ( .A(G50GAT), .B(n519), .Z(G1331GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n521) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U578 ( .A(n521), .B(n520), .ZN(n526) );
  INV_X1 U579 ( .A(n385), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n523), .A2(n522), .ZN(n533) );
  OR2_X1 U581 ( .A1(n533), .A2(n524), .ZN(n529) );
  NOR2_X1 U582 ( .A1(n535), .A2(n529), .ZN(n525) );
  XOR2_X1 U583 ( .A(n526), .B(n525), .Z(G1332GAT) );
  NOR2_X1 U584 ( .A1(n537), .A2(n529), .ZN(n527) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n527), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n547), .A2(n529), .ZN(n528) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n528), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n545), .A2(n529), .ZN(n531) );
  XNOR2_X1 U589 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n530) );
  XNOR2_X1 U590 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U591 ( .A(G78GAT), .B(n532), .Z(G1335GAT) );
  OR2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U593 ( .A1(n535), .A2(n540), .ZN(n536) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n536), .Z(G1336GAT) );
  NOR2_X1 U595 ( .A1(n537), .A2(n540), .ZN(n538) );
  XOR2_X1 U596 ( .A(G92GAT), .B(n538), .Z(G1337GAT) );
  NOR2_X1 U597 ( .A1(n547), .A2(n540), .ZN(n539) );
  XOR2_X1 U598 ( .A(G99GAT), .B(n539), .Z(G1338GAT) );
  NOR2_X1 U599 ( .A1(n545), .A2(n540), .ZN(n541) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(n541), .Z(n542) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n542), .ZN(G1339GAT) );
  NOR2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n559) );
  NAND2_X1 U603 ( .A1(n545), .A2(n559), .ZN(n546) );
  NOR2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n553) );
  NAND2_X1 U605 ( .A1(n571), .A2(n553), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .Z(n550) );
  NAND2_X1 U608 ( .A1(n553), .A2(n522), .ZN(n549) );
  XNOR2_X1 U609 ( .A(n550), .B(n549), .ZN(G1341GAT) );
  NAND2_X1 U610 ( .A1(n553), .A2(n589), .ZN(n551) );
  XNOR2_X1 U611 ( .A(n551), .B(KEYINPUT50), .ZN(n552) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U614 ( .A1(n553), .A2(n390), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT116), .Z(n556) );
  XNOR2_X1 U617 ( .A(n557), .B(n556), .ZN(G1343GAT) );
  INV_X1 U618 ( .A(n579), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n560), .B(KEYINPUT117), .ZN(n569) );
  NAND2_X1 U621 ( .A1(n569), .A2(n385), .ZN(n561) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(n561), .ZN(G1344GAT) );
  NAND2_X1 U623 ( .A1(n569), .A2(n522), .ZN(n567) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n563) );
  XNOR2_X1 U625 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT52), .Z(n564) );
  XNOR2_X1 U628 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U629 ( .A(n567), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n569), .A2(n589), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n390), .A2(n569), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U634 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n577), .A2(n522), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT56), .Z(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n589), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT125), .Z(n582) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n591) );
  NAND2_X1 U645 ( .A1(n591), .A2(n385), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n587) );
  NAND2_X1 U650 ( .A1(n591), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n588), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n591), .A2(n589), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U655 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n593) );
  NAND2_X1 U656 ( .A1(n591), .A2(n487), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

