

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X2 U325 ( .A(n359), .B(n358), .ZN(n582) );
  XNOR2_X1 U326 ( .A(n481), .B(n480), .ZN(n568) );
  NOR2_X1 U327 ( .A1(n450), .A2(n449), .ZN(n451) );
  NOR2_X1 U328 ( .A1(n586), .A2(n453), .ZN(n454) );
  XOR2_X1 U329 ( .A(KEYINPUT38), .B(n455), .Z(n505) );
  INV_X1 U330 ( .A(KEYINPUT83), .ZN(n406) );
  XNOR2_X1 U331 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U332 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U333 ( .A(n425), .B(n408), .ZN(n409) );
  INV_X1 U334 ( .A(KEYINPUT64), .ZN(n474) );
  XNOR2_X1 U335 ( .A(n339), .B(n338), .ZN(n341) );
  XNOR2_X1 U336 ( .A(n475), .B(n474), .ZN(n573) );
  XNOR2_X1 U337 ( .A(n420), .B(n419), .ZN(n532) );
  XNOR2_X1 U338 ( .A(G183GAT), .B(KEYINPUT126), .ZN(n482) );
  XNOR2_X1 U339 ( .A(n456), .B(G43GAT), .ZN(n457) );
  XNOR2_X1 U340 ( .A(n483), .B(n482), .ZN(G1350GAT) );
  XNOR2_X1 U341 ( .A(n458), .B(n457), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT68), .B(KEYINPUT73), .Z(n294) );
  XNOR2_X1 U343 ( .A(KEYINPUT70), .B(KEYINPUT67), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n307) );
  XOR2_X1 U345 ( .A(G15GAT), .B(G197GAT), .Z(n296) );
  XNOR2_X1 U346 ( .A(G50GAT), .B(G36GAT), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U348 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n298) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT30), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U351 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U352 ( .A(G141GAT), .B(G22GAT), .Z(n399) );
  XOR2_X1 U353 ( .A(G169GAT), .B(G8GAT), .Z(n431) );
  XOR2_X1 U354 ( .A(G1GAT), .B(KEYINPUT72), .Z(n348) );
  XOR2_X1 U355 ( .A(n431), .B(n348), .Z(n302) );
  NAND2_X1 U356 ( .A1(G229GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n399), .B(n303), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U361 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n309) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(G29GAT), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U364 ( .A(KEYINPUT8), .B(n310), .ZN(n340) );
  XNOR2_X1 U365 ( .A(n311), .B(n340), .ZN(n574) );
  INV_X1 U366 ( .A(n574), .ZN(n546) );
  XOR2_X1 U367 ( .A(KEYINPUT13), .B(KEYINPUT74), .Z(n313) );
  XNOR2_X1 U368 ( .A(G71GAT), .B(G57GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n351) );
  XOR2_X1 U370 ( .A(G99GAT), .B(G85GAT), .Z(n325) );
  XOR2_X1 U371 ( .A(n351), .B(n325), .Z(n315) );
  NAND2_X1 U372 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U374 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n317) );
  XNOR2_X1 U375 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U377 ( .A(n319), .B(n318), .Z(n324) );
  XNOR2_X1 U378 ( .A(G106GAT), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n320), .B(G148GAT), .ZN(n390) );
  XOR2_X1 U380 ( .A(G64GAT), .B(G92GAT), .Z(n322) );
  XNOR2_X1 U381 ( .A(G176GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n428) );
  XNOR2_X1 U383 ( .A(n390), .B(n428), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n578) );
  NOR2_X1 U385 ( .A1(n546), .A2(n578), .ZN(n488) );
  XOR2_X1 U386 ( .A(KEYINPUT10), .B(n325), .Z(n327) );
  XOR2_X1 U387 ( .A(G50GAT), .B(G162GAT), .Z(n398) );
  XNOR2_X1 U388 ( .A(G218GAT), .B(n398), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n333) );
  XNOR2_X1 U390 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n328), .B(KEYINPUT76), .ZN(n424) );
  INV_X1 U392 ( .A(KEYINPUT75), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n424), .B(n329), .ZN(n331) );
  NAND2_X1 U394 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U396 ( .A(n333), .B(n332), .Z(n339) );
  XOR2_X1 U397 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n335) );
  XNOR2_X1 U398 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n337) );
  XNOR2_X1 U400 ( .A(G134GAT), .B(G106GAT), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n559) );
  XNOR2_X1 U402 ( .A(KEYINPUT36), .B(n559), .ZN(n586) );
  XOR2_X1 U403 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n343) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U405 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U406 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n345) );
  XNOR2_X1 U407 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n359) );
  XOR2_X1 U410 ( .A(G183GAT), .B(KEYINPUT77), .Z(n430) );
  XOR2_X1 U411 ( .A(n430), .B(G78GAT), .Z(n350) );
  XNOR2_X1 U412 ( .A(n348), .B(G155GAT), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n355) );
  XOR2_X1 U414 ( .A(G15GAT), .B(G127GAT), .Z(n414) );
  XOR2_X1 U415 ( .A(n351), .B(n414), .Z(n353) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U418 ( .A(n355), .B(n354), .Z(n357) );
  XNOR2_X1 U419 ( .A(G22GAT), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U421 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n361) );
  XNOR2_X1 U422 ( .A(KEYINPUT5), .B(KEYINPUT94), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U424 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n363) );
  XNOR2_X1 U425 ( .A(G1GAT), .B(KEYINPUT89), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U427 ( .A(n365), .B(n364), .Z(n371) );
  XNOR2_X1 U428 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n366), .B(KEYINPUT2), .ZN(n391) );
  XOR2_X1 U430 ( .A(G85GAT), .B(n391), .Z(n368) );
  NAND2_X1 U431 ( .A1(G225GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U433 ( .A(G29GAT), .B(n369), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U435 ( .A(G162GAT), .B(G148GAT), .Z(n373) );
  XNOR2_X1 U436 ( .A(G141GAT), .B(G127GAT), .ZN(n372) );
  XNOR2_X1 U437 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U438 ( .A(n375), .B(n374), .Z(n383) );
  XOR2_X1 U439 ( .A(KEYINPUT82), .B(G134GAT), .Z(n377) );
  XNOR2_X1 U440 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U442 ( .A(G113GAT), .B(n378), .Z(n410) );
  XOR2_X1 U443 ( .A(G57GAT), .B(KEYINPUT92), .Z(n380) );
  XNOR2_X1 U444 ( .A(KEYINPUT6), .B(KEYINPUT91), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n410), .B(n381), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n383), .B(n382), .ZN(n520) );
  XOR2_X1 U448 ( .A(KEYINPUT21), .B(G218GAT), .Z(n385) );
  XNOR2_X1 U449 ( .A(KEYINPUT87), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U451 ( .A(G197GAT), .B(n386), .Z(n434) );
  XOR2_X1 U452 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n388) );
  NAND2_X1 U453 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U455 ( .A(n389), .B(KEYINPUT22), .Z(n393) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U458 ( .A(G204GAT), .B(KEYINPUT85), .Z(n395) );
  XNOR2_X1 U459 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U461 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n434), .B(n402), .ZN(n476) );
  XOR2_X1 U465 ( .A(KEYINPUT84), .B(KEYINPUT65), .Z(n404) );
  XNOR2_X1 U466 ( .A(G169GAT), .B(G71GAT), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n420) );
  XNOR2_X1 U468 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n405), .B(KEYINPUT17), .ZN(n425) );
  NAND2_X1 U470 ( .A1(G227GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n418) );
  XOR2_X1 U472 ( .A(G176GAT), .B(G183GAT), .Z(n412) );
  XNOR2_X1 U473 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U475 ( .A(n413), .B(G99GAT), .Z(n416) );
  XNOR2_X1 U476 ( .A(G43GAT), .B(n414), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  INV_X1 U479 ( .A(n532), .ZN(n440) );
  XOR2_X1 U480 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n422) );
  NAND2_X1 U481 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U483 ( .A(n423), .B(KEYINPUT97), .Z(n427) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U486 ( .A(n429), .B(n428), .Z(n433) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n522) );
  INV_X1 U490 ( .A(n522), .ZN(n470) );
  NOR2_X1 U491 ( .A1(n440), .A2(n470), .ZN(n436) );
  XNOR2_X1 U492 ( .A(KEYINPUT100), .B(n436), .ZN(n437) );
  NOR2_X1 U493 ( .A1(n476), .A2(n437), .ZN(n439) );
  XNOR2_X1 U494 ( .A(KEYINPUT101), .B(KEYINPUT25), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n445) );
  NAND2_X1 U496 ( .A1(n476), .A2(n440), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n441), .B(KEYINPUT26), .ZN(n572) );
  XOR2_X1 U498 ( .A(n470), .B(KEYINPUT27), .Z(n447) );
  INV_X1 U499 ( .A(n447), .ZN(n442) );
  NOR2_X1 U500 ( .A1(n442), .A2(n572), .ZN(n443) );
  XOR2_X1 U501 ( .A(KEYINPUT99), .B(n443), .Z(n444) );
  NOR2_X1 U502 ( .A1(n445), .A2(n444), .ZN(n446) );
  NOR2_X1 U503 ( .A1(n520), .A2(n446), .ZN(n450) );
  NAND2_X1 U504 ( .A1(n447), .A2(n520), .ZN(n448) );
  XOR2_X1 U505 ( .A(KEYINPUT98), .B(n448), .Z(n544) );
  XOR2_X1 U506 ( .A(KEYINPUT28), .B(n476), .Z(n496) );
  NAND2_X1 U507 ( .A1(n544), .A2(n496), .ZN(n530) );
  NOR2_X1 U508 ( .A1(n530), .A2(n532), .ZN(n449) );
  XNOR2_X1 U509 ( .A(KEYINPUT102), .B(n451), .ZN(n486) );
  NOR2_X1 U510 ( .A1(n582), .A2(n486), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n452), .B(KEYINPUT107), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT37), .B(n454), .Z(n517) );
  NAND2_X1 U513 ( .A1(n488), .A2(n517), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n505), .A2(n532), .ZN(n458) );
  XOR2_X1 U515 ( .A(KEYINPUT40), .B(KEYINPUT109), .Z(n456) );
  INV_X1 U516 ( .A(KEYINPUT124), .ZN(n481) );
  XOR2_X1 U517 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n463) );
  XNOR2_X1 U518 ( .A(KEYINPUT41), .B(n578), .ZN(n549) );
  NOR2_X1 U519 ( .A1(n546), .A2(n549), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n459), .B(KEYINPUT46), .ZN(n460) );
  NOR2_X1 U521 ( .A1(n582), .A2(n460), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n461), .A2(n559), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n463), .B(n462), .ZN(n468) );
  INV_X1 U524 ( .A(n582), .ZN(n555) );
  NOR2_X1 U525 ( .A1(n586), .A2(n555), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n464), .B(KEYINPUT45), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n465), .A2(n546), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n578), .A2(n466), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT48), .ZN(n543) );
  NOR2_X1 U531 ( .A1(n470), .A2(n543), .ZN(n472) );
  INV_X1 U532 ( .A(KEYINPUT54), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U534 ( .A1(n473), .A2(n520), .ZN(n475) );
  NOR2_X1 U535 ( .A1(n573), .A2(n476), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n532), .A2(n479), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n568), .A2(n582), .ZN(n483) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n485) );
  NAND2_X1 U541 ( .A1(n582), .A2(n559), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(n487) );
  NOR2_X1 U543 ( .A1(n487), .A2(n486), .ZN(n509) );
  AND2_X1 U544 ( .A1(n488), .A2(n509), .ZN(n497) );
  NAND2_X1 U545 ( .A1(n497), .A2(n520), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n489), .B(KEYINPUT34), .ZN(n490) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n490), .ZN(G1324GAT) );
  XOR2_X1 U548 ( .A(G8GAT), .B(KEYINPUT103), .Z(n492) );
  NAND2_X1 U549 ( .A1(n497), .A2(n522), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n494) );
  NAND2_X1 U552 ( .A1(n497), .A2(n532), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(n495), .ZN(G1326GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n499) );
  INV_X1 U556 ( .A(n496), .ZN(n526) );
  NAND2_X1 U557 ( .A1(n497), .A2(n526), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U559 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  XOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .Z(n502) );
  NAND2_X1 U561 ( .A1(n520), .A2(n505), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n505), .A2(n522), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT108), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G36GAT), .B(n504), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n505), .A2(n526), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT110), .B(KEYINPUT112), .Z(n508) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(n511) );
  XNOR2_X1 U571 ( .A(KEYINPUT111), .B(n549), .ZN(n563) );
  AND2_X1 U572 ( .A1(n546), .A2(n563), .ZN(n518) );
  AND2_X1 U573 ( .A1(n518), .A2(n509), .ZN(n514) );
  NAND2_X1 U574 ( .A1(n514), .A2(n520), .ZN(n510) );
  XOR2_X1 U575 ( .A(n511), .B(n510), .Z(G1332GAT) );
  NAND2_X1 U576 ( .A1(n522), .A2(n514), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n532), .A2(n514), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U581 ( .A1(n514), .A2(n526), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(KEYINPUT113), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n527), .A2(n520), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n527), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n532), .A2(n527), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT114), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n543), .A2(n530), .ZN(n531) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U597 ( .A(KEYINPUT116), .B(n533), .Z(n540) );
  NAND2_X1 U598 ( .A1(n540), .A2(n574), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n536) );
  NAND2_X1 U601 ( .A1(n563), .A2(n540), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n582), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  INV_X1 U608 ( .A(n559), .ZN(n569) );
  NAND2_X1 U609 ( .A1(n569), .A2(n540), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n572), .A2(n543), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n558) );
  NOR2_X1 U613 ( .A1(n546), .A2(n558), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT118), .B(n547), .Z(n548) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n558), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(KEYINPUT53), .B(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n558), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT122), .B(n560), .Z(n561) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n568), .A2(n574), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n563), .A2(n568), .ZN(n565) );
  XOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT125), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n584) );
  NAND2_X1 U640 ( .A1(n584), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n584), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U649 ( .A(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

