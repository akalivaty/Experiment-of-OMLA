//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1286, new_n1287, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(KEYINPUT68), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT66), .B(G77), .Z(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT67), .B(G244), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n212), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n211), .A2(KEYINPUT68), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT69), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n208), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n226), .B(new_n232), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n223), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT70), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT16), .ZN(new_n252));
  INV_X1    g0052(.A(G68), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n230), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n257), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n253), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G58), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n253), .ZN(new_n264));
  OAI21_X1  g0064(.A(G20), .B1(new_n264), .B2(new_n201), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G159), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n252), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT80), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n229), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n260), .A2(new_n261), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n268), .B1(new_n275), .B2(G68), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n274), .B1(new_n276), .B2(KEYINPUT16), .ZN(new_n277));
  OAI211_X1 g0077(.A(KEYINPUT80), .B(new_n252), .C1(new_n262), .C2(new_n268), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT72), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n263), .A2(KEYINPUT72), .A3(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G1), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n273), .B1(new_n285), .B2(G20), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(G13), .A3(G20), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  INV_X1    g0092(.A(G226), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G1698), .ZN(new_n294));
  AND2_X1   g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n294), .B1(G223), .B2(G1698), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G87), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n292), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G41), .ZN(new_n300));
  INV_X1    g0100(.A(G45), .ZN(new_n301));
  AOI21_X1  g0101(.A(G1), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(new_n292), .A3(G274), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n285), .B1(G41), .B2(G45), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n292), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n236), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G200), .B2(new_n307), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n279), .A2(new_n290), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT17), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n279), .A2(KEYINPUT17), .A3(new_n310), .A4(new_n290), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT18), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n279), .A2(new_n290), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n297), .A2(new_n298), .ZN(new_n319));
  INV_X1    g0119(.A(new_n292), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n306), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G179), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n299), .A2(new_n306), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n316), .B1(new_n317), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g0128(.A(KEYINPUT18), .B(new_n326), .C1(new_n279), .C2(new_n290), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n315), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n292), .A2(G238), .A3(new_n304), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n303), .A2(new_n333), .A3(KEYINPUT78), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT78), .B1(new_n303), .B2(new_n333), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n293), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n236), .A2(G1698), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n338), .B(new_n339), .C1(new_n295), .C2(new_n296), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(KEYINPUT77), .A3(new_n341), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(new_n320), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n336), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n336), .B2(new_n346), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n332), .B(G169), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT79), .ZN(new_n351));
  INV_X1    g0151(.A(new_n345), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT77), .B1(new_n340), .B2(new_n341), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n352), .A2(new_n353), .A3(new_n292), .ZN(new_n354));
  INV_X1    g0154(.A(new_n335), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n303), .A2(new_n333), .A3(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT13), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n336), .A2(new_n346), .A3(new_n347), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT79), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(new_n332), .A4(G169), .ZN(new_n362));
  OAI21_X1  g0162(.A(G169), .B1(new_n348), .B2(new_n349), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT14), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n358), .A2(G179), .A3(new_n359), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n351), .A2(new_n362), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n286), .A2(G68), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT12), .ZN(new_n368));
  INV_X1    g0168(.A(new_n288), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n253), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n288), .A2(KEYINPUT12), .A3(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n253), .ZN(new_n373));
  INV_X1    g0173(.A(G77), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n230), .A2(G33), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n376), .A2(KEYINPUT11), .A3(new_n273), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT11), .B1(new_n376), .B2(new_n273), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n372), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n366), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n360), .A2(G200), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n358), .A2(G190), .A3(new_n359), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n305), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G226), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n303), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT71), .ZN(new_n389));
  AOI21_X1  g0189(.A(G1698), .B1(new_n256), .B2(new_n257), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G222), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n256), .A2(new_n257), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(G223), .A3(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n391), .B(new_n393), .C1(new_n213), .C2(new_n392), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n320), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT71), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n387), .A2(new_n396), .A3(new_n303), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G200), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n389), .A2(new_n395), .A3(G190), .A4(new_n397), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT10), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT9), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n288), .A2(G50), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n286), .B2(G50), .ZN(new_n406));
  INV_X1    g0206(.A(new_n375), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n282), .A2(new_n407), .A3(new_n283), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n266), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n404), .B(new_n406), .C1(new_n410), .C2(new_n274), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n274), .B1(new_n408), .B2(new_n409), .ZN(new_n412));
  INV_X1    g0212(.A(new_n406), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT9), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n399), .A2(new_n415), .A3(new_n400), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n403), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n401), .A3(new_n402), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n398), .A2(new_n318), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n406), .B1(new_n410), .B2(new_n274), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(G179), .C2(new_n398), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n392), .A2(G238), .A3(G1698), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n392), .A2(G232), .A3(new_n337), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT73), .B(G107), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n424), .B(new_n425), .C1(new_n392), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n320), .ZN(new_n428));
  INV_X1    g0228(.A(G274), .ZN(new_n429));
  AND2_X1   g0229(.A1(G1), .A2(G13), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(new_n291), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n386), .A2(new_n215), .B1(new_n302), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n428), .A2(new_n324), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(G169), .B1(new_n428), .B2(new_n432), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n213), .A2(new_n230), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n263), .A2(KEYINPUT8), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT8), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G58), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT74), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT74), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n280), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n436), .B1(new_n444), .B2(new_n266), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT15), .B(G87), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n445), .A2(KEYINPUT75), .B1(new_n407), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n440), .A2(KEYINPUT74), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n280), .A2(new_n442), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n266), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n436), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT75), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n274), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n286), .A2(G77), .B1(new_n213), .B2(new_n369), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n435), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n451), .A2(KEYINPUT75), .A3(new_n452), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n447), .A2(new_n407), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n445), .A2(KEYINPUT75), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n273), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n428), .A2(new_n432), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G200), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n428), .A2(G190), .A3(new_n432), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n457), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  NOR4_X1   g0269(.A1(new_n331), .A2(new_n385), .A3(new_n423), .A4(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n285), .A2(G33), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n288), .A2(new_n472), .A3(new_n229), .A4(new_n272), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G116), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(G116), .B2(new_n369), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  AOI221_X4 g0276(.A(KEYINPUT86), .B1(new_n476), .B2(G20), .C1(new_n272), .C2(new_n229), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT86), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(G20), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n273), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n482), .B(new_n230), .C1(G33), .C2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n255), .A2(G97), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(KEYINPUT87), .A3(new_n230), .A4(new_n482), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n481), .A2(KEYINPUT20), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT20), .B1(new_n481), .B2(new_n489), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n475), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n301), .A2(G1), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G270), .A3(new_n292), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT84), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n500), .A3(G270), .A4(new_n292), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G264), .B(G1698), .C1(new_n295), .C2(new_n296), .ZN(new_n503));
  OAI211_X1 g0303(.A(G257), .B(new_n337), .C1(new_n295), .C2(new_n296), .ZN(new_n504));
  INV_X1    g0304(.A(G303), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n503), .B(new_n504), .C1(new_n505), .C2(new_n392), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n320), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n292), .A2(G274), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n497), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n502), .A2(G179), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n493), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n502), .A2(new_n507), .A3(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n499), .B2(new_n501), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT85), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n507), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n514), .A2(new_n492), .A3(G169), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT88), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n512), .B1(new_n519), .B2(KEYINPUT21), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT88), .ZN(new_n521));
  AND4_X1   g0321(.A1(new_n516), .A2(new_n502), .A3(new_n507), .A4(new_n510), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n516), .B1(new_n515), .B2(new_n507), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n480), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n273), .A2(new_n478), .A3(new_n479), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n489), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n481), .A2(KEYINPUT20), .A3(new_n489), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n318), .B1(new_n531), .B2(new_n475), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n521), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n514), .A2(G200), .A3(new_n517), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n536), .B(new_n493), .C1(new_n524), .C2(new_n308), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n520), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(G257), .B(G1698), .C1(new_n295), .C2(new_n296), .ZN(new_n539));
  OAI211_X1 g0339(.A(G250), .B(new_n337), .C1(new_n295), .C2(new_n296), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G294), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n320), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n497), .A2(G264), .A3(new_n292), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n510), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G169), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT89), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n497), .A2(new_n548), .A3(G264), .A4(new_n292), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n509), .B1(new_n320), .B2(new_n542), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n546), .B1(new_n324), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n230), .B(G87), .C1(new_n295), .C2(new_n296), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT22), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n392), .A2(new_n557), .A3(new_n230), .A4(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(G107), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G20), .ZN(new_n561));
  OAI22_X1  g0361(.A1(KEYINPUT23), .A2(new_n561), .B1(new_n375), .B2(new_n476), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n426), .A2(G20), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(KEYINPUT23), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n554), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(new_n564), .A3(new_n554), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n274), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(G13), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n561), .A2(G1), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n570), .B(KEYINPUT25), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT81), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n274), .A2(new_n572), .A3(new_n288), .A4(new_n472), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n473), .A2(KEYINPUT81), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n574), .A3(G107), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n553), .B1(new_n568), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n567), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n273), .B1(new_n578), .B2(new_n565), .ZN(new_n579));
  INV_X1    g0379(.A(new_n576), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n545), .A2(G190), .ZN(new_n581));
  AOI21_X1  g0381(.A(G200), .B1(new_n550), .B2(new_n551), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n573), .A2(new_n574), .A3(G97), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n369), .A2(new_n483), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n266), .A2(G77), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT6), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n589), .A2(new_n483), .A3(G107), .ZN(new_n590));
  XNOR2_X1  g0390(.A(G97), .B(G107), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n588), .B1(new_n592), .B2(new_n230), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n426), .B1(new_n260), .B2(new_n261), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n273), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G250), .B(G1698), .C1(new_n295), .C2(new_n296), .ZN(new_n597));
  OAI211_X1 g0397(.A(G244), .B(new_n337), .C1(new_n295), .C2(new_n296), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n482), .B(new_n597), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT4), .B1(new_n390), .B2(G244), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n320), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n497), .A2(G257), .A3(new_n292), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n510), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n596), .B1(G200), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n603), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n598), .A2(new_n599), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n392), .A2(KEYINPUT4), .A3(G244), .A4(new_n337), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n482), .A4(new_n597), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n606), .B1(new_n609), .B2(new_n320), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(G190), .A3(new_n510), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n324), .A3(new_n510), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n318), .A2(new_n604), .B1(new_n587), .B2(new_n595), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n605), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  OR2_X1    g0415(.A1(G238), .A2(G1698), .ZN(new_n616));
  INV_X1    g0416(.A(G244), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G1698), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n616), .B(new_n618), .C1(new_n295), .C2(new_n296), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G116), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n292), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G250), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n285), .B2(G45), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n292), .ZN(new_n624));
  INV_X1    g0424(.A(new_n494), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n624), .B1(new_n508), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n615), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n431), .A2(new_n494), .B1(new_n292), .B2(new_n623), .ZN(new_n629));
  INV_X1    g0429(.A(new_n620), .ZN(new_n630));
  NOR2_X1   g0430(.A1(G238), .A2(G1698), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n617), .B2(G1698), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n630), .B1(new_n632), .B2(new_n392), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n629), .B(KEYINPUT82), .C1(new_n633), .C2(new_n292), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n318), .B1(new_n628), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n627), .A2(new_n634), .A3(new_n324), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT83), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT83), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n627), .A2(new_n634), .A3(new_n639), .A4(new_n324), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n392), .A2(new_n230), .A3(G68), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n375), .A2(new_n483), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(KEYINPUT19), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(G87), .A2(G97), .ZN(new_n644));
  NAND3_X1  g0444(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n426), .A2(new_n644), .B1(new_n230), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n273), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n446), .A2(new_n369), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n573), .A2(new_n574), .A3(new_n447), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n636), .A2(new_n638), .A3(new_n640), .A4(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(G200), .B1(new_n628), .B2(new_n635), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n573), .A2(new_n574), .A3(G87), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n627), .A2(new_n634), .A3(G190), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n584), .A2(new_n614), .A3(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n471), .A2(new_n538), .A3(new_n658), .ZN(G372));
  NOR2_X1   g0459(.A1(new_n328), .A2(new_n329), .ZN(new_n660));
  INV_X1    g0460(.A(new_n459), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n366), .B2(new_n380), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n313), .A2(new_n314), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n384), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n418), .A3(new_n419), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n422), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n604), .A2(new_n318), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n669), .A2(new_n612), .A3(new_n596), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n651), .A3(new_n656), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT26), .ZN(new_n672));
  INV_X1    g0472(.A(new_n621), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n629), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT90), .B1(new_n674), .B2(new_n318), .ZN(new_n675));
  OAI211_X1 g0475(.A(KEYINPUT90), .B(new_n318), .C1(new_n621), .C2(new_n626), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n650), .B(new_n637), .C1(new_n675), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(G200), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n654), .A2(new_n655), .A3(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(new_n670), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n672), .A2(new_n683), .A3(new_n678), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT91), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n577), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n553), .B(KEYINPUT91), .C1(new_n568), .C2(new_n576), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n520), .A2(new_n688), .A3(new_n535), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n614), .A2(new_n583), .A3(new_n681), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n684), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n668), .B1(new_n471), .B2(new_n691), .ZN(G369));
  INV_X1    g0492(.A(G330), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n285), .A2(new_n230), .A3(G13), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT92), .ZN(new_n696));
  OAI21_X1  g0496(.A(G213), .B1(new_n694), .B2(KEYINPUT27), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n492), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n512), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n533), .B2(new_n534), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n518), .A2(KEYINPUT88), .A3(new_n534), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n520), .A2(new_n535), .A3(new_n537), .A4(new_n702), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n693), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n584), .ZN(new_n710));
  INV_X1    g0510(.A(new_n701), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n579), .B2(new_n580), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n710), .A2(new_n712), .B1(new_n577), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n686), .A2(new_n687), .A3(new_n711), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n701), .B1(new_n520), .B2(new_n535), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n584), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n714), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n224), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n228), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n426), .A2(new_n476), .A3(new_n644), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G1), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n722), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n627), .A2(new_n550), .A3(new_n551), .A4(new_n634), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n602), .A2(new_n603), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n729), .A2(new_n511), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n728), .B1(new_n731), .B2(KEYINPUT93), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT93), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n550), .A2(new_n551), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(new_n610), .A3(new_n627), .A4(new_n634), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n733), .B(KEYINPUT30), .C1(new_n735), .C2(new_n511), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n324), .B1(new_n621), .B2(new_n626), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n551), .B2(new_n550), .ZN(new_n739));
  AND4_X1   g0539(.A1(new_n514), .A2(new_n517), .A3(new_n604), .A4(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n711), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n742), .A2(KEYINPUT94), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT94), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n740), .B1(new_n732), .B2(new_n736), .ZN(new_n747));
  INV_X1    g0547(.A(new_n744), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n743), .B1(new_n747), .B2(new_n711), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n745), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n538), .A2(new_n658), .A3(new_n701), .ZN(new_n752));
  OAI21_X1  g0552(.A(G330), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n678), .A2(new_n680), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n613), .A2(new_n612), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT26), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n670), .A2(new_n651), .A3(new_n682), .A4(new_n656), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(new_n678), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n520), .A2(new_n535), .A3(new_n577), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(new_n690), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT29), .B1(new_n760), .B2(new_n701), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT29), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n614), .A2(new_n583), .A3(new_n681), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n534), .B1(new_n518), .B2(KEYINPUT88), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n706), .A2(new_n764), .A3(new_n512), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n763), .B1(new_n765), .B2(new_n688), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n762), .B(new_n711), .C1(new_n766), .C2(new_n684), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n753), .A2(new_n761), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n727), .B1(new_n769), .B2(G1), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT95), .Z(G364));
  INV_X1    g0571(.A(new_n721), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n569), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n285), .B1(new_n773), .B2(G45), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n772), .A2(KEYINPUT96), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT96), .ZN(new_n776));
  INV_X1    g0576(.A(new_n774), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n721), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n224), .A2(new_n392), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(G116), .B2(new_n224), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n392), .B(new_n720), .C1(new_n301), .C2(new_n228), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n784), .A2(KEYINPUT97), .B1(G45), .B2(new_n250), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n229), .B1(G20), .B2(new_n318), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n780), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n230), .A2(G179), .ZN(new_n795));
  INV_X1    g0595(.A(G200), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n795), .A2(new_n308), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n392), .B1(new_n798), .B2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n230), .A2(new_n796), .A3(G179), .A4(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n799), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n230), .A2(new_n324), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n805), .A2(new_n796), .A3(G190), .ZN(new_n806));
  INV_X1    g0606(.A(G317), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT33), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n807), .A2(KEYINPUT33), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n324), .A2(new_n796), .A3(G190), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n803), .B(new_n815), .C1(G326), .C2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n795), .A2(G190), .A3(G200), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT101), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G303), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n796), .B1(new_n804), .B2(KEYINPUT98), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(KEYINPUT98), .B2(new_n804), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n308), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n826), .A2(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(KEYINPUT100), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G322), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n825), .A2(G190), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT99), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT99), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n822), .B1(new_n823), .B2(new_n830), .C1(new_n831), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n798), .A2(G159), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT32), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n802), .A2(new_n560), .B1(new_n202), .B2(new_n816), .ZN(new_n839));
  INV_X1    g0639(.A(new_n806), .ZN(new_n840));
  INV_X1    g0640(.A(G87), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n840), .A2(new_n253), .B1(new_n819), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n392), .B1(new_n813), .B2(new_n483), .ZN(new_n843));
  NOR4_X1   g0643(.A1(new_n838), .A2(new_n839), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n835), .B2(new_n263), .C1(new_n213), .C2(new_n830), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n836), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n794), .B1(new_n846), .B2(new_n791), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n707), .A2(new_n708), .ZN(new_n848));
  INV_X1    g0648(.A(new_n790), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(G330), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n779), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n848), .A2(G330), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(G396));
  OAI21_X1  g0654(.A(new_n701), .B1(new_n456), .B2(new_n458), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n459), .A2(new_n855), .A3(new_n468), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT103), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n661), .A2(new_n701), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n459), .A2(new_n855), .A3(new_n468), .A4(KEYINPUT103), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n691), .B2(new_n701), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n863));
  INV_X1    g0663(.A(new_n753), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n858), .A2(new_n860), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n711), .B(new_n865), .C1(new_n766), .C2(new_n684), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT104), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n867), .B(new_n861), .C1(new_n691), .C2(new_n701), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n863), .A2(new_n864), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n779), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT105), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n869), .A2(new_n872), .A3(new_n779), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n863), .A2(new_n866), .A3(new_n868), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n871), .B(new_n873), .C1(new_n864), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n791), .A2(new_n788), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n780), .B1(G77), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n392), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n879), .B1(new_n797), .B2(new_n823), .C1(new_n813), .C2(new_n483), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n801), .A2(G87), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n881), .B1(new_n505), .B2(new_n816), .C1(new_n840), .C2(new_n800), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n880), .B(new_n882), .C1(G107), .C2(new_n820), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n883), .B1(new_n814), .B2(new_n835), .C1(new_n476), .C2(new_n830), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n879), .B1(new_n798), .B2(G132), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n885), .B1(new_n263), .B2(new_n813), .C1(new_n253), .C2(new_n802), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(G50), .B2(new_n820), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n806), .A2(G150), .B1(new_n817), .B2(G137), .ZN(new_n888));
  INV_X1    g0688(.A(G143), .ZN(new_n889));
  INV_X1    g0689(.A(G159), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n888), .B1(new_n835), .B2(new_n889), .C1(new_n830), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT34), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n887), .B1(new_n893), .B2(KEYINPUT102), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n884), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n878), .B1(new_n897), .B2(new_n791), .ZN(new_n898));
  INV_X1    g0698(.A(new_n861), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n898), .B1(new_n789), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n875), .A2(new_n900), .ZN(G384));
  INV_X1    g0701(.A(new_n592), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(KEYINPUT35), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(KEYINPUT35), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n903), .A2(G116), .A3(new_n231), .A4(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT36), .Z(new_n906));
  OR3_X1    g0706(.A1(new_n213), .A2(new_n227), .A3(new_n264), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n202), .A2(G68), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n285), .B(G13), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n277), .A2(new_n269), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n698), .B1(new_n913), .B2(new_n289), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n663), .B2(new_n660), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n913), .A2(new_n289), .B1(new_n327), .B2(new_n698), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n917), .B2(new_n311), .ZN(new_n918));
  INV_X1    g0718(.A(new_n311), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n326), .B1(new_n279), .B2(new_n290), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n699), .B1(new_n279), .B2(new_n290), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n918), .B1(new_n922), .B2(new_n916), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n912), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n317), .A2(new_n327), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n317), .A2(new_n698), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n925), .A2(new_n926), .A3(new_n916), .A4(new_n311), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n917), .A2(new_n311), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n916), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(KEYINPUT38), .C1(new_n330), .C2(new_n914), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n924), .A2(KEYINPUT106), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(new_n912), .C1(new_n915), .C2(new_n923), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n711), .A2(new_n379), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n381), .A2(new_n384), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n384), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n380), .B(new_n701), .C1(new_n366), .C2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n861), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n614), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n577), .A2(new_n583), .A3(new_n651), .A4(new_n656), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n943), .A2(new_n765), .A3(new_n537), .A4(new_n711), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n742), .A2(new_n744), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(new_n945), .A3(new_n750), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n911), .B1(new_n934), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n940), .A2(new_n946), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n925), .A2(new_n926), .A3(new_n311), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT37), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n951), .A2(new_n927), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n926), .B1(new_n663), .B2(new_n660), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n912), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n911), .B1(new_n954), .B2(new_n930), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT108), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n470), .A2(new_n946), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n693), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n691), .A2(KEYINPUT29), .A3(new_n701), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n759), .A2(new_n690), .ZN(new_n964));
  INV_X1    g0764(.A(new_n758), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n762), .B1(new_n966), .B2(new_n711), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n470), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n668), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT107), .Z(new_n970));
  NAND3_X1  g0770(.A1(new_n931), .A2(KEYINPUT39), .A3(new_n933), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT39), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n954), .A2(new_n972), .A3(new_n930), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n381), .A2(new_n701), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n660), .A2(new_n698), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n931), .A2(new_n933), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n937), .A2(new_n939), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n459), .A2(new_n701), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n979), .B1(new_n866), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n977), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n976), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n970), .B(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n962), .A2(new_n985), .B1(new_n285), .B2(new_n773), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT109), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n962), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(KEYINPUT109), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n910), .B1(new_n989), .B2(new_n990), .ZN(G367));
  NAND2_X1  g0791(.A1(new_n701), .A2(new_n596), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n614), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(new_n577), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n701), .B1(new_n994), .B2(new_n755), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n670), .A2(new_n701), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n717), .A2(new_n584), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n995), .B1(KEYINPUT42), .B2(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(KEYINPUT42), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n711), .A2(new_n654), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(new_n678), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n681), .A2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n999), .A2(new_n1000), .B1(KEYINPUT43), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(KEYINPUT43), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1005), .B(new_n1006), .Z(new_n1007));
  INV_X1    g0807(.A(new_n997), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n714), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1007), .B(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n721), .B(KEYINPUT41), .Z(new_n1011));
  INV_X1    g0811(.A(KEYINPUT111), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n584), .B(new_n711), .C1(new_n705), .C2(new_n706), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n713), .B2(new_n717), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n851), .B(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1012), .B1(new_n1015), .B2(new_n768), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n963), .A2(new_n967), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1014), .B(new_n709), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1017), .A2(new_n1018), .A3(KEYINPUT111), .A4(new_n753), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n709), .A2(KEYINPUT110), .A3(new_n713), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT44), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n718), .B2(new_n997), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1013), .A2(new_n715), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(KEYINPUT44), .A3(new_n1008), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT45), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1023), .B2(new_n1008), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n718), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1020), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n1025), .A2(new_n1029), .A3(new_n1020), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1016), .B(new_n1019), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1011), .B1(new_n1032), .B2(new_n769), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n774), .B1(new_n1033), .B2(KEYINPUT112), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT112), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1035), .B(new_n1011), .C1(new_n1032), .C2(new_n769), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1010), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT113), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT113), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1010), .B(new_n1039), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n830), .A2(new_n800), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n879), .B1(new_n807), .B2(new_n797), .C1(new_n802), .C2(new_n483), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n813), .A2(new_n426), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n840), .A2(new_n814), .B1(new_n816), .B2(new_n823), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT46), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n820), .B2(G116), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n819), .A2(KEYINPUT46), .A3(new_n476), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1046), .B1(new_n505), .B2(new_n835), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n879), .B1(new_n214), .B2(new_n801), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT115), .ZN(new_n1052));
  INV_X1    g0852(.A(G137), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n813), .A2(new_n253), .B1(new_n1053), .B2(new_n797), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n819), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n806), .A2(G159), .B1(G58), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n889), .B2(new_n816), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1052), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(G150), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n835), .B2(new_n1059), .C1(new_n202), .C2(new_n830), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1050), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT47), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1050), .A2(KEYINPUT47), .A3(new_n1060), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n791), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1002), .A2(new_n790), .A3(new_n1003), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n720), .A2(new_n392), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n243), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n792), .C1(new_n224), .C2(new_n446), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n780), .A2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT114), .Z(new_n1071));
  NAND3_X1  g0871(.A1(new_n1065), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1041), .A2(new_n1072), .ZN(G387));
  NAND2_X1  g0873(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1074), .B(new_n721), .C1(new_n769), .C2(new_n1018), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n392), .B1(new_n1059), .B2(new_n797), .C1(new_n802), .C2(new_n483), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n813), .A2(new_n446), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n213), .A2(new_n819), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n890), .B2(new_n816), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n284), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1076), .B(new_n1080), .C1(new_n1081), .C2(new_n806), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n202), .B2(new_n835), .C1(new_n253), .C2(new_n830), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n392), .B1(new_n798), .B2(G326), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n806), .A2(G311), .B1(new_n817), .B2(G322), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n835), .B2(new_n807), .C1(new_n830), .C2(new_n505), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1055), .A2(G294), .B1(new_n812), .B2(G283), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT49), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1084), .B1(new_n476), .B2(new_n802), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1091), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(KEYINPUT49), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1083), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1096), .A2(new_n791), .ZN(new_n1097));
  AOI21_X1  g0897(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n444), .A2(new_n202), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1100));
  OAI211_X1 g0900(.A(new_n724), .B(new_n1098), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1067), .B1(new_n1101), .B2(new_n1102), .C1(new_n301), .C2(new_n239), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(G107), .B2(new_n224), .C1(new_n724), .C2(new_n781), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n779), .B1(new_n1104), .B2(new_n792), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n713), .B2(new_n849), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1075), .B1(new_n774), .B2(new_n1015), .C1(new_n1097), .C2(new_n1106), .ZN(G393));
  AND2_X1   g0907(.A1(new_n1032), .A2(new_n721), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(new_n714), .Z(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1074), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n792), .B1(new_n224), .B2(new_n483), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1067), .B2(new_n247), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n835), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1115), .A2(G159), .B1(G150), .B2(new_n817), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n1117));
  OR2_X1    g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n806), .A2(G50), .B1(G77), .B2(new_n812), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n879), .B1(new_n798), .B2(G143), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1055), .A2(G68), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1120), .A2(new_n881), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n829), .B2(new_n444), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1118), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n835), .A2(new_n823), .B1(new_n807), .B2(new_n816), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT52), .Z(new_n1127));
  OAI22_X1  g0927(.A1(new_n840), .A2(new_n505), .B1(new_n476), .B2(new_n813), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n879), .B1(new_n831), .B2(new_n797), .C1(new_n802), .C2(new_n560), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(G283), .C2(new_n1055), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n830), .B2(new_n814), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n779), .B(new_n1114), .C1(new_n1132), .C2(new_n791), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1008), .A2(new_n790), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT117), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1110), .B2(new_n774), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1112), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(G390));
  NAND3_X1  g0939(.A1(new_n946), .A2(G330), .A3(new_n899), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n979), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n760), .A2(new_n701), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n980), .B1(new_n1142), .B2(new_n865), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n940), .B(G330), .C1(new_n752), .C2(new_n751), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n946), .A2(G330), .ZN(new_n1146));
  OAI211_X1 g0946(.A(G330), .B(new_n899), .C1(new_n751), .C2(new_n752), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1146), .A2(new_n940), .B1(new_n1147), .B2(new_n979), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n866), .A2(new_n981), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1145), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n470), .A2(G330), .A3(new_n946), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n968), .A2(new_n668), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n971), .B(new_n973), .C1(new_n975), .C2(new_n982), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n975), .B1(new_n954), .B2(new_n930), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1143), .B2(new_n979), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1156), .A2(new_n1158), .A3(new_n1144), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n940), .A2(new_n946), .A3(G330), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1155), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n979), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n975), .B1(new_n1149), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1158), .B1(new_n974), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1160), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1147), .A2(new_n979), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1160), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1149), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1153), .B1(new_n1170), .B2(new_n1145), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1156), .A2(new_n1158), .A3(new_n1144), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1162), .A2(new_n1173), .A3(new_n721), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n974), .A2(new_n789), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n879), .B1(new_n814), .B2(new_n797), .C1(new_n802), .C2(new_n253), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n817), .A2(G283), .B1(G77), .B2(new_n812), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n426), .B2(new_n840), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(G87), .C2(new_n820), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n835), .B2(new_n476), .C1(new_n483), .C2(new_n830), .ZN(new_n1180));
  INV_X1    g0980(.A(G132), .ZN(new_n1181));
  INV_X1    g0981(.A(G128), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n835), .A2(new_n1181), .B1(new_n1182), .B2(new_n816), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT120), .Z(new_n1184));
  OAI21_X1  g0984(.A(new_n392), .B1(new_n802), .B2(new_n202), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT119), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n819), .A2(new_n1059), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT53), .Z(new_n1188));
  AOI22_X1  g0988(.A1(new_n798), .A2(G125), .B1(G159), .B2(new_n812), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n840), .B2(new_n1053), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1186), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n830), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1180), .B1(new_n1184), .B2(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1194), .A2(new_n791), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n780), .B1(new_n1081), .B2(new_n877), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1175), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n777), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1174), .A2(new_n1199), .ZN(G378));
  AOI21_X1  g1000(.A(new_n693), .B1(new_n949), .B2(new_n955), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n421), .A2(new_n698), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT55), .Z(new_n1203));
  XNOR2_X1  g1003(.A(new_n423), .B(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1205));
  XNOR2_X1  g1005(.A(new_n1204), .B(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n948), .A2(new_n1201), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n948), .B2(new_n1201), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1208), .A2(new_n984), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1149), .A2(new_n1163), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1211), .A2(new_n934), .B1(new_n660), .B2(new_n698), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n975), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n971), .B2(new_n973), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n948), .A2(new_n1201), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1206), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n948), .A2(new_n1201), .A3(new_n1207), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n777), .B1(new_n1210), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1192), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n817), .A2(G125), .B1(new_n1055), .B2(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n1059), .B2(new_n813), .C1(new_n1181), .C2(new_n840), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n835), .A2(new_n1182), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G137), .C2(new_n829), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT59), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT121), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1229), .A2(G124), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(G124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n798), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(G33), .A2(G41), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(new_n890), .C2(new_n802), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1227), .A2(new_n1228), .A3(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G50), .B(new_n1233), .C1(new_n879), .C2(new_n300), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G41), .B(new_n392), .C1(new_n798), .C2(G283), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n253), .B2(new_n813), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n840), .A2(new_n483), .B1(new_n263), .B2(new_n802), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n816), .A2(new_n476), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1078), .A4(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n835), .B2(new_n560), .C1(new_n446), .C2(new_n830), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT58), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1236), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1243), .B2(new_n1242), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n791), .B1(new_n1235), .B2(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT122), .Z(new_n1247));
  OAI21_X1  g1047(.A(new_n780), .B1(G50), .B2(new_n877), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1206), .A2(new_n788), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1220), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1173), .A2(new_n1154), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n984), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1217), .A2(new_n1215), .A3(new_n1218), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT57), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n772), .B1(new_n1260), .B2(new_n1253), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1252), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(G375));
  AND2_X1   g1063(.A1(new_n1144), .A2(new_n1143), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1264), .A2(new_n1141), .B1(new_n1169), .B2(new_n1149), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1153), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1011), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1155), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n979), .A2(new_n788), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n780), .B1(G68), .B2(new_n877), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n392), .B1(new_n801), .B2(G77), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT124), .Z(new_n1272));
  AOI21_X1  g1072(.A(new_n1077), .B1(G303), .B2(new_n798), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1273), .B1(new_n476), .B2(new_n840), .C1(new_n814), .C2(new_n816), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1272), .B(new_n1274), .C1(G97), .C2(new_n820), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n800), .B2(new_n835), .C1(new_n426), .C2(new_n830), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n392), .B1(new_n1182), .B2(new_n797), .C1(new_n802), .C2(new_n263), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n806), .A2(new_n1221), .B1(G50), .B2(new_n812), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1181), .B2(new_n816), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1277), .B(new_n1279), .C1(G159), .C2(new_n820), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1280), .B1(new_n835), .B2(new_n1053), .C1(new_n1059), .C2(new_n830), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1276), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1270), .B1(new_n1282), .B2(new_n791), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1151), .A2(new_n777), .B1(new_n1269), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1268), .A2(new_n1284), .ZN(G381));
  NOR3_X1   g1085(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(new_n1138), .A3(new_n1284), .A4(new_n1268), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G387), .A2(new_n1287), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1088(.A(G378), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1262), .A2(new_n700), .A3(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G407), .A2(G213), .A3(new_n1290), .ZN(G409));
  INV_X1    g1091(.A(KEYINPUT126), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G390), .B1(new_n1041), .B2(new_n1072), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1072), .ZN(new_n1294));
  AOI211_X1 g1094(.A(new_n1294), .B(new_n1138), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1292), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G393), .B(G396), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1292), .B(new_n1297), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  INV_X1    g1102(.A(G213), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1303), .A2(G343), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1256), .A2(new_n777), .B1(new_n1250), .B2(new_n1249), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1253), .A2(new_n1256), .A3(KEYINPUT57), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n721), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G378), .B(new_n1305), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1253), .A2(new_n1256), .A3(new_n1267), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1289), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1304), .B1(new_n1309), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1304), .A2(G2897), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1265), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1153), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1170), .A2(new_n1153), .A3(KEYINPUT60), .A4(new_n1145), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT60), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n772), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1316), .A2(new_n1319), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1323), .A2(G384), .A3(new_n1284), .ZN(new_n1324));
  AOI21_X1  g1124(.A(G384), .B1(new_n1323), .B2(new_n1284), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1315), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1284), .ZN(new_n1327));
  INV_X1    g1127(.A(G384), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1323), .A2(G384), .A3(new_n1284), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1314), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1302), .B1(new_n1313), .B2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1309), .A2(new_n1312), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1304), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1334), .A2(new_n1335), .A3(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1313), .A2(KEYINPUT62), .A3(new_n1337), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1333), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1301), .A2(new_n1342), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1344));
  AOI21_X1  g1144(.A(G378), .B1(new_n1305), .B2(new_n1310), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1345), .B1(new_n1262), .B2(G378), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1344), .B1(new_n1346), .B2(new_n1304), .ZN(new_n1347));
  AOI211_X1 g1147(.A(new_n1304), .B(new_n1336), .C1(new_n1309), .C2(new_n1312), .ZN(new_n1348));
  OAI211_X1 g1148(.A(new_n1347), .B(new_n1302), .C1(new_n1348), .C2(KEYINPUT63), .ZN(new_n1349));
  AND3_X1   g1149(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1337), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1299), .B(new_n1300), .C1(new_n1349), .C2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT127), .ZN(new_n1352));
  AND3_X1   g1152(.A1(new_n1343), .A2(new_n1351), .A3(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1352), .B1(new_n1343), .B2(new_n1351), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1353), .A2(new_n1354), .ZN(G405));
  NAND2_X1  g1155(.A1(G375), .A2(new_n1289), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1309), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1301), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1299), .A2(new_n1300), .A3(new_n1357), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1336), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1359), .A2(new_n1337), .A3(new_n1360), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(G402));
endmodule


