//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  OR4_X1    g031(.A1(G237), .A2(G238), .A3(G236), .A4(G235), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n461), .B1(G2104), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR3_X1   g039(.A1(new_n464), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n465));
  OAI21_X1  g040(.A(G101), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n464), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n462), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(G136), .B2(new_n483), .ZN(G162));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n462), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n467), .A2(new_n489), .A3(G138), .A4(new_n462), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n462), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT69), .A4(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n478), .A2(G126), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n500), .B2(new_n502), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n491), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT71), .B1(new_n508), .B2(G62), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(G75), .B2(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(KEYINPUT71), .A3(G62), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(new_n508), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n512), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n520));
  XOR2_X1   g095(.A(new_n520), .B(KEYINPUT72), .Z(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  INV_X1    g099(.A(G89), .ZN(new_n525));
  OAI221_X1 g100(.A(new_n523), .B1(new_n516), .B2(new_n524), .C1(new_n525), .C2(new_n514), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n521), .A2(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n514), .A2(new_n529), .B1(new_n516), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n507), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(G171));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT5), .B(G543), .Z(new_n536));
  INV_X1    g111(.A(G56), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n507), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n540), .B1(new_n539), .B2(new_n538), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n513), .A2(new_n508), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n513), .A2(G543), .ZN(new_n543));
  AOI22_X1  g118(.A1(G81), .A2(new_n542), .B1(new_n543), .B2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  XNOR2_X1  g126(.A(new_n508), .B(KEYINPUT75), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n507), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n542), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n514), .A2(KEYINPUT74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(G91), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n543), .A2(new_n559), .A3(G53), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n516), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n554), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G166), .ZN(G303));
  INV_X1    g143(.A(G49), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n516), .A2(KEYINPUT77), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT77), .B1(new_n516), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n556), .A2(new_n557), .ZN(new_n575));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  OR3_X1    g151(.A1(new_n575), .A2(KEYINPUT76), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT76), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n536), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(new_n543), .B2(G48), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n575), .B2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(G85), .A2(new_n542), .B1(new_n543), .B2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n507), .B2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n556), .A2(G92), .A3(new_n557), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT10), .Z(new_n592));
  NAND2_X1  g167(.A1(new_n552), .A2(G66), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n507), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(G54), .B2(new_n543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n590), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n590), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G868), .B2(new_n565), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(G868), .B2(new_n565), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n598), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n598), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g184(.A1(new_n463), .A2(new_n465), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n467), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n483), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n478), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n462), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n629), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT78), .Z(new_n641));
  NOR2_X1   g216(.A1(G2072), .A2(G2078), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n444), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(KEYINPUT17), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n639), .B(new_n640), .C1(new_n444), .C2(new_n642), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n645), .A2(new_n641), .A3(new_n639), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  AND2_X1   g236(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT80), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n655), .A2(new_n658), .A3(new_n662), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1981), .B(G1986), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G23), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n579), .B2(new_n673), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT33), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(G22), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G166), .B2(new_n673), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(G1971), .Z(new_n680));
  MUX2_X1   g255(.A(G6), .B(G305), .S(G16), .Z(new_n681));
  XOR2_X1   g256(.A(KEYINPUT32), .B(G1981), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT81), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT34), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  MUX2_X1   g263(.A(G24), .B(G290), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G1986), .Z(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n483), .A2(G131), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n478), .A2(G119), .ZN(new_n694));
  OR2_X1    g269(.A1(G95), .A2(G2105), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n695), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n692), .B1(new_n698), .B2(new_n691), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT35), .B(G1991), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n687), .A2(new_n688), .A3(new_n690), .A4(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT82), .B(KEYINPUT36), .Z(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT94), .B(KEYINPUT23), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n673), .A2(G20), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n565), .B2(new_n673), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1956), .ZN(new_n710));
  OAI21_X1  g285(.A(KEYINPUT89), .B1(G16), .B2(G21), .ZN(new_n711));
  NOR2_X1   g286(.A1(G286), .A2(new_n673), .ZN(new_n712));
  MUX2_X1   g287(.A(new_n711), .B(KEYINPUT89), .S(new_n712), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1966), .ZN(new_n714));
  NOR2_X1   g289(.A1(G29), .A2(G35), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G162), .B2(G29), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G2090), .ZN(new_n719));
  NAND2_X1  g294(.A1(G160), .A2(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(KEYINPUT24), .A2(G34), .ZN(new_n721));
  NOR2_X1   g296(.A1(KEYINPUT24), .A2(G34), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n691), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT85), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT86), .ZN(new_n726));
  INV_X1    g301(.A(G2084), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n714), .A2(new_n719), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n718), .A2(G2090), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT93), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n673), .A2(G19), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n546), .B2(new_n673), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1341), .Z(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT30), .B(G28), .ZN(new_n735));
  OR2_X1    g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  NAND2_X1  g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n735), .A2(new_n691), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n691), .A2(G32), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  AOI22_X1  g317(.A1(G129), .A2(new_n478), .B1(new_n483), .B2(G141), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n610), .A2(G105), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n738), .B1(new_n691), .B2(new_n621), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n750));
  OR3_X1    g325(.A1(new_n750), .A2(G5), .A3(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(G5), .B2(G16), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n751), .B(new_n752), .C1(G301), .C2(new_n673), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n483), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n478), .A2(G128), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n462), .A2(G116), .ZN(new_n757));
  OAI21_X1  g332(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n691), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n734), .A2(new_n749), .A3(new_n754), .A4(new_n765), .ZN(new_n766));
  OR4_X1    g341(.A1(new_n710), .A2(new_n729), .A3(new_n731), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n691), .A2(G27), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n691), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT91), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(new_n443), .ZN(new_n771));
  NOR2_X1   g346(.A1(G29), .A2(G33), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n483), .A2(G139), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT83), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT84), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n467), .A2(G127), .ZN(new_n780));
  INV_X1    g355(.A(G115), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n464), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n779), .B1(G2105), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n772), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(new_n442), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n726), .A2(new_n727), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT87), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n673), .A2(G4), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n598), .B2(new_n673), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n785), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n767), .A2(new_n771), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n704), .A2(new_n705), .A3(new_n793), .ZN(G150));
  INV_X1    g369(.A(G150), .ZN(G311));
  NOR2_X1   g370(.A1(new_n597), .A2(new_n604), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT38), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n542), .A2(G93), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n543), .A2(G55), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(new_n507), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT95), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n802), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n804), .A2(new_n805), .A3(new_n799), .A4(new_n798), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n803), .A2(new_n806), .A3(new_n541), .A4(new_n544), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n803), .A2(new_n806), .B1(new_n541), .B2(new_n544), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n797), .B(new_n810), .Z(new_n811));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n812));
  AOI21_X1  g387(.A(G860), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n812), .B2(new_n811), .ZN(new_n814));
  OAI21_X1  g389(.A(G860), .B1(new_n800), .B2(new_n802), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(G145));
  NAND2_X1  g392(.A1(new_n483), .A2(G142), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n478), .A2(G130), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n462), .A2(G118), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n612), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n697), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT96), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n745), .B(new_n759), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n783), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n783), .A2(new_n826), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n495), .A2(new_n499), .B1(new_n478), .B2(G126), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n491), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n831), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n783), .A2(new_n826), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n827), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n825), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n831), .B1(new_n828), .B2(new_n829), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(new_n833), .A3(new_n827), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(KEYINPUT97), .A3(new_n825), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n841), .A2(new_n825), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(G160), .B(new_n621), .Z(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(G162), .Z(new_n847));
  AOI21_X1  g422(.A(G37), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n838), .B2(new_n842), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(KEYINPUT98), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n839), .A2(new_n840), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(new_n852), .A3(new_n824), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n849), .A2(KEYINPUT99), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT99), .B1(new_n849), .B2(new_n853), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n848), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g432(.A1(new_n800), .A2(new_n802), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(G868), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n606), .B(KEYINPUT100), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n810), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n565), .B1(new_n592), .B2(new_n596), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n592), .A2(new_n565), .A3(new_n596), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n867));
  INV_X1    g442(.A(new_n864), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n862), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(KEYINPUT41), .A3(new_n864), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n866), .B1(new_n871), .B2(new_n861), .ZN(new_n872));
  XNOR2_X1  g447(.A(G290), .B(KEYINPUT101), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n579), .ZN(new_n874));
  XOR2_X1   g449(.A(G166), .B(G305), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT42), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G868), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(new_n872), .B2(new_n878), .ZN(new_n881));
  AOI211_X1 g456(.A(KEYINPUT102), .B(new_n859), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n879), .A2(new_n881), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(KEYINPUT102), .B2(new_n883), .ZN(G295));
  AOI21_X1  g459(.A(new_n882), .B1(KEYINPUT102), .B2(new_n883), .ZN(G331));
  OAI21_X1  g460(.A(G171), .B1(new_n808), .B2(new_n809), .ZN(new_n886));
  INV_X1    g461(.A(new_n809), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(G301), .A3(new_n807), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(G286), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n888), .A3(G168), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n871), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n892), .A2(new_n865), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n871), .A2(new_n892), .A3(KEYINPUT103), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n895), .A2(new_n876), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n892), .A2(new_n865), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n869), .A2(new_n870), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n891), .B2(new_n890), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n902), .B2(KEYINPUT103), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n876), .A4(new_n895), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  INV_X1    g481(.A(new_n876), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n896), .A2(new_n897), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT103), .B1(new_n871), .B2(new_n892), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n899), .A2(new_n905), .A3(new_n906), .A4(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G37), .B1(new_n898), .B2(KEYINPUT104), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n907), .B1(new_n902), .B2(new_n900), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n905), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n913), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT44), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n911), .A2(new_n919), .A3(KEYINPUT43), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n911), .B2(KEYINPUT43), .ZN(new_n921));
  AND4_X1   g496(.A1(new_n912), .A2(new_n914), .A3(new_n905), .A4(new_n915), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n918), .B1(new_n923), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g499(.A1(G160), .A2(G40), .ZN(new_n925));
  AOI21_X1  g500(.A(G1384), .B1(new_n491), .B2(new_n830), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n925), .A2(KEYINPUT45), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n928), .A2(G1986), .A3(G290), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n930));
  INV_X1    g505(.A(G1996), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n745), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n759), .B(new_n764), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n697), .B(new_n700), .Z(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI22_X1  g511(.A1(new_n929), .A2(new_n930), .B1(new_n936), .B2(new_n928), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n930), .B2(new_n929), .ZN(new_n938));
  INV_X1    g513(.A(new_n933), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n927), .B1(new_n939), .B2(new_n745), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n927), .A2(new_n931), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(KEYINPUT46), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT47), .Z(new_n945));
  NAND2_X1  g520(.A1(new_n698), .A2(new_n700), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n934), .A2(new_n946), .B1(G2067), .B2(new_n759), .ZN(new_n947));
  AOI211_X1 g522(.A(new_n938), .B(new_n945), .C1(new_n927), .C2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT127), .ZN(new_n949));
  INV_X1    g524(.A(G8), .ZN(new_n950));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT115), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT115), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n505), .A2(new_n954), .A3(KEYINPUT45), .A4(new_n951), .ZN(new_n955));
  INV_X1    g530(.A(G40), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n470), .A2(new_n473), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n926), .B2(KEYINPUT45), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1966), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n505), .B2(new_n951), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n831), .A2(new_n951), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n957), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n964), .A2(new_n966), .A3(G2084), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n950), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(G286), .A2(G8), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT126), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n969), .A2(KEYINPUT51), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n962), .A2(KEYINPUT125), .A3(new_n968), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT125), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n958), .B1(new_n952), .B2(KEYINPUT115), .ZN(new_n975));
  AOI21_X1  g550(.A(G1966), .B1(new_n975), .B2(new_n955), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n976), .B2(new_n967), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n977), .A3(new_n971), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n978), .A2(KEYINPUT51), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n973), .A2(new_n977), .A3(G8), .ZN(new_n980));
  INV_X1    g555(.A(new_n971), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n949), .B(new_n972), .C1(new_n979), .C2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(KEYINPUT51), .A3(new_n978), .ZN(new_n984));
  INV_X1    g559(.A(new_n972), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT127), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT62), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n980), .A2(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n978), .A2(KEYINPUT51), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n949), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT62), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(KEYINPUT127), .A3(new_n985), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n579), .A2(G1976), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n925), .A2(new_n965), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(new_n950), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n579), .B2(G1976), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n584), .B1(new_n585), .B2(new_n514), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G1981), .ZN(new_n1003));
  INV_X1    g578(.A(G1981), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n584), .C1(new_n575), .C2(new_n585), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(KEYINPUT49), .A3(new_n1005), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n997), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n1011), .B(new_n574), .C1(new_n577), .C2(new_n578), .ZN(new_n1012));
  INV_X1    g587(.A(new_n997), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT52), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1001), .A2(new_n1010), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n925), .B1(KEYINPUT45), .B2(new_n926), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n505), .A2(new_n951), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n957), .B1(new_n965), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n505), .A2(new_n951), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT106), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT107), .B(G1971), .Z(new_n1026));
  NAND3_X1  g601(.A1(new_n1020), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n964), .A2(new_n966), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1029), .A2(G2090), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n950), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G166), .A2(new_n950), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1015), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n957), .B1(new_n926), .B2(new_n963), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n505), .A2(new_n963), .A3(new_n951), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n957), .B(KEYINPUT113), .C1(new_n926), .C2(new_n963), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(G2090), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1027), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n950), .B1(new_n1046), .B2(KEYINPUT114), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1027), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1034), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1029), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1053));
  AOI21_X1  g628(.A(G2078), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1054));
  OAI221_X1 g629(.A(new_n1052), .B1(new_n960), .B2(new_n1053), .C1(new_n1054), .C2(KEYINPUT53), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G171), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1038), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n987), .A2(new_n994), .A3(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n969), .A2(G168), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1037), .B(new_n1059), .C1(new_n1060), .C2(new_n1034), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT63), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1001), .A2(KEYINPUT110), .A3(new_n1010), .A4(new_n1014), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT110), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1014), .A2(new_n1010), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n998), .A2(new_n1000), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1036), .A2(new_n1031), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1069), .A2(KEYINPUT63), .A3(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(new_n1059), .C1(new_n1034), .C2(new_n1031), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1005), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G288), .A2(G1976), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n1010), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1075), .A2(KEYINPUT111), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(KEYINPUT111), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n997), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1069), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n1070), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1078), .B(KEYINPUT112), .C1(new_n1079), .C2(new_n1070), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1063), .A2(new_n1072), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1058), .A2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT116), .B(G1956), .Z(new_n1086));
  NAND2_X1  g661(.A1(new_n1044), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1024), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n564), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(new_n1091), .C1(new_n507), .C2(new_n553), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT57), .B1(new_n554), .B2(new_n564), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1087), .A2(new_n1089), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1044), .A2(new_n1086), .B1(new_n1024), .B2(new_n1088), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(KEYINPUT117), .A3(new_n1094), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1094), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1097), .A2(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1016), .B(new_n931), .C1(new_n1017), .C2(KEYINPUT45), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT121), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1024), .A2(new_n1108), .A3(new_n931), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n996), .A2(KEYINPUT118), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n996), .A2(KEYINPUT118), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1105), .B1(new_n1114), .B2(new_n546), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1114), .A2(new_n1105), .A3(new_n546), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1102), .A2(new_n1104), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1095), .A2(KEYINPUT61), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1101), .B1(new_n1098), .B2(KEYINPUT119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1100), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1094), .B1(new_n1100), .B2(new_n1121), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1098), .A2(KEYINPUT119), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(KEYINPUT120), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1118), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT123), .B1(new_n1117), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1118), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1120), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT117), .B1(new_n1098), .B2(new_n1094), .ZN(new_n1134));
  AND4_X1   g709(.A1(KEYINPUT117), .A2(new_n1087), .A3(new_n1089), .A4(new_n1094), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1114), .A2(new_n546), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1114), .A2(new_n1105), .A3(new_n546), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1136), .A2(new_n1103), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1132), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(G2067), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n790), .B2(new_n1029), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT60), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(new_n598), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(KEYINPUT60), .B2(new_n1144), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1128), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1130), .A2(new_n1131), .B1(new_n597), .B2(new_n1144), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1038), .A2(new_n1050), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1054), .A2(KEYINPUT53), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1051), .B2(new_n1029), .ZN(new_n1155));
  XOR2_X1   g730(.A(G171), .B(KEYINPUT54), .Z(new_n1156));
  AOI21_X1  g731(.A(new_n1053), .B1(new_n926), .B2(KEYINPUT45), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n959), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1155), .A2(new_n1158), .B1(new_n1055), .B2(new_n1156), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1153), .B(new_n1159), .C1(new_n983), .C2(new_n986), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(KEYINPUT124), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1085), .B1(new_n1152), .B2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(G290), .B(G1986), .Z(new_n1164));
  AOI21_X1  g739(.A(new_n928), .B1(new_n936), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n948), .B1(new_n1163), .B2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g741(.A1(new_n652), .A2(G319), .ZN(new_n1168));
  NOR3_X1   g742(.A1(G229), .A2(G401), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n856), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n923), .A2(new_n1170), .ZN(G308));
  OR2_X1    g745(.A1(new_n921), .A2(new_n922), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n856), .B(new_n1169), .C1(new_n1172), .C2(new_n920), .ZN(G225));
endmodule


