//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  AOI21_X1  g011(.A(G146), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n190), .B(new_n193), .C1(new_n198), .C2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n195), .A2(new_n197), .A3(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G143), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n191), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n200), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G146), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n190), .B1(new_n208), .B2(new_n193), .ZN(new_n209));
  OAI21_X1  g023(.A(G125), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n202), .A2(G128), .A3(new_n213), .A4(new_n203), .ZN(new_n214));
  INV_X1    g028(.A(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n195), .A2(new_n197), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n200), .B1(new_n216), .B2(new_n199), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(new_n203), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n214), .B(new_n215), .C1(new_n217), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G224), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G953), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT7), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G110), .B(G122), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n228), .B(KEYINPUT8), .Z(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  INV_X1    g044(.A(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G107), .ZN(new_n232));
  INV_X1    g046(.A(G107), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT3), .A3(G104), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT74), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n233), .B2(G104), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(KEYINPUT74), .A3(G107), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(new_n236), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n231), .A2(G107), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n233), .A2(G104), .ZN(new_n242));
  OAI21_X1  g056(.A(G101), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G113), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G119), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT5), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G119), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G116), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(G119), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT5), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n245), .A2(KEYINPUT2), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G113), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G116), .B(G119), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n244), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n249), .A2(new_n253), .B1(new_n259), .B2(new_n258), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n240), .A3(new_n243), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n229), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI211_X1 g081(.A(KEYINPUT83), .B(new_n229), .C1(new_n262), .C2(new_n264), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n227), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT82), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n210), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n193), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT65), .B1(new_n217), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n204), .A3(new_n201), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT82), .A3(G125), .ZN(new_n275));
  INV_X1    g089(.A(new_n203), .ZN(new_n276));
  OAI21_X1  g090(.A(G128), .B1(new_n213), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n207), .B2(G146), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n219), .A2(new_n218), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n208), .A2(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n226), .B1(new_n280), .B2(new_n215), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n271), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n189), .B1(new_n269), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n233), .A2(KEYINPUT3), .A3(G104), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT3), .B1(new_n233), .B2(G104), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n238), .B(new_n239), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n236), .A2(KEYINPUT75), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n240), .A2(KEYINPUT4), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n287), .A2(KEYINPUT4), .A3(new_n288), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n258), .A2(new_n259), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n260), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n264), .B(new_n228), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n265), .B(new_n266), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n296), .A2(KEYINPUT84), .A3(new_n282), .A4(new_n227), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n284), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n271), .A2(new_n275), .A3(new_n221), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n224), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n271), .A2(new_n275), .A3(new_n221), .A4(new_n225), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n228), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n240), .A2(KEYINPUT4), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n287), .A2(new_n288), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n287), .A2(KEYINPUT4), .A3(new_n288), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n294), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n264), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT6), .A3(new_n295), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n313), .B(new_n304), .C1(new_n309), .C2(new_n310), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n299), .B1(new_n303), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n188), .B1(new_n298), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n312), .A2(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n301), .A2(new_n302), .ZN(new_n319));
  AOI21_X1  g133(.A(G902), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n284), .A2(new_n297), .A3(new_n295), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n187), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n317), .A2(KEYINPUT85), .A3(new_n322), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n320), .A2(new_n321), .A3(new_n187), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT85), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(G113), .B(G122), .Z(new_n329));
  XOR2_X1   g143(.A(KEYINPUT90), .B(G104), .Z(new_n330));
  XOR2_X1   g144(.A(new_n329), .B(new_n330), .Z(new_n331));
  INV_X1    g145(.A(G237), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G214), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n195), .B(new_n197), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(G143), .A2(G214), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT86), .ZN(new_n338));
  NOR2_X1   g152(.A1(G237), .A2(G953), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n338), .B1(new_n337), .B2(new_n339), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT18), .A2(G131), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n199), .ZN(new_n346));
  INV_X1    g160(.A(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n215), .A2(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G146), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n342), .A2(new_n344), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n343), .B(KEYINPUT87), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(new_n336), .C1(new_n340), .C2(new_n341), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n342), .A2(G131), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n357));
  INV_X1    g171(.A(G131), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n336), .B(new_n358), .C1(new_n340), .C2(new_n341), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT16), .ZN(new_n361));
  OR3_X1    g175(.A1(new_n215), .A2(KEYINPUT16), .A3(G140), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(G146), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G146), .B1(new_n361), .B2(new_n362), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n342), .A2(KEYINPUT17), .A3(G131), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n331), .B(new_n355), .C1(new_n360), .C2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n356), .A2(new_n359), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n366), .B(new_n367), .C1(new_n371), .C2(KEYINPUT17), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n331), .B1(new_n372), .B2(new_n355), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n299), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G475), .ZN(new_n375));
  INV_X1    g189(.A(new_n331), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT19), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT88), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n377), .B1(new_n350), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n345), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n364), .B1(new_n381), .B2(new_n199), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n371), .A2(new_n382), .B1(new_n352), .B2(new_n354), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n376), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n371), .A2(new_n382), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n386), .A2(new_n384), .A3(new_n355), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n369), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n389));
  NOR2_X1   g203(.A1(G475), .A2(G902), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n375), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT91), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n386), .A2(new_n355), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n331), .B1(new_n396), .B2(KEYINPUT89), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n383), .A2(new_n384), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n370), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n390), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n391), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT91), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n375), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT15), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G478), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT9), .B(G234), .ZN(new_n407));
  INV_X1    g221(.A(G217), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n407), .A2(new_n408), .A3(G953), .ZN(new_n409));
  XNOR2_X1  g223(.A(G116), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n233), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n207), .A2(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n218), .A2(G143), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n412), .A2(KEYINPUT13), .A3(new_n413), .ZN(new_n415));
  OAI21_X1  g229(.A(G134), .B1(new_n412), .B2(KEYINPUT13), .ZN(new_n416));
  OAI221_X1 g230(.A(new_n411), .B1(new_n414), .B2(G134), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n246), .A2(G122), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n233), .B1(new_n418), .B2(KEYINPUT14), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(new_n410), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n414), .A2(G134), .ZN(new_n421));
  INV_X1    g235(.A(G134), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n412), .B2(new_n413), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n420), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n409), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n424), .A3(new_n409), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n406), .B1(new_n428), .B2(new_n299), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n299), .A3(new_n406), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(G234), .A2(G237), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n433), .A2(G952), .A3(new_n333), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n433), .A2(G902), .A3(G953), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(G898), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n395), .A2(new_n404), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n328), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G137), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT72), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT23), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(KEYINPUT23), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n218), .A2(G119), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G119), .B(G128), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n449), .B1(new_n450), .B2(new_n446), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G110), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT24), .B(G110), .Z(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n450), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n452), .B(new_n454), .C1(new_n364), .C2(new_n365), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n363), .A2(new_n346), .ZN(new_n456));
  INV_X1    g270(.A(G110), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n449), .B(new_n457), .C1(new_n450), .C2(new_n446), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n453), .A2(new_n450), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n455), .B1(new_n460), .B2(KEYINPUT73), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n363), .A3(new_n346), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT73), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n444), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n464), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n460), .A2(KEYINPUT73), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n455), .A4(new_n443), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n466), .A2(new_n299), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n466), .A2(KEYINPUT25), .A3(new_n469), .A4(new_n299), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n408), .B1(G234), .B2(new_n299), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n466), .A2(new_n469), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n475), .A2(G902), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT71), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT31), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT11), .B1(new_n422), .B2(G137), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT11), .ZN(new_n484));
  INV_X1    g298(.A(G137), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(G134), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT66), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n485), .B2(G134), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n422), .A2(KEYINPUT66), .A3(G137), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n487), .A2(new_n358), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n422), .A2(G137), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n485), .A2(G134), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n214), .B1(new_n217), .B2(new_n220), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n293), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n483), .A2(new_n486), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n489), .A2(new_n490), .ZN(new_n500));
  OAI21_X1  g314(.A(G131), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n491), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n502), .A2(new_n273), .A3(new_n204), .A4(new_n201), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n332), .A2(new_n333), .A3(G210), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT27), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT26), .B(G101), .Z(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT68), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n511), .B(new_n508), .C1(new_n498), .C2(new_n503), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n496), .A2(new_n497), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n503), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT30), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n503), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n294), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n482), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n501), .A2(new_n491), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n274), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n294), .B1(new_n280), .B2(new_n495), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n509), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n511), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n504), .A2(KEYINPUT68), .A3(new_n509), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n518), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n517), .B1(new_n503), .B2(new_n514), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n293), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(KEYINPUT31), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n504), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n294), .B1(new_n503), .B2(new_n514), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT28), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n503), .A2(KEYINPUT70), .A3(new_n514), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT70), .B1(new_n503), .B2(new_n514), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n536), .A2(new_n537), .A3(new_n293), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n534), .B1(new_n538), .B2(KEYINPUT28), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n508), .B(KEYINPUT69), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n520), .A2(new_n531), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(G472), .A2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n481), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n293), .B1(new_n515), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT28), .B1(new_n546), .B2(new_n535), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  INV_X1    g362(.A(new_n533), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n549), .B2(new_n504), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n540), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n513), .A2(new_n482), .A3(new_n519), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT31), .B1(new_n527), .B2(new_n530), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(KEYINPUT71), .A3(new_n542), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT32), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n544), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n520), .A2(new_n531), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n543), .B1(new_n558), .B2(new_n551), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT29), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n508), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n534), .B(new_n561), .C1(new_n538), .C2(KEYINPUT28), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n516), .A2(new_n518), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n532), .B1(new_n563), .B2(new_n293), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n560), .B1(new_n564), .B2(new_n509), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n547), .A2(new_n550), .A3(new_n540), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n562), .B(new_n299), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n559), .A2(KEYINPUT32), .B1(new_n567), .B2(G472), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n480), .B1(new_n557), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G221), .B1(new_n407), .B2(G902), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G140), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n333), .A2(G227), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n240), .A2(new_n243), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT79), .B1(new_n579), .B2(new_n497), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT79), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n280), .A2(new_n581), .A3(new_n244), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n196), .A2(G143), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n194), .A2(KEYINPUT64), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n199), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n218), .B1(new_n586), .B2(KEYINPUT1), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n214), .B1(new_n587), .B2(new_n278), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT77), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n579), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n579), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT77), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n583), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n521), .A2(KEYINPUT78), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n578), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n588), .A2(new_n589), .A3(new_n579), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n589), .B1(new_n588), .B2(new_n579), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n580), .B(new_n582), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n577), .A3(new_n594), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT76), .B1(new_n291), .B2(new_n274), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n205), .A2(new_n209), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT76), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n603), .B(new_n604), .C1(new_n289), .C2(new_n290), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n597), .B2(new_n598), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n497), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n606), .A2(new_n608), .A3(new_n521), .A4(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n574), .B1(new_n601), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n502), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n613), .A2(new_n574), .A3(new_n610), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT80), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT80), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n574), .A3(new_n610), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n600), .A2(new_n596), .B1(new_n618), .B2(new_n521), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n616), .B(new_n617), .C1(new_n619), .C2(new_n574), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n615), .A2(G469), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT81), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n599), .A2(new_n577), .A3(new_n594), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n577), .B1(new_n599), .B2(new_n594), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n610), .A2(new_n574), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n596), .A2(KEYINPUT81), .A3(new_n600), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n613), .A2(new_n610), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n573), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(G469), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n299), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n299), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n621), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n440), .A2(new_n569), .A3(new_n570), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  OAI21_X1  g452(.A(G472), .B1(new_n541), .B2(G902), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n544), .A2(new_n639), .A3(new_n555), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n480), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n641), .A2(new_n636), .A3(new_n642), .A4(new_n570), .ZN(new_n643));
  INV_X1    g457(.A(new_n427), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n425), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(G902), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT92), .B1(new_n646), .B2(G478), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT92), .ZN(new_n648));
  INV_X1    g462(.A(G478), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n648), .B(new_n649), .C1(new_n645), .C2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n428), .B(KEYINPUT33), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n649), .A2(G902), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n403), .B1(new_n402), .B2(new_n375), .ZN(new_n656));
  INV_X1    g470(.A(G475), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n355), .B1(new_n360), .B2(new_n368), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n376), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n369), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n657), .B1(new_n660), .B2(new_n299), .ZN(new_n661));
  AOI211_X1 g475(.A(KEYINPUT91), .B(new_n661), .C1(new_n401), .C2(new_n391), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n655), .B1(new_n656), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n437), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n187), .B1(new_n320), .B2(new_n321), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n327), .B(new_n664), .C1(new_n324), .C2(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n643), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT34), .B(G104), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NAND3_X1  g483(.A1(new_n401), .A2(KEYINPUT93), .A3(new_n391), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT93), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n388), .A2(new_n671), .A3(new_n389), .A4(new_n390), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(new_n375), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n432), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n643), .A2(new_n666), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT35), .B(G107), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n461), .A2(new_n465), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n444), .A2(KEYINPUT36), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n679), .B(new_n680), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n478), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n476), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n640), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n440), .A2(new_n570), .A3(new_n636), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  INV_X1    g502(.A(new_n327), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n317), .B2(new_n322), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n434), .B1(new_n435), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n432), .A2(new_n670), .A3(new_n673), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n690), .A2(new_n694), .A3(new_n683), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n557), .B2(new_n568), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n636), .A2(new_n570), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT94), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n327), .B(new_n683), .C1(new_n324), .C2(new_n665), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n670), .A2(new_n673), .A3(new_n432), .A4(new_n693), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n557), .A2(new_n568), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n636), .A2(new_n570), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT94), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  NOR2_X1   g522(.A1(new_n513), .A2(new_n519), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n549), .A2(new_n504), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(new_n540), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n299), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n559), .A2(KEYINPUT32), .B1(G472), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n557), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT95), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n323), .A2(new_n326), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT38), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n395), .A2(new_n404), .B1(new_n430), .B2(new_n431), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n327), .A3(new_n684), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n692), .B(KEYINPUT39), .Z(new_n721));
  NAND2_X1  g535(.A1(new_n697), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n216), .ZN(G45));
  OAI21_X1  g540(.A(KEYINPUT96), .B1(new_n663), .B2(new_n692), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n647), .A2(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n395), .B2(new_n404), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT96), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n693), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n700), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n703), .A2(new_n636), .A3(new_n570), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G146), .ZN(G48));
  AOI21_X1  g551(.A(new_n632), .B1(new_n631), .B2(new_n299), .ZN(new_n738));
  AOI211_X1 g552(.A(G469), .B(G902), .C1(new_n628), .C2(new_n630), .ZN(new_n739));
  INV_X1    g553(.A(new_n570), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n663), .A2(new_n666), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n569), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT41), .B(G113), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G15));
  NOR2_X1   g559(.A1(new_n666), .A2(new_n675), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n569), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR2_X1   g562(.A1(new_n439), .A2(new_n684), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n741), .A2(new_n703), .A3(new_n690), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  OAI21_X1  g565(.A(new_n432), .B1(new_n656), .B2(new_n662), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n666), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n554), .A2(new_n542), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n639), .A2(new_n642), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n741), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT97), .B(G122), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G24));
  AND2_X1   g572(.A1(new_n727), .A2(new_n731), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n631), .A2(new_n299), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(G469), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n570), .A3(new_n633), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n327), .B1(new_n324), .B2(new_n665), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n639), .A2(new_n754), .A3(new_n683), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT98), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n639), .A2(new_n754), .A3(KEYINPUT98), .A4(new_n683), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n759), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n727), .A2(new_n731), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n569), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n610), .B1(new_n623), .B2(new_n624), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n775), .A2(new_n573), .B1(new_n626), .B2(new_n613), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n634), .B1(new_n776), .B2(G469), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n740), .B1(new_n633), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n689), .B1(new_n323), .B2(new_n326), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n773), .A2(new_n774), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n780), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n754), .A2(new_n556), .ZN(new_n783));
  AOI211_X1 g597(.A(KEYINPUT99), .B(new_n480), .C1(new_n568), .C2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT99), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n568), .A2(new_n783), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n786), .B2(new_n642), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n759), .B(new_n782), .C1(new_n784), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n781), .B1(new_n788), .B2(KEYINPUT42), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NAND4_X1  g604(.A1(new_n569), .A2(new_n694), .A3(new_n779), .A4(new_n778), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  NOR2_X1   g606(.A1(new_n656), .A2(new_n662), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n655), .ZN(new_n794));
  NAND2_X1  g608(.A1(KEYINPUT100), .A2(KEYINPUT43), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(new_n655), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n640), .A3(new_n683), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n779), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT101), .Z(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT45), .B1(new_n615), .B2(new_n620), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n776), .A2(KEYINPUT45), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(G469), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n804), .B1(new_n808), .B2(new_n634), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT46), .B(new_n635), .C1(new_n805), .C2(new_n807), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n633), .A3(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n811), .A2(new_n570), .A3(new_n721), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n800), .A2(new_n801), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n803), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT102), .B(G137), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(G39));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n570), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n811), .A2(KEYINPUT47), .A3(new_n570), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n716), .A2(new_n327), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n703), .A3(new_n642), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n759), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n752), .A2(new_n763), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n476), .A2(new_n682), .A3(new_n693), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT109), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT109), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n476), .A2(new_n682), .A3(new_n831), .A4(new_n693), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n828), .A2(new_n714), .A3(new_n778), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n833), .A2(new_n718), .A3(new_n690), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(KEYINPUT110), .A3(new_n714), .A4(new_n778), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n736), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT94), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n770), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n827), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n767), .A2(new_n768), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n732), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n764), .A2(new_n846), .B1(new_n699), .B2(new_n706), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n836), .A2(new_n838), .B1(new_n733), .B2(new_n735), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(KEYINPUT52), .A3(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n569), .B(new_n741), .C1(new_n742), .C2(new_n746), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n750), .A3(new_n756), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT106), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT106), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n851), .A2(new_n750), .A3(new_n854), .A4(new_n756), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT107), .ZN(new_n857));
  INV_X1    g671(.A(new_n431), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n429), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n430), .A2(KEYINPUT107), .A3(new_n431), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n404), .A3(new_n395), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n437), .B1(new_n862), .B2(new_n663), .ZN(new_n863));
  INV_X1    g677(.A(new_n328), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n637), .B(new_n686), .C1(new_n643), .C2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n769), .A2(new_n731), .A3(new_n727), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n791), .B1(new_n867), .B2(new_n780), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n670), .A2(new_n673), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n861), .A2(new_n684), .A3(new_n870), .A4(new_n692), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n735), .A2(KEYINPUT108), .A3(new_n779), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT108), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n779), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n734), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n856), .A2(new_n869), .A3(new_n789), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n826), .B1(new_n850), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT112), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n844), .A2(new_n849), .ZN(new_n881));
  INV_X1    g695(.A(new_n852), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n789), .A2(KEYINPUT53), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT111), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n872), .A2(new_n875), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n865), .A2(new_n643), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n759), .A2(new_n769), .A3(new_n782), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n697), .B(new_n440), .C1(new_n569), .C2(new_n685), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n791), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n885), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n869), .A2(KEYINPUT111), .A3(new_n876), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n881), .A2(new_n884), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n877), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n881), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n891), .A2(new_n892), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n883), .B1(new_n844), .B2(new_n849), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n897), .A2(new_n826), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n879), .B1(new_n900), .B2(new_n880), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n896), .A2(KEYINPUT53), .A3(new_n881), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n880), .B1(new_n878), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n895), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n762), .A2(new_n822), .A3(KEYINPUT116), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT116), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n741), .B2(new_n779), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n799), .B(new_n434), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n787), .A2(new_n784), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT48), .Z(new_n912));
  OAI21_X1  g726(.A(new_n434), .B1(new_n906), .B2(new_n908), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n715), .A2(new_n642), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT118), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n434), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT116), .B1(new_n762), .B2(new_n822), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n741), .A2(new_n907), .A3(new_n779), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n642), .A4(new_n715), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n729), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(G952), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n799), .A2(new_n434), .A3(new_n755), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n923), .B(G953), .C1(new_n924), .C2(new_n764), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n912), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n655), .A2(new_n656), .A3(new_n662), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n915), .A2(new_n921), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT117), .B1(new_n909), .B2(new_n845), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n919), .A2(new_n930), .A3(new_n769), .A4(new_n799), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT114), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT113), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n741), .A2(new_n936), .A3(new_n689), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n717), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n741), .B2(new_n689), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n939), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(KEYINPUT114), .A3(new_n717), .A4(new_n937), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n942), .A3(new_n924), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT115), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT50), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT50), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n761), .A2(new_n633), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT104), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n950), .A2(new_n740), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n779), .B(new_n924), .C1(new_n821), .C2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n934), .A2(new_n945), .A3(new_n948), .A4(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT51), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n926), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT120), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT119), .B1(new_n928), .B2(new_n932), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n928), .A2(new_n932), .A3(KEYINPUT119), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n948), .A2(new_n952), .A3(KEYINPUT51), .A4(new_n945), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n956), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n928), .A2(new_n932), .A3(KEYINPUT119), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n957), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n965), .A2(new_n961), .A3(KEYINPUT120), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n955), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  OAI22_X1  g781(.A1(new_n905), .A2(new_n967), .B1(G952), .B2(G953), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT49), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n950), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT105), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n480), .A2(new_n740), .A3(new_n689), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT103), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(new_n794), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n715), .A2(new_n974), .A3(new_n717), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n971), .B(new_n975), .C1(new_n969), .C2(new_n950), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n968), .A2(new_n976), .ZN(G75));
  NOR2_X1   g791(.A1(new_n333), .A2(G952), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n299), .B1(new_n878), .B2(new_n893), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT56), .B1(new_n980), .B2(G210), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n315), .B(new_n319), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT55), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n979), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n983), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT121), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n981), .A2(KEYINPUT121), .A3(new_n983), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(G51));
  XNOR2_X1  g803(.A(new_n634), .B(KEYINPUT57), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n877), .B1(new_n844), .B2(new_n849), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n893), .B(new_n880), .C1(new_n991), .C2(KEYINPUT53), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n880), .B1(new_n878), .B2(new_n893), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n631), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n808), .B(KEYINPUT122), .Z(new_n997));
  NAND2_X1  g811(.A1(new_n980), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n978), .B1(new_n996), .B2(new_n998), .ZN(G54));
  NAND2_X1  g813(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT123), .Z(new_n1001));
  AOI21_X1  g815(.A(new_n388), .B1(new_n980), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n980), .A2(new_n388), .A3(new_n1001), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT124), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n980), .A2(KEYINPUT124), .A3(new_n388), .A4(new_n1001), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n978), .B(new_n1002), .C1(new_n1005), .C2(new_n1006), .ZN(G60));
  NAND2_X1  g821(.A1(G478), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT59), .Z(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n992), .A2(KEYINPUT112), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n894), .B(new_n1010), .C1(new_n1011), .C2(new_n903), .ZN(new_n1012));
  INV_X1    g826(.A(new_n652), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1013), .A2(new_n1009), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n893), .ZN(new_n1017));
  AOI21_X1  g831(.A(KEYINPUT53), .B1(new_n896), .B2(new_n881), .ZN(new_n1018));
  OAI21_X1  g832(.A(KEYINPUT54), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1016), .B1(new_n1019), .B2(new_n992), .ZN(new_n1020));
  OAI21_X1  g834(.A(KEYINPUT125), .B1(new_n1020), .B2(new_n978), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n993), .B2(new_n994), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT125), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1022), .A2(new_n1023), .A3(new_n979), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1014), .A2(new_n1021), .A3(new_n1024), .ZN(G63));
  NAND2_X1  g839(.A1(G217), .A2(G902), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT60), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n681), .B(new_n1028), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n900), .A2(new_n1027), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n979), .B(new_n1029), .C1(new_n1030), .C2(new_n477), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT61), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(G66));
  AOI21_X1  g847(.A(new_n866), .B1(new_n853), .B2(new_n855), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT126), .Z(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n333), .ZN(new_n1036));
  OAI21_X1  g850(.A(G953), .B1(new_n436), .B2(new_n223), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n315), .B1(G898), .B2(new_n333), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(G69));
  NAND3_X1  g854(.A1(new_n725), .A2(new_n736), .A3(new_n847), .ZN(new_n1041));
  OR2_X1    g855(.A1(new_n1041), .A2(KEYINPUT62), .ZN(new_n1042));
  AND2_X1   g856(.A1(new_n862), .A2(new_n663), .ZN(new_n1043));
  NOR4_X1   g857(.A1(new_n722), .A2(new_n774), .A3(new_n822), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1044), .B1(new_n1041), .B2(KEYINPUT62), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n814), .A2(new_n1042), .A3(new_n824), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n333), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n563), .B(new_n381), .Z(new_n1048));
  NAND2_X1  g862(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AND4_X1   g863(.A1(new_n736), .A2(new_n789), .A3(new_n791), .A4(new_n847), .ZN(new_n1050));
  OAI211_X1 g864(.A(new_n812), .B(new_n828), .C1(new_n784), .C2(new_n787), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n1052), .A2(new_n814), .A3(new_n333), .A4(new_n824), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1048), .B1(G900), .B2(G953), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n333), .B1(G227), .B2(G900), .ZN(new_n1055));
  AOI22_X1  g869(.A1(new_n1053), .A2(new_n1054), .B1(KEYINPUT127), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1049), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1055), .A2(KEYINPUT127), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g873(.A(new_n1057), .B(new_n1059), .ZN(G72));
  NAND2_X1  g874(.A1(G472), .A2(G902), .ZN(new_n1061));
  XOR2_X1   g875(.A(new_n1061), .B(KEYINPUT63), .Z(new_n1062));
  NAND3_X1  g876(.A1(new_n1052), .A2(new_n814), .A3(new_n824), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n1062), .B1(new_n1063), .B2(new_n1035), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1064), .A2(new_n508), .A3(new_n564), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n878), .A2(new_n902), .ZN(new_n1066));
  NOR2_X1   g880(.A1(new_n564), .A2(new_n509), .ZN(new_n1067));
  OAI211_X1 g881(.A(new_n1066), .B(new_n1062), .C1(new_n709), .C2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g882(.A1(new_n1065), .A2(new_n1068), .A3(new_n979), .ZN(new_n1069));
  OAI21_X1  g883(.A(new_n1062), .B1(new_n1046), .B2(new_n1035), .ZN(new_n1070));
  NOR2_X1   g884(.A1(new_n564), .A2(new_n508), .ZN(new_n1071));
  AOI21_X1  g885(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(G57));
endmodule


