//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  OR3_X1    g012(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n199), .A2(new_n200), .B1(KEYINPUT2), .B2(G113), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n189), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n193), .A2(new_n197), .A3(new_n201), .A4(KEYINPUT71), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(new_n202), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G137), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT11), .B1(new_n208), .B2(G134), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n209), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n210), .B2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n209), .A2(new_n211), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n212), .A2(new_n213), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(new_n225), .B2(G143), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n232), .A2(new_n235), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n208), .A2(G134), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n222), .B1(new_n239), .B2(new_n211), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT1), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n228), .A2(G146), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n231), .A3(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n226), .A2(new_n229), .B1(G143), .B2(new_n225), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n242), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n241), .A2(new_n223), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n207), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT30), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT30), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n251), .B1(new_n257), .B2(new_n207), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n188), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n251), .A2(KEYINPUT28), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n264), .B(KEYINPUT72), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n207), .A2(new_n250), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT73), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n207), .A2(new_n271), .A3(new_n250), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n251), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n267), .B(new_n268), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT29), .ZN(new_n276));
  INV_X1    g090(.A(new_n264), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n203), .A2(new_n204), .B1(new_n202), .B2(new_n198), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n255), .B2(new_n256), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT74), .B(new_n277), .C1(new_n279), .C2(new_n251), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n265), .A2(new_n275), .A3(new_n276), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n238), .A3(new_n249), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n269), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n266), .B1(new_n283), .B2(KEYINPUT28), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n277), .A2(new_n276), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n187), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n257), .A2(new_n207), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n282), .A3(new_n264), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n258), .A2(KEYINPUT31), .A3(new_n264), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n267), .B1(new_n273), .B2(new_n274), .ZN(new_n293));
  INV_X1    g107(.A(new_n268), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT32), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n294), .ZN(new_n299));
  INV_X1    g113(.A(new_n292), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT31), .B1(new_n258), .B2(new_n264), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT32), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(new_n296), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n287), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G217), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(G234), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G125), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT75), .A3(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(KEYINPUT16), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT16), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n314), .B2(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G146), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n311), .A2(new_n225), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n190), .A2(G128), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n190), .A2(G128), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT24), .B(G110), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n242), .A2(KEYINPUT23), .A3(G119), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n329), .B(new_n324), .C1(new_n322), .C2(KEYINPUT23), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n326), .A2(new_n328), .B1(new_n330), .B2(G110), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n321), .A3(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(KEYINPUT76), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n316), .A2(new_n225), .A3(new_n318), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n320), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n326), .A2(new_n328), .B1(G110), .B2(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(KEYINPUT76), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT77), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT22), .B(G137), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n333), .A2(new_n343), .A3(new_n337), .A4(new_n338), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n310), .B1(new_n347), .B2(G902), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n345), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n346), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n309), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n347), .A2(G902), .A3(new_n308), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n305), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G110), .B(G122), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G107), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(G104), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(KEYINPUT3), .ZN(new_n360));
  INV_X1    g174(.A(G104), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G107), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n358), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT79), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(KEYINPUT79), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n357), .A2(G104), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G101), .ZN(new_n371));
  INV_X1    g185(.A(G101), .ZN(new_n372));
  INV_X1    g186(.A(new_n358), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n360), .A2(new_n362), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n368), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n372), .B1(new_n363), .B2(new_n368), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n278), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G101), .B1(new_n362), .B2(new_n358), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n193), .A2(new_n197), .A3(KEYINPUT5), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n191), .A2(KEYINPUT5), .ZN(new_n383));
  INV_X1    g197(.A(G113), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n205), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n356), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n203), .A2(new_n204), .B1(new_n382), .B2(new_n385), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n381), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n390), .B(new_n355), .C1(new_n278), .C2(new_n378), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n391), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n248), .A2(G125), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n314), .B2(new_n237), .ZN(new_n394));
  INV_X1    g208(.A(G224), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G953), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT85), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n394), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n399), .B(new_n356), .C1(new_n379), .C2(new_n387), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n392), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT7), .B1(new_n395), .B2(G953), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n402), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n393), .B(new_n404), .C1(new_n314), .C2(new_n237), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n378), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n207), .A2(new_n407), .B1(new_n389), .B2(new_n381), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n406), .B1(new_n408), .B2(new_n355), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n355), .B(KEYINPUT8), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n389), .A2(new_n381), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(new_n387), .ZN(new_n412));
  AOI21_X1  g226(.A(G902), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G210), .B1(G237), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n401), .A2(new_n415), .A3(new_n413), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G214), .B1(G237), .B2(G902), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n259), .A2(new_n260), .A3(G214), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(G143), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(G131), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OR3_X1    g241(.A1(new_n424), .A2(new_n426), .A3(new_n222), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n427), .A2(new_n320), .A3(new_n334), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G113), .B(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT86), .B(G104), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n430), .B(new_n431), .Z(new_n432));
  NAND2_X1  g246(.A1(KEYINPUT18), .A2(G131), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n424), .B(new_n433), .Z(new_n434));
  NAND2_X1  g248(.A1(new_n313), .A2(new_n315), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n321), .B1(new_n435), .B2(new_n225), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n424), .B(new_n222), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n311), .A2(KEYINPUT19), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n435), .B2(KEYINPUT19), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n439), .B(new_n320), .C1(G146), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n437), .ZN(new_n443));
  INV_X1    g257(.A(new_n432), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(G475), .A2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT20), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n446), .A2(new_n451), .A3(new_n448), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n438), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n432), .B1(new_n429), .B2(new_n437), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n307), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G475), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(G234), .A2(G237), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n459), .A2(G952), .A3(new_n260), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n459), .A2(G902), .A3(G953), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(G898), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G116), .B(G122), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT14), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n194), .A2(KEYINPUT14), .A3(G122), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(G107), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT87), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n464), .A2(new_n357), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n228), .A2(G128), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n242), .A2(G143), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n210), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G134), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n470), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT13), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n472), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n471), .A2(new_n478), .ZN(new_n481));
  OAI21_X1  g295(.A(G134), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n464), .A2(new_n357), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n482), .B(new_n473), .C1(new_n483), .C2(new_n470), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT9), .B(G234), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n486), .A2(new_n306), .A3(G953), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n477), .A2(new_n484), .A3(new_n487), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n494), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n458), .A2(new_n463), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n422), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n371), .B(new_n237), .C1(new_n376), .C2(new_n377), .ZN(new_n502));
  INV_X1    g316(.A(new_n224), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n248), .A2(KEYINPUT10), .A3(new_n375), .A4(new_n380), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n245), .B1(new_n247), .B2(new_n236), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n375), .A2(new_n505), .A3(new_n380), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT10), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n502), .A2(new_n503), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT80), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n375), .A2(KEYINPUT10), .A3(new_n380), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n512), .A2(new_n248), .B1(new_n506), .B2(new_n507), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n513), .A2(KEYINPUT80), .A3(new_n503), .A4(new_n502), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n503), .B1(new_n513), .B2(new_n502), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G110), .B(G140), .ZN(new_n519));
  INV_X1    g333(.A(G227), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(G953), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n519), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n511), .B2(new_n514), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n248), .B1(new_n375), .B2(new_n380), .ZN(new_n525));
  INV_X1    g339(.A(new_n506), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n224), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT12), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(KEYINPUT12), .B(new_n224), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n523), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT84), .B(G469), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n307), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT83), .ZN(new_n537));
  INV_X1    g351(.A(new_n522), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n515), .A2(new_n531), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT81), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n515), .A2(KEYINPUT81), .A3(new_n531), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT82), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n515), .B2(new_n538), .ZN(new_n545));
  AOI211_X1 g359(.A(KEYINPUT82), .B(new_n522), .C1(new_n511), .C2(new_n514), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n545), .A2(new_n546), .A3(new_n516), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n537), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n515), .A2(KEYINPUT81), .A3(new_n531), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT81), .B1(new_n515), .B2(new_n531), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n522), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n545), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n516), .B1(new_n524), .B2(new_n544), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n554), .A3(KEYINPUT83), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n548), .A2(new_n307), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n536), .B1(new_n556), .B2(G469), .ZN(new_n557));
  OAI21_X1  g371(.A(G221), .B1(new_n486), .B2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n354), .A2(new_n501), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G101), .ZN(G3));
  OAI21_X1  g376(.A(G472), .B1(new_n295), .B2(G902), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n302), .A2(new_n296), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR4_X1   g379(.A1(new_n557), .A2(new_n565), .A3(new_n353), .A4(new_n559), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT88), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n417), .A2(new_n567), .A3(new_n418), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n401), .A2(new_n413), .A3(KEYINPUT88), .A4(new_n415), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n569), .A2(new_n420), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n491), .B2(G478), .ZN(new_n573));
  OR3_X1    g387(.A1(new_n491), .A2(new_n572), .A3(G478), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n489), .A2(new_n490), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT33), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n492), .A2(G902), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n573), .A2(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n458), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n571), .A2(new_n580), .A3(new_n463), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n566), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT90), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT34), .B(G104), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G6));
  INV_X1    g399(.A(new_n463), .ZN(new_n586));
  AND4_X1   g400(.A1(new_n457), .A2(new_n453), .A3(new_n586), .A4(new_n498), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n587), .A2(new_n568), .A3(new_n570), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n566), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT35), .B(G107), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G9));
  NOR2_X1   g405(.A1(new_n344), .A2(KEYINPUT36), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n339), .B(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n308), .A2(G902), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n350), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(new_n499), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n598), .A2(new_n422), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n557), .A2(new_n565), .A3(new_n559), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT91), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT37), .B(G110), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G12));
  NOR3_X1   g418(.A1(new_n305), .A2(new_n571), .A3(new_n596), .ZN(new_n605));
  INV_X1    g419(.A(new_n497), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(new_n495), .ZN(new_n607));
  INV_X1    g421(.A(G900), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n461), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n460), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n458), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n605), .A2(new_n560), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G128), .ZN(G30));
  XNOR2_X1  g429(.A(new_n611), .B(KEYINPUT39), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n560), .A2(new_n616), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n617), .A2(KEYINPUT40), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(KEYINPUT40), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n298), .A2(new_n304), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n283), .A2(new_n294), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n289), .A2(G472), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(G472), .A2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT93), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n607), .B1(new_n453), .B2(new_n457), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n596), .A2(new_n420), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT92), .B(KEYINPUT38), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n419), .B(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n627), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n618), .A2(new_n619), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G143), .ZN(G45));
  NOR2_X1   g448(.A1(new_n580), .A2(new_n612), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n605), .A2(new_n560), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT94), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n605), .A2(new_n638), .A3(new_n560), .A4(new_n635), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G146), .ZN(G48));
  AOI21_X1  g455(.A(G902), .B1(new_n523), .B2(new_n532), .ZN(new_n642));
  INV_X1    g456(.A(G469), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n535), .B(new_n558), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT95), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n646), .A2(new_n647), .A3(new_n558), .A4(new_n535), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n354), .A2(new_n581), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT41), .B(G113), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G15));
  INV_X1    g466(.A(new_n287), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n620), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n654), .A2(new_n649), .A3(new_n352), .A4(new_n588), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT96), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT96), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n354), .A2(new_n657), .A3(new_n588), .A4(new_n649), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G116), .ZN(G18));
  NOR2_X1   g474(.A1(new_n571), .A2(new_n644), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n654), .A2(new_n598), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G119), .ZN(G21));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n568), .A2(new_n570), .A3(new_n628), .A4(new_n586), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n649), .A2(new_n666), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n300), .A2(new_n301), .B1(new_n268), .B2(new_n284), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT97), .B1(new_n668), .B2(new_n296), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n284), .A2(new_n268), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n291), .B2(new_n292), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT97), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n671), .A2(new_n672), .A3(new_n297), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n352), .B(new_n563), .C1(new_n669), .C2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n664), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n674), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(KEYINPUT98), .A3(new_n649), .A4(new_n666), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G122), .ZN(G24));
  AOI21_X1  g493(.A(new_n187), .B1(new_n302), .B2(new_n307), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n672), .B1(new_n671), .B2(new_n297), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n668), .A2(KEYINPUT97), .A3(new_n296), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n661), .A3(new_n597), .A4(new_n635), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G125), .ZN(G27));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n654), .A2(new_n352), .ZN(new_n687));
  INV_X1    g501(.A(new_n420), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n419), .A2(new_n559), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n515), .A2(new_n544), .A3(new_n538), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n517), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n690), .B1(new_n692), .B2(new_n545), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT100), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n551), .A2(KEYINPUT99), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT99), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n522), .C1(new_n549), .C2(new_n550), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n643), .B1(new_n699), .B2(new_n307), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n689), .B1(new_n700), .B2(new_n536), .ZN(new_n701));
  INV_X1    g515(.A(new_n635), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n687), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n686), .B1(new_n703), .B2(KEYINPUT101), .ZN(new_n704));
  INV_X1    g518(.A(new_n701), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n354), .A3(new_n635), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n707), .A3(KEYINPUT42), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n222), .ZN(G33));
  NAND3_X1  g524(.A1(new_n705), .A2(new_n354), .A3(new_n613), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G134), .ZN(G36));
  NOR2_X1   g526(.A1(new_n458), .A2(new_n578), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT43), .B1(new_n458), .B2(new_n578), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n565), .A2(new_n715), .A3(new_n597), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n718));
  OR3_X1    g532(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT44), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n717), .B2(KEYINPUT44), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n419), .A2(new_n688), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n717), .B2(KEYINPUT44), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n719), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n616), .A2(new_n558), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n548), .A2(new_n728), .A3(new_n555), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n695), .A2(KEYINPUT45), .A3(new_n696), .A4(new_n698), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(G469), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n730), .A3(KEYINPUT102), .A4(G469), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n643), .A2(new_n307), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n736), .A2(new_n739), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n536), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  AOI211_X1 g556(.A(new_n726), .B(new_n727), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n735), .A2(new_n741), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n736), .B1(new_n733), .B2(new_n734), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n744), .B(new_n535), .C1(KEYINPUT46), .C2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n727), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT103), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n725), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  NAND2_X1  g564(.A1(new_n744), .A2(new_n535), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n558), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT47), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n746), .A2(new_n755), .A3(new_n558), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n702), .A2(new_n654), .A3(new_n352), .A4(new_n722), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  AND3_X1   g573(.A1(new_n715), .A2(new_n460), .A3(new_n716), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n676), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n644), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n631), .A2(new_n688), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT50), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n764), .B(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n765), .B2(KEYINPUT50), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n721), .A2(new_n762), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n683), .A2(new_n597), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT110), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n626), .A2(new_n769), .A3(new_n353), .A4(new_n610), .ZN(new_n775));
  INV_X1    g589(.A(new_n458), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n578), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n768), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n761), .A2(new_n722), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT108), .Z(new_n780));
  AND2_X1   g594(.A1(new_n754), .A2(new_n756), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n646), .A2(new_n535), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n558), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n780), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT51), .B1(new_n778), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n771), .A2(new_n687), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT48), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n775), .A2(new_n458), .A3(new_n579), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n676), .A2(new_n760), .A3(new_n661), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(G952), .A3(new_n260), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT112), .Z(new_n793));
  NOR2_X1   g607(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n778), .A2(new_n785), .A3(KEYINPUT51), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(KEYINPUT111), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(KEYINPUT111), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n498), .B(KEYINPUT106), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n580), .B1(new_n800), .B2(new_n458), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n801), .A2(new_n422), .A3(new_n586), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n656), .A2(new_n658), .B1(new_n566), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n675), .A2(new_n677), .B1(new_n599), .B2(new_n600), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n561), .A2(new_n650), .A3(new_n662), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n772), .A2(new_n702), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n721), .A2(new_n776), .A3(new_n611), .A4(new_n800), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n807), .A2(new_n305), .A3(new_n596), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n806), .A2(new_n705), .B1(new_n808), .B2(new_n560), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n704), .A2(new_n708), .A3(new_n711), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n614), .A2(new_n684), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n568), .A2(new_n570), .A3(new_n628), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n815), .A2(new_n597), .A3(new_n559), .A4(new_n612), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n816), .B(new_n626), .C1(new_n536), .C2(new_n700), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n640), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n813), .B1(new_n639), .B2(new_n637), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n817), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n813), .A3(new_n817), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n812), .A2(new_n819), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n812), .A2(new_n819), .A3(KEYINPUT53), .A4(new_n822), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n799), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(KEYINPUT107), .B(KEYINPUT54), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n824), .A2(KEYINPUT53), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n812), .A2(new_n819), .A3(new_n825), .A4(new_n822), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  OAI22_X1  g648(.A1(new_n798), .A2(new_n834), .B1(G952), .B2(G953), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n783), .A2(KEYINPUT49), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT105), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n559), .A2(new_n688), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n713), .A2(new_n352), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n783), .A2(KEYINPUT49), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n627), .A2(new_n631), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n835), .B1(new_n837), .B2(new_n841), .ZN(G75));
  NAND2_X1  g656(.A1(new_n831), .A2(new_n832), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n307), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(G210), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n392), .A2(new_n400), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT113), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT55), .Z(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n398), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n845), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n845), .B2(new_n846), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n260), .A2(G952), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G51));
  NAND2_X1  g668(.A1(new_n843), .A2(new_n829), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n831), .A2(new_n830), .A3(new_n832), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n737), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n533), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n844), .A2(new_n733), .A3(new_n734), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n853), .B1(new_n861), .B2(new_n862), .ZN(G54));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  AND2_X1   g678(.A1(KEYINPUT58), .A2(G475), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n844), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n866), .B2(new_n447), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n853), .B1(new_n866), .B2(new_n447), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n844), .A2(KEYINPUT115), .A3(new_n446), .A4(new_n865), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G60));
  NAND2_X1  g684(.A1(G478), .A2(G902), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT59), .Z(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n828), .B2(new_n833), .ZN(new_n874));
  INV_X1    g688(.A(new_n576), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n853), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n872), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n857), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n831), .A2(new_n830), .A3(new_n832), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n877), .B(new_n878), .C1(new_n880), .C2(new_n833), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n876), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(G63));
  NAND2_X1  g698(.A1(G217), .A2(G902), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n831), .A2(new_n593), .A3(new_n832), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n853), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(KEYINPUT117), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n890), .A2(KEYINPUT61), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n831), .A2(new_n832), .A3(new_n887), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n347), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n888), .A2(new_n889), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n891), .B(new_n895), .ZN(G66));
  OAI21_X1  g710(.A(G953), .B1(new_n462), .B2(new_n395), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT118), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(G953), .ZN(new_n901));
  MUX2_X1   g715(.A(new_n898), .B(KEYINPUT118), .S(new_n901), .Z(new_n902));
  INV_X1    g716(.A(G898), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n848), .B1(new_n903), .B2(G953), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n902), .B(new_n904), .Z(G69));
  XOR2_X1   g719(.A(new_n257), .B(KEYINPUT119), .Z(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(new_n441), .Z(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT120), .Z(new_n908));
  OAI221_X1 g722(.A(G953), .B1(new_n520), .B2(new_n608), .C1(new_n908), .C2(KEYINPUT124), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n907), .B1(G900), .B2(G953), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n687), .A2(new_n815), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n743), .B2(new_n748), .ZN(new_n914));
  INV_X1    g728(.A(new_n811), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n758), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n726), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n746), .A2(KEYINPUT103), .A3(new_n747), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n724), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n820), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n749), .A2(KEYINPUT122), .A3(new_n820), .ZN(new_n924));
  AOI211_X1 g738(.A(KEYINPUT123), .B(new_n916), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n924), .ZN(new_n927));
  INV_X1    g741(.A(new_n916), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n912), .B1(new_n930), .B2(new_n260), .ZN(new_n931));
  INV_X1    g745(.A(new_n908), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n820), .A2(new_n633), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n354), .A2(new_n721), .A3(new_n801), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n933), .A2(KEYINPUT62), .B1(new_n617), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n921), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n758), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n932), .B1(new_n941), .B2(new_n260), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n910), .B1(new_n931), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n260), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n908), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n927), .A2(new_n928), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT123), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n927), .A2(new_n926), .A3(new_n928), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n260), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n911), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n945), .A2(new_n950), .A3(new_n909), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n943), .A2(new_n951), .ZN(G72));
  XNOR2_X1  g766(.A(new_n258), .B(KEYINPUT125), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n937), .A2(new_n940), .A3(new_n899), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n623), .B(KEYINPUT63), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n264), .B(new_n953), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n826), .A2(new_n827), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n265), .A2(new_n289), .A3(new_n280), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n955), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT126), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n853), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n930), .A2(new_n900), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n955), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n953), .A2(new_n264), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G57));
endmodule


