//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0' ..
//Module:
 module locked_locked_c3540( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41,
    G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132,
    G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226,
    G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311,
    G317, G322, G326, G329, G330, G343, G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  , KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64);
input KEYINPUT64;
input KEYINPUT65;
input KEYINPUT66;
input KEYINPUT67;
input KEYINPUT68;
input KEYINPUT69;
input KEYINPUT70;
input KEYINPUT71;
input KEYINPUT72;
input KEYINPUT73;
input KEYINPUT74;
input KEYINPUT75;
input KEYINPUT76;
input KEYINPUT77;
input KEYINPUT78;
input KEYINPUT79;
input KEYINPUT80;
input KEYINPUT81;
input KEYINPUT82;
input KEYINPUT83;
input KEYINPUT84;
input KEYINPUT85;
input KEYINPUT86;
input KEYINPUT87;
input KEYINPUT88;
input KEYINPUT89;
input KEYINPUT90;
input KEYINPUT91;
input KEYINPUT92;
input KEYINPUT93;
input KEYINPUT94;
input KEYINPUT95;
input KEYINPUT96;
input KEYINPUT97;
input KEYINPUT98;
input KEYINPUT99;
input KEYINPUT100;
input KEYINPUT101;
input KEYINPUT102;
input KEYINPUT103;
input KEYINPUT104;
input KEYINPUT105;
input KEYINPUT106;
input KEYINPUT107;
input KEYINPUT108;
input KEYINPUT109;
input KEYINPUT110;
input KEYINPUT111;
input KEYINPUT112;
input KEYINPUT113;
input KEYINPUT114;
input KEYINPUT115;
input KEYINPUT116;
input KEYINPUT117;
input KEYINPUT118;
input KEYINPUT119;
input KEYINPUT120;
input KEYINPUT121;
input KEYINPUT122;
input KEYINPUT123;
input KEYINPUT124;
input KEYINPUT125;
input KEYINPUT126;
input KEYINPUT127;
//Header:
   input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13,
    G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124,
    G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213,
    G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283,
    G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137, new_n138, new_n139, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n172, new_n174, new_n175,
    new_n176, new_n177, new_n178, new_n179, new_n181, new_n182, new_n183,
    new_n184, new_n185, new_n186, new_n187, new_n188, new_n189, new_n190,
    new_n191, new_n192, new_n193, new_n194, new_n195, new_n196, new_n197,
    new_n198, new_n199, new_n200, new_n201, new_n202, new_n203, new_n204,
    new_n205, new_n206, new_n207, new_n208, new_n209, new_n210, new_n211,
    new_n212, new_n213, new_n214, new_n215, new_n216, new_n217, new_n218,
    new_n219, new_n220, new_n221, new_n222, new_n223, new_n224, new_n225,
    new_n226, new_n227, new_n228, new_n229, new_n230, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n262, new_n263, new_n264, new_n265, new_n266, new_n267,
    new_n268, new_n269, new_n270, new_n271, new_n272, new_n273, new_n274,
    new_n275, new_n276, new_n277, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n313, new_n314, new_n315, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n371, new_n372,
    new_n373, new_n374, new_n375, new_n376, new_n377, new_n378, new_n379,
    new_n380, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n400,
    new_n401, new_n402, new_n403, new_n404, new_n405, new_n406, new_n407,
    new_n408, new_n409, new_n410, new_n411, new_n412, new_n413, new_n414,
    new_n415, new_n416, new_n417, new_n418, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n425, new_n426, new_n427, new_n428,
    new_n429, new_n430, new_n431, new_n432, new_n433, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n461, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475, new_n476, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n514,
    new_n515, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041;
wire RLL_wire_A_64;
wire RLL_wire_A_65;
wire RLL_wire_A_66;
wire RLL_wire_A_67;
wire RLL_wire_A_68;
wire RLL_wire_A_69;
wire RLL_wire_A_70;
wire RLL_wire_A_71;
wire RLL_wire_A_72;
wire RLL_wire_A_73;
wire RLL_wire_A_74;
wire RLL_wire_A_75;
wire RLL_wire_A_76;
wire RLL_wire_A_77;
wire RLL_wire_A_78;
wire RLL_wire_A_79;
wire RLL_wire_A_80;
wire RLL_wire_A_81;
wire RLL_wire_A_82;
wire RLL_wire_A_83;
wire RLL_wire_A_84;
wire RLL_wire_A_85;
wire RLL_wire_A_86;
wire RLL_wire_A_87;
wire RLL_wire_A_88;
wire RLL_wire_A_89;
wire RLL_wire_A_90;
wire RLL_wire_A_91;
wire RLL_wire_A_92;
wire RLL_wire_A_93;
wire RLL_wire_A_94;
wire RLL_wire_A_95;
wire RLL_wire_A_96;
wire RLL_wire_A_97;
wire RLL_wire_A_98;
wire RLL_wire_A_99;
wire RLL_wire_A_100;
wire RLL_wire_A_101;
wire RLL_wire_A_102;
wire RLL_wire_A_103;
wire RLL_wire_A_104;
wire RLL_wire_A_105;
wire RLL_wire_A_106;
wire RLL_wire_A_107;
wire RLL_wire_A_108;
wire RLL_wire_A_109;
wire RLL_wire_A_110;
wire RLL_wire_A_111;
wire RLL_wire_A_112;
wire RLL_wire_A_113;
wire RLL_wire_A_114;
wire RLL_wire_A_115;
wire RLL_wire_A_116;
wire RLL_wire_A_117;
wire RLL_wire_A_118;
wire RLL_wire_A_119;
wire RLL_wire_A_120;
wire RLL_wire_A_121;
wire RLL_wire_A_122;
wire RLL_wire_A_123;
wire RLL_wire_A_124;
wire RLL_wire_A_125;
wire RLL_wire_A_126;
wire RLL_wire_A_127;

//Body:
  NOR2_X1   g000(.A1(G58), .A2(G68), .ZN(new_n137));
  INV_X1    g001(.A(G50), .ZN(new_n138));
  NAND2_X1  g002(.A1(new_n137), .A2(new_n138), .ZN(new_n139));
  NOR2_X1   g003(.A1(new_n139), .A2(G77), .ZN(RLL_wire_A_64));
  XNOR2_X1 RLL_XNOR_64 (.A(RLL_wire_A_64), .B(KEYINPUT64), .ZN(G353) );
  OAI21_X1  g004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g005(.A1(G1), .A2(G20), .ZN(new_n142));
  NOR2_X1   g006(.A1(new_n142), .A2(G13), .ZN(new_n143));
  OAI211_X1 g007(.A(new_n143), .B(G250), .C1(G257), .C2(G264), .ZN(new_n144));
  XOR2_X1   g008(.A(new_n144), .B(KEYINPUT0), .Z(new_n145));
  NAND2_X1  g009(.A1(G1), .A2(G13), .ZN(new_n146));
  INV_X1    g010(.A(G20), .ZN(new_n147));
  NOR2_X1   g011(.A1(new_n146), .A2(new_n147), .ZN(RLL_wire_A_65));
  XNOR2_X1 RLL_XNOR_65 (.A(RLL_wire_A_65), .B(KEYINPUT65), .ZN(new_n148) );
  INV_X1    g012(.A(new_n137), .ZN(new_n149));
  NAND2_X1  g013(.A1(new_n149), .A2(G50), .ZN(new_n150));
  INV_X1    g014(.A(new_n150), .ZN(new_n151));
  AOI21_X1  g015(.A(new_n145), .B1(new_n148), .B2(new_n151), .ZN(new_n152));
  AOI22_X1  g016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n153));
  INV_X1    g017(.A(G68), .ZN(new_n154));
  INV_X1    g018(.A(G238), .ZN(new_n155));
  INV_X1    g019(.A(G77), .ZN(new_n156));
  INV_X1    g020(.A(G244), .ZN(new_n157));
  OAI221_X1 g021(.A(new_n153), .B1(new_n154), .B2(new_n155), .C1(new_n156), .C2(new_n157), .ZN(new_n158));
  AOI22_X1  g022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n159));
  AOI22_X1  g023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n160));
  NAND2_X1  g024(.A1(new_n159), .A2(new_n160), .ZN(new_n161));
  OAI21_X1  g025(.A(new_n142), .B1(new_n158), .B2(new_n161), .ZN(new_n162));
  OR2_X1    g026(.A1(new_n162), .A2(KEYINPUT1), .ZN(new_n163));
  NAND2_X1  g027(.A1(new_n162), .A2(KEYINPUT1), .ZN(new_n164));
  AND3_X1   g028(.A1(new_n152), .A2(new_n163), .A3(new_n164), .ZN(G361));
  XOR2_X1   g029(.A(G238), .B(G244), .Z(new_n166));
  XNOR2_X1  g030(.A(new_n166), .B(KEYINPUT2), .ZN(new_n167));
  XOR2_X1   g031(.A(G226), .B(G232), .Z(new_n168));
  XNOR2_X1  g032(.A(new_n167), .B(new_n168), .ZN(new_n169));
  XOR2_X1   g033(.A(G250), .B(G257), .Z(new_n170));
  XNOR2_X1  g034(.A(G264), .B(G270), .ZN(new_n171));
  XNOR2_X1  g035(.A(new_n170), .B(new_n171), .ZN(new_n172));
  XNOR2_X1  g036(.A(new_n169), .B(new_n172), .ZN(G358));
  XOR2_X1   g037(.A(G68), .B(G77), .Z(new_n174));
  XOR2_X1   g038(.A(G50), .B(G58), .Z(new_n175));
  XNOR2_X1  g039(.A(new_n174), .B(new_n175), .ZN(new_n176));
  XOR2_X1   g040(.A(G87), .B(G97), .Z(new_n177));
  XNOR2_X1  g041(.A(G107), .B(G116), .ZN(new_n178));
  XNOR2_X1  g042(.A(new_n177), .B(new_n178), .ZN(new_n179));
  XOR2_X1   g043(.A(new_n176), .B(new_n179), .Z(G351));
  INV_X1    g044(.A(G41), .ZN(new_n181));
  INV_X1    g045(.A(G45), .ZN(new_n182));
  AOI21_X1  g046(.A(G1), .B1(new_n181), .B2(new_n182), .ZN(new_n183));
  NAND2_X1  g047(.A1(G33), .A2(G41), .ZN(new_n184));
  NAND3_X1  g048(.A1(new_n184), .A2(G1), .A3(G13), .ZN(new_n185));
  NAND3_X1  g049(.A1(new_n183), .A2(new_n185), .A3(G274), .ZN(new_n186));
  INV_X1    g050(.A(G226), .ZN(new_n187));
  INV_X1    g051(.A(G1), .ZN(new_n188));
  OAI21_X1  g052(.A(new_n188), .B1(G41), .B2(G45), .ZN(new_n189));
  NAND2_X1  g053(.A1(new_n185), .A2(new_n189), .ZN(new_n190));
  OAI21_X1  g054(.A(new_n186), .B1(new_n187), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G33), .ZN(new_n192));
  INV_X1    g056(.A(G1698), .ZN(new_n193));
  NAND3_X1  g057(.A1(new_n192), .A2(G222), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g058(.A1(new_n192), .A2(G1698), .ZN(new_n195));
  INV_X1    g059(.A(G223), .ZN(new_n196));
  OAI221_X1 g060(.A(new_n194), .B1(new_n156), .B2(new_n192), .C1(new_n195), .C2(new_n196), .ZN(RLL_wire_A_66));
  XOR2_X1 RLL_XOR_66 (.A(RLL_wire_A_66), .B(KEYINPUT66), .Z(new_n197) );
  AOI21_X1  g061(.A(new_n146), .B1(G33), .B2(G41), .ZN(new_n198));
  AOI21_X1  g062(.A(new_n191), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND3_X1  g063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n200));
  NAND2_X1  g064(.A1(new_n200), .A2(new_n146), .ZN(new_n201));
  INV_X1    g065(.A(new_n201), .ZN(new_n202));
  INV_X1    g066(.A(G58), .ZN(new_n203));
  NAND2_X1  g067(.A1(new_n203), .A2(KEYINPUT8), .ZN(new_n204));
  INV_X1    g068(.A(KEYINPUT8), .ZN(new_n205));
  NAND2_X1  g069(.A1(new_n205), .A2(G58), .ZN(new_n206));
  NAND2_X1  g070(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g071(.A1(new_n147), .A2(G33), .ZN(new_n208));
  INV_X1    g072(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g073(.A1(G20), .A2(G33), .ZN(new_n210));
  AOI22_X1  g074(.A1(new_n207), .A2(new_n209), .B1(G150), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g075(.A1(new_n139), .A2(G20), .ZN(new_n212));
  AOI21_X1  g076(.A(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g077(.A1(new_n188), .A2(G13), .A3(G20), .ZN(RLL_wire_A_67));
  XOR2_X1 RLL_XOR_67 (.A(RLL_wire_A_67), .B(KEYINPUT67), .Z(new_n214) );
  NAND2_X1  g078(.A1(new_n202), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g079(.A1(new_n188), .A2(G20), .ZN(new_n216));
  NAND2_X1  g080(.A1(new_n216), .A2(G50), .ZN(new_n217));
  OAI22_X1  g081(.A1(new_n215), .A2(new_n217), .B1(G50), .B2(new_n214), .ZN(new_n218));
  OAI22_X1  g082(.A1(new_n199), .A2(G169), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  INV_X1    g083(.A(G179), .ZN(new_n220));
  AND2_X1   g084(.A1(new_n199), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g085(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g086(.A(new_n186), .B1(new_n157), .B2(new_n190), .ZN(new_n223));
  NAND3_X1  g087(.A1(new_n192), .A2(G232), .A3(new_n193), .ZN(new_n224));
  INV_X1    g088(.A(G107), .ZN(new_n225));
  OAI221_X1 g089(.A(new_n224), .B1(new_n225), .B2(new_n192), .C1(new_n195), .C2(new_n155), .ZN(new_n226));
  AOI21_X1  g090(.A(new_n223), .B1(new_n226), .B2(new_n198), .ZN(RLL_wire_A_68));
  XNOR2_X1 RLL_XNOR_68 (.A(RLL_wire_A_68), .B(KEYINPUT68), .ZN(new_n227) );
  AND2_X1   g091(.A1(new_n227), .A2(G190), .ZN(new_n228));
  XNOR2_X1  g092(.A(KEYINPUT8), .B(G58), .ZN(RLL_wire_A_69));
  XOR2_X1 RLL_XOR_69 (.A(RLL_wire_A_69), .B(KEYINPUT69), .Z(new_n229) );
  INV_X1    g093(.A(new_n210), .ZN(RLL_wire_A_70));
  XNOR2_X1 RLL_XNOR_70 (.A(RLL_wire_A_70), .B(KEYINPUT70), .ZN(new_n230) );
  OAI22_X1  g094(.A1(new_n229), .A2(new_n230), .B1(new_n147), .B2(new_n156), .ZN(new_n231));
  XNOR2_X1  g095(.A(KEYINPUT15), .B(G87), .ZN(new_n232));
  NOR2_X1   g096(.A1(new_n232), .A2(new_n208), .ZN(new_n233));
  OAI21_X1  g097(.A(new_n201), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g098(.A(new_n214), .ZN(new_n235));
  NAND2_X1  g099(.A1(new_n235), .A2(new_n156), .ZN(new_n236));
  NOR2_X1   g100(.A1(new_n235), .A2(new_n201), .ZN(new_n237));
  NAND3_X1  g101(.A1(new_n237), .A2(G77), .A3(new_n216), .ZN(new_n238));
  NAND3_X1  g102(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g103(.A(new_n239), .ZN(new_n240));
  INV_X1    g104(.A(G200), .ZN(RLL_wire_A_71));
  XNOR2_X1 RLL_XNOR_71 (.A(RLL_wire_A_71), .B(KEYINPUT71), .ZN(new_n241) );
  OAI21_X1  g105(.A(new_n240), .B1(new_n227), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g106(.A1(new_n227), .A2(new_n220), .ZN(new_n243));
  OAI21_X1  g107(.A(new_n239), .B1(new_n227), .B2(G169), .ZN(new_n244));
  OAI22_X1  g108(.A1(new_n228), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g109(.A1(new_n213), .A2(new_n218), .ZN(new_n246));
  OR2_X1    g110(.A1(new_n246), .A2(KEYINPUT9), .ZN(RLL_wire_A_72));
  XOR2_X1 RLL_XOR_72 (.A(RLL_wire_A_72), .B(KEYINPUT72), .Z(new_n247) );
  NAND2_X1  g111(.A1(new_n246), .A2(KEYINPUT9), .ZN(new_n248));
  AND2_X1   g112(.A1(new_n247), .A2(new_n248), .ZN(RLL_wire_A_73));
  XOR2_X1 RLL_XOR_73 (.A(RLL_wire_A_73), .B(KEYINPUT73), .Z(new_n249) );
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n250));
  NOR2_X1   g114(.A1(new_n199), .A2(new_n241), .ZN(new_n251));
  INV_X1    g115(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g116(.A1(new_n199), .A2(G190), .ZN(new_n253));
  NAND4_X1  g117(.A1(new_n249), .A2(new_n250), .A3(new_n252), .A4(new_n253), .ZN(new_n254));
  NAND3_X1  g118(.A1(new_n247), .A2(new_n253), .A3(new_n248), .ZN(new_n255));
  OAI21_X1  g119(.A(KEYINPUT10), .B1(new_n255), .B2(new_n251), .ZN(new_n256));
  AOI211_X1 g120(.A(new_n222), .B(new_n245), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g121(.A1(new_n192), .A2(G226), .A3(new_n193), .ZN(new_n258));
  NAND3_X1  g122(.A1(new_n192), .A2(G232), .A3(G1698), .ZN(new_n259));
  NAND2_X1  g123(.A1(G33), .A2(G97), .ZN(new_n260));
  NAND3_X1  g124(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(RLL_wire_A_74));
  XOR2_X1 RLL_XOR_74 (.A(RLL_wire_A_74), .B(KEYINPUT74), .Z(new_n261) );
  NAND2_X1  g125(.A1(new_n261), .A2(new_n198), .ZN(new_n262));
  INV_X1    g126(.A(new_n186), .ZN(new_n263));
  INV_X1    g127(.A(new_n190), .ZN(new_n264));
  AOI21_X1  g128(.A(new_n263), .B1(G238), .B2(new_n264), .ZN(new_n265));
  INV_X1    g129(.A(KEYINPUT13), .ZN(new_n266));
  AND3_X1   g130(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g131(.A(new_n266), .B1(new_n262), .B2(new_n265), .ZN(new_n268));
  OAI21_X1  g132(.A(G200), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g133(.A1(new_n262), .A2(new_n265), .ZN(new_n270));
  NAND2_X1  g134(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n271));
  NAND3_X1  g135(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n272));
  NAND3_X1  g136(.A1(new_n271), .A2(G190), .A3(new_n272), .ZN(new_n273));
  AOI22_X1  g137(.A1(new_n209), .A2(G77), .B1(G20), .B2(new_n154), .ZN(new_n274));
  NAND2_X1  g138(.A1(new_n210), .A2(G50), .ZN(new_n275));
  AOI21_X1  g139(.A(new_n202), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g140(.A(new_n276), .B(KEYINPUT11), .ZN(new_n277));
  NAND3_X1  g141(.A1(new_n237), .A2(G68), .A3(new_n216), .ZN(new_n278));
  NOR3_X1   g142(.A1(new_n214), .A2(KEYINPUT12), .A3(G68), .ZN(new_n279));
  INV_X1    g143(.A(KEYINPUT12), .ZN(new_n280));
  AOI21_X1  g144(.A(new_n280), .B1(new_n235), .B2(new_n154), .ZN(new_n281));
  OAI21_X1  g145(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(RLL_wire_A_75));
  XOR2_X1 RLL_XOR_75 (.A(RLL_wire_A_75), .B(KEYINPUT75), .Z(new_n282) );
  NOR2_X1   g146(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g147(.A1(new_n269), .A2(new_n273), .A3(new_n283), .ZN(new_n284));
  INV_X1    g148(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g149(.A(G169), .B1(new_n267), .B2(new_n268), .ZN(new_n286));
  NAND2_X1  g150(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n287));
  INV_X1    g151(.A(KEYINPUT14), .ZN(new_n288));
  OAI211_X1 g152(.A(new_n288), .B(G169), .C1(new_n267), .C2(new_n268), .ZN(new_n289));
  NAND3_X1  g153(.A1(new_n271), .A2(G179), .A3(new_n272), .ZN(new_n290));
  NAND3_X1  g154(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g155(.A(new_n283), .ZN(new_n292));
  AOI21_X1  g156(.A(new_n285), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g157(.A(G33), .ZN(new_n294));
  NAND2_X1  g158(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n295));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g160(.A1(new_n296), .A2(G33), .ZN(new_n297));
  NAND2_X1  g161(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g162(.A(KEYINPUT7), .B1(new_n298), .B2(new_n147), .ZN(new_n299));
  INV_X1    g163(.A(KEYINPUT7), .ZN(new_n300));
  AOI211_X1 g164(.A(new_n300), .B(G20), .C1(new_n295), .C2(new_n297), .ZN(new_n301));
  OAI21_X1  g165(.A(G68), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g166(.A1(new_n203), .A2(new_n154), .ZN(new_n303));
  OAI21_X1  g167(.A(G20), .B1(new_n303), .B2(new_n137), .ZN(new_n304));
  NAND2_X1  g168(.A1(new_n210), .A2(G159), .ZN(new_n305));
  NAND2_X1  g169(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g170(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g171(.A1(new_n302), .A2(KEYINPUT16), .A3(new_n307), .ZN(new_n308));
  INV_X1    g172(.A(KEYINPUT16), .ZN(new_n309));
  OAI21_X1  g173(.A(new_n300), .B1(new_n192), .B2(G20), .ZN(new_n310));
  NOR2_X1   g174(.A1(new_n296), .A2(G33), .ZN(new_n311));
  NOR2_X1   g175(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n312));
  OAI211_X1 g176(.A(KEYINPUT7), .B(new_n147), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  AOI21_X1  g177(.A(new_n154), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g178(.A(new_n309), .B1(new_n314), .B2(new_n306), .ZN(new_n315));
  NAND3_X1  g179(.A1(new_n308), .A2(new_n315), .A3(new_n201), .ZN(new_n316));
  NAND2_X1  g180(.A1(new_n207), .A2(new_n216), .ZN(new_n317));
  OAI22_X1  g181(.A1(new_n215), .A2(new_n317), .B1(new_n214), .B2(new_n207), .ZN(new_n318));
  INV_X1    g182(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g183(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g184(.A1(new_n295), .A2(new_n297), .A3(G226), .A4(G1698), .ZN(new_n321));
  NAND4_X1  g185(.A1(new_n295), .A2(new_n297), .A3(G223), .A4(new_n193), .ZN(new_n322));
  NAND2_X1  g186(.A1(G33), .A2(G87), .ZN(new_n323));
  NAND3_X1  g187(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g188(.A1(new_n324), .A2(new_n198), .ZN(new_n325));
  NAND3_X1  g189(.A1(new_n185), .A2(G232), .A3(new_n189), .ZN(new_n326));
  NAND2_X1  g190(.A1(new_n186), .A2(new_n326), .ZN(new_n327));
  INV_X1    g191(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g192(.A1(new_n325), .A2(new_n220), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g193(.A(new_n327), .B1(new_n198), .B2(new_n324), .ZN(new_n330));
  OAI21_X1  g194(.A(new_n329), .B1(G169), .B2(new_n330), .ZN(new_n331));
  INV_X1    g195(.A(new_n331), .ZN(new_n332));
  AND3_X1   g196(.A1(new_n320), .A2(new_n332), .A3(KEYINPUT18), .ZN(new_n333));
  AOI21_X1  g197(.A(KEYINPUT18), .B1(new_n320), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g198(.A1(new_n333), .A2(new_n334), .ZN(RLL_wire_A_76));
  XOR2_X1 RLL_XOR_76 (.A(RLL_wire_A_76), .B(KEYINPUT76), .Z(new_n335) );
  INV_X1    g199(.A(G190), .ZN(new_n336));
  NAND3_X1  g200(.A1(new_n325), .A2(new_n336), .A3(new_n328), .ZN(new_n337));
  OAI21_X1  g201(.A(new_n337), .B1(G200), .B2(new_n330), .ZN(new_n338));
  NAND3_X1  g202(.A1(new_n316), .A2(new_n319), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g203(.A1(new_n339), .A2(KEYINPUT17), .ZN(new_n340));
  INV_X1    g204(.A(KEYINPUT17), .ZN(RLL_wire_A_77));
  XNOR2_X1 RLL_XNOR_77 (.A(RLL_wire_A_77), .B(KEYINPUT77), .ZN(new_n341) );
  NAND4_X1  g205(.A1(new_n316), .A2(new_n338), .A3(new_n341), .A4(new_n319), .ZN(RLL_wire_A_78));
  XNOR2_X1 RLL_XNOR_78 (.A(RLL_wire_A_78), .B(KEYINPUT78), .ZN(new_n342) );
  AND2_X1   g206(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g207(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  AND3_X1   g208(.A1(new_n257), .A2(new_n293), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g209(.A1(new_n210), .A2(G77), .ZN(new_n346));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n347));
  INV_X1    g211(.A(G97), .ZN(new_n348));
  NOR3_X1   g212(.A1(new_n347), .A2(new_n348), .A3(G107), .ZN(new_n349));
  XNOR2_X1  g213(.A(G97), .B(G107), .ZN(new_n350));
  AOI21_X1  g214(.A(new_n349), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g215(.A(new_n346), .B1(new_n351), .B2(new_n147), .ZN(new_n352));
  AOI21_X1  g216(.A(new_n225), .B1(new_n310), .B2(new_n313), .ZN(new_n353));
  OAI21_X1  g217(.A(new_n201), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g218(.A1(new_n214), .A2(G97), .ZN(new_n355));
  NAND2_X1  g219(.A1(new_n188), .A2(G33), .ZN(RLL_wire_A_79));
  XOR2_X1 RLL_XOR_79 (.A(RLL_wire_A_79), .B(KEYINPUT79), .Z(new_n356) );
  AND3_X1   g220(.A1(new_n202), .A2(new_n214), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g221(.A(new_n355), .B1(new_n357), .B2(G97), .ZN(new_n358));
  AND2_X1   g222(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g223(.A1(new_n295), .A2(new_n297), .A3(G244), .A4(new_n193), .ZN(new_n360));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n361));
  NAND2_X1  g225(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g226(.A1(new_n192), .A2(KEYINPUT4), .A3(G244), .A4(new_n193), .ZN(new_n363));
  NAND2_X1  g227(.A1(G33), .A2(G283), .ZN(new_n364));
  NAND3_X1  g228(.A1(new_n192), .A2(G250), .A3(G1698), .ZN(new_n365));
  NAND4_X1  g229(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g230(.A1(new_n366), .A2(new_n198), .ZN(RLL_wire_A_80));
  XOR2_X1 RLL_XOR_80 (.A(RLL_wire_A_80), .B(KEYINPUT80), .Z(new_n367) );
  OAI211_X1 g231(.A(new_n188), .B(G45), .C1(new_n181), .C2(KEYINPUT5), .ZN(new_n368));
  INV_X1    g232(.A(new_n368), .ZN(new_n369));
  INV_X1    g233(.A(KEYINPUT5), .ZN(new_n370));
  NOR2_X1   g234(.A1(new_n370), .A2(G41), .ZN(new_n371));
  INV_X1    g235(.A(new_n371), .ZN(new_n372));
  NAND4_X1  g236(.A1(new_n369), .A2(G274), .A3(new_n185), .A4(new_n372), .ZN(new_n373));
  OAI211_X1 g237(.A(G257), .B(new_n185), .C1(new_n368), .C2(new_n371), .ZN(new_n374));
  NAND2_X1  g238(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g239(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g240(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g241(.A1(new_n377), .A2(G200), .ZN(new_n378));
  AOI21_X1  g242(.A(new_n375), .B1(new_n366), .B2(new_n198), .ZN(new_n379));
  NAND2_X1  g243(.A1(new_n379), .A2(G190), .ZN(new_n380));
  NAND3_X1  g244(.A1(new_n359), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g245(.A1(new_n354), .A2(new_n358), .ZN(new_n382));
  NAND3_X1  g246(.A1(new_n367), .A2(new_n220), .A3(new_n376), .ZN(new_n383));
  OAI211_X1 g247(.A(new_n382), .B(new_n383), .C1(G169), .C2(new_n379), .ZN(new_n384));
  NAND2_X1  g248(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g249(.A1(new_n185), .A2(new_n188), .A3(G45), .A4(G274), .ZN(new_n386));
  NAND2_X1  g250(.A1(new_n188), .A2(G45), .ZN(new_n387));
  NAND3_X1  g251(.A1(new_n185), .A2(G250), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g252(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g253(.A1(new_n295), .A2(new_n297), .A3(G238), .A4(new_n193), .ZN(new_n390));
  NAND4_X1  g254(.A1(new_n295), .A2(new_n297), .A3(G244), .A4(G1698), .ZN(new_n391));
  INV_X1    g255(.A(G116), .ZN(new_n392));
  OAI211_X1 g256(.A(new_n390), .B(new_n391), .C1(new_n294), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g257(.A(new_n389), .B1(new_n393), .B2(new_n198), .ZN(new_n394));
  NAND2_X1  g258(.A1(new_n394), .A2(new_n220), .ZN(new_n395));
  OAI21_X1  g259(.A(new_n395), .B1(G169), .B2(new_n394), .ZN(new_n396));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n397));
  OAI21_X1  g261(.A(new_n147), .B1(new_n260), .B2(new_n397), .ZN(new_n398));
  INV_X1    g262(.A(G87), .ZN(new_n399));
  NAND3_X1  g263(.A1(new_n399), .A2(new_n348), .A3(new_n225), .ZN(new_n400));
  NAND2_X1  g264(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g265(.A1(new_n295), .A2(new_n297), .A3(new_n147), .A4(G68), .ZN(new_n402));
  OAI21_X1  g266(.A(new_n397), .B1(new_n208), .B2(new_n348), .ZN(new_n403));
  NAND3_X1  g267(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI22_X1  g268(.A1(new_n404), .A2(new_n201), .B1(new_n235), .B2(new_n232), .ZN(new_n405));
  INV_X1    g269(.A(new_n232), .ZN(new_n406));
  NAND2_X1  g270(.A1(new_n357), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g271(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g272(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g273(.A1(new_n357), .A2(G87), .ZN(new_n410));
  OAI211_X1 g274(.A(new_n405), .B(new_n410), .C1(new_n394), .C2(new_n241), .ZN(new_n411));
  NAND2_X1  g275(.A1(new_n394), .A2(G190), .ZN(new_n412));
  INV_X1    g276(.A(new_n412), .ZN(new_n413));
  OAI22_X1  g277(.A1(new_n396), .A2(new_n409), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g278(.A1(new_n385), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g279(.A(G270), .B(new_n185), .C1(new_n368), .C2(new_n371), .ZN(new_n416));
  AND2_X1   g280(.A1(new_n373), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g281(.A1(new_n295), .A2(new_n297), .A3(G257), .A4(new_n193), .ZN(new_n418));
  NAND4_X1  g282(.A1(new_n295), .A2(new_n297), .A3(G264), .A4(G1698), .ZN(new_n419));
  INV_X1    g283(.A(G303), .ZN(new_n420));
  OAI211_X1 g284(.A(new_n418), .B(new_n419), .C1(new_n420), .C2(new_n192), .ZN(new_n421));
  NAND2_X1  g285(.A1(new_n421), .A2(new_n198), .ZN(new_n422));
  NAND2_X1  g286(.A1(new_n417), .A2(new_n422), .ZN(RLL_wire_A_81));
  XNOR2_X1 RLL_XNOR_81 (.A(RLL_wire_A_81), .B(KEYINPUT81), .ZN(new_n423) );
  NAND3_X1  g287(.A1(new_n237), .A2(G116), .A3(new_n356), .ZN(new_n424));
  NAND2_X1  g288(.A1(new_n235), .A2(new_n392), .ZN(new_n425));
  AOI22_X1  g289(.A1(new_n200), .A2(new_n146), .B1(G20), .B2(new_n392), .ZN(new_n426));
  OAI211_X1 g290(.A(new_n364), .B(new_n147), .C1(G33), .C2(new_n348), .ZN(new_n427));
  AND3_X1   g291(.A1(new_n426), .A2(KEYINPUT20), .A3(new_n427), .ZN(RLL_wire_A_82));
  XOR2_X1 RLL_XOR_82 (.A(RLL_wire_A_82), .B(KEYINPUT82), .Z(new_n428) );
  AOI21_X1  g292(.A(KEYINPUT20), .B1(new_n426), .B2(new_n427), .ZN(new_n429));
  OAI211_X1 g293(.A(new_n424), .B(new_n425), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND4_X1  g294(.A1(new_n423), .A2(KEYINPUT21), .A3(G169), .A4(new_n430), .ZN(new_n431));
  NAND4_X1  g295(.A1(new_n430), .A2(G179), .A3(new_n422), .A4(new_n417), .ZN(new_n432));
  AND2_X1   g296(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g297(.A1(new_n423), .A2(G169), .A3(new_n430), .ZN(new_n434));
  INV_X1    g298(.A(KEYINPUT21), .ZN(new_n435));
  NAND2_X1  g299(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g300(.A(new_n430), .B1(new_n423), .B2(G200), .ZN(new_n437));
  OAI21_X1  g301(.A(new_n437), .B1(new_n336), .B2(new_n423), .ZN(new_n438));
  AND3_X1   g302(.A1(new_n433), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g303(.A1(new_n295), .A2(new_n297), .A3(new_n147), .A4(G87), .ZN(new_n440));
  NAND2_X1  g304(.A1(new_n440), .A2(KEYINPUT22), .ZN(RLL_wire_A_83));
  XNOR2_X1 RLL_XNOR_83 (.A(RLL_wire_A_83), .B(KEYINPUT83), .ZN(new_n441) );
  INV_X1    g305(.A(KEYINPUT22), .ZN(new_n442));
  NAND4_X1  g306(.A1(new_n192), .A2(new_n442), .A3(new_n147), .A4(G87), .ZN(new_n443));
  NAND2_X1  g307(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g308(.A(KEYINPUT24), .ZN(new_n445));
  NOR3_X1   g309(.A1(new_n294), .A2(new_n392), .A3(G20), .ZN(new_n446));
  INV_X1    g310(.A(KEYINPUT23), .ZN(new_n447));
  AOI21_X1  g311(.A(new_n447), .B1(G20), .B2(new_n225), .ZN(new_n448));
  NOR3_X1   g312(.A1(new_n147), .A2(KEYINPUT23), .A3(G107), .ZN(new_n449));
  NOR3_X1   g313(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND3_X1   g314(.A1(new_n444), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g315(.A(new_n445), .B1(new_n444), .B2(new_n450), .ZN(RLL_wire_A_84));
  XNOR2_X1 RLL_XNOR_84 (.A(RLL_wire_A_84), .B(KEYINPUT84), .ZN(new_n452) );
  OAI21_X1  g316(.A(new_n201), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g317(.A(KEYINPUT25), .ZN(new_n454));
  NOR3_X1   g318(.A1(new_n214), .A2(new_n454), .A3(G107), .ZN(RLL_wire_A_85));
  XNOR2_X1 RLL_XNOR_85 (.A(RLL_wire_A_85), .B(KEYINPUT85), .ZN(new_n455) );
  INV_X1    g319(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g320(.A(new_n454), .B1(new_n214), .B2(G107), .ZN(new_n457));
  AOI22_X1  g321(.A1(new_n357), .A2(G107), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g322(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g323(.A1(new_n295), .A2(new_n297), .A3(G257), .A4(G1698), .ZN(new_n460));
  NAND4_X1  g324(.A1(new_n295), .A2(new_n297), .A3(G250), .A4(new_n193), .ZN(RLL_wire_A_86));
  XOR2_X1 RLL_XOR_86 (.A(RLL_wire_A_86), .B(KEYINPUT86), .Z(new_n461) );
  INV_X1    g325(.A(G294), .ZN(new_n462));
  OAI211_X1 g326(.A(new_n460), .B(new_n461), .C1(new_n294), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g327(.A1(new_n463), .A2(new_n198), .ZN(new_n464));
  OAI211_X1 g328(.A(G264), .B(new_n185), .C1(new_n368), .C2(new_n371), .ZN(new_n465));
  NAND3_X1  g329(.A1(new_n464), .A2(new_n373), .A3(new_n465), .ZN(RLL_wire_A_87));
  XOR2_X1 RLL_XOR_87 (.A(RLL_wire_A_87), .B(KEYINPUT87), .Z(new_n466) );
  NAND2_X1  g330(.A1(new_n466), .A2(G169), .ZN(new_n467));
  INV_X1    g331(.A(new_n465), .ZN(new_n468));
  AOI21_X1  g332(.A(new_n468), .B1(new_n463), .B2(new_n198), .ZN(RLL_wire_A_88));
  XOR2_X1 RLL_XOR_88 (.A(RLL_wire_A_88), .B(KEYINPUT88), .Z(new_n469) );
  NAND3_X1  g333(.A1(new_n469), .A2(G179), .A3(new_n373), .ZN(new_n470));
  NAND2_X1  g334(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g335(.A1(new_n459), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g336(.A1(new_n466), .A2(G190), .ZN(new_n473));
  AOI21_X1  g337(.A(G200), .B1(new_n469), .B2(new_n373), .ZN(new_n474));
  OAI211_X1 g338(.A(new_n453), .B(new_n458), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  AND2_X1   g339(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AND4_X1   g340(.A1(new_n345), .A2(new_n415), .A3(new_n439), .A4(new_n476), .ZN(G372));
  NAND2_X1  g341(.A1(new_n393), .A2(new_n198), .ZN(new_n478));
  INV_X1    g342(.A(new_n389), .ZN(new_n479));
  AOI21_X1  g343(.A(G169), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g344(.A(new_n480), .B1(new_n220), .B2(new_n394), .ZN(new_n481));
  AOI21_X1  g345(.A(new_n241), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  NAND2_X1  g346(.A1(new_n405), .A2(new_n410), .ZN(new_n483));
  NOR2_X1   g347(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g348(.A1(new_n481), .A2(new_n408), .B1(new_n484), .B2(new_n412), .ZN(new_n485));
  NAND4_X1  g349(.A1(new_n485), .A2(new_n384), .A3(new_n381), .A4(new_n475), .ZN(new_n486));
  NAND3_X1  g350(.A1(new_n436), .A2(new_n432), .A3(new_n431), .ZN(new_n487));
  AOI22_X1  g351(.A1(new_n453), .A2(new_n458), .B1(new_n467), .B2(new_n470), .ZN(new_n488));
  NOR2_X1   g352(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g353(.A1(new_n486), .A2(new_n489), .ZN(RLL_wire_A_89));
  XOR2_X1 RLL_XOR_89 (.A(RLL_wire_A_89), .B(KEYINPUT89), .Z(new_n490) );
  NAND2_X1  g354(.A1(new_n481), .A2(new_n408), .ZN(new_n491));
  OAI21_X1  g355(.A(new_n383), .B1(G169), .B2(new_n379), .ZN(new_n492));
  NOR2_X1   g356(.A1(new_n492), .A2(new_n359), .ZN(new_n493));
  AOI21_X1  g357(.A(KEYINPUT26), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  INV_X1    g358(.A(KEYINPUT26), .ZN(new_n495));
  NOR3_X1   g359(.A1(new_n414), .A2(new_n384), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g360(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g361(.A(new_n345), .B1(new_n490), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g362(.A(new_n331), .B1(new_n316), .B2(new_n319), .ZN(new_n499));
  XNOR2_X1  g363(.A(new_n499), .B(KEYINPUT18), .ZN(new_n500));
  NOR2_X1   g364(.A1(new_n243), .A2(new_n244), .ZN(new_n501));
  AOI22_X1  g365(.A1(new_n291), .A2(new_n292), .B1(new_n284), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g366(.A(new_n500), .B1(new_n502), .B2(new_n343), .ZN(new_n503));
  NAND2_X1  g367(.A1(new_n254), .A2(new_n256), .ZN(new_n504));
  AOI21_X1  g368(.A(new_n222), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g369(.A1(new_n498), .A2(new_n505), .ZN(G369));
  NAND3_X1  g370(.A1(new_n188), .A2(new_n147), .A3(G13), .ZN(new_n507));
  OR2_X1    g371(.A1(new_n507), .A2(KEYINPUT27), .ZN(RLL_wire_A_90));
  XOR2_X1 RLL_XOR_90 (.A(RLL_wire_A_90), .B(KEYINPUT90), .Z(new_n508) );
  NAND2_X1  g372(.A1(new_n507), .A2(KEYINPUT27), .ZN(RLL_wire_A_91));
  XOR2_X1 RLL_XOR_91 (.A(RLL_wire_A_91), .B(KEYINPUT91), .Z(new_n509) );
  NAND3_X1  g373(.A1(new_n508), .A2(G213), .A3(new_n509), .ZN(new_n510));
  INV_X1    g374(.A(G343), .ZN(new_n511));
  NOR2_X1   g375(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g376(.A1(new_n430), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g377(.A1(new_n487), .A2(new_n513), .ZN(new_n514));
  INV_X1    g378(.A(new_n439), .ZN(new_n515));
  OAI21_X1  g379(.A(new_n514), .B1(new_n515), .B2(new_n513), .ZN(new_n516));
  INV_X1    g380(.A(new_n516), .ZN(new_n517));
  INV_X1    g381(.A(G330), .ZN(new_n518));
  NOR2_X1   g382(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g383(.A1(new_n459), .A2(new_n512), .ZN(new_n520));
  NAND2_X1  g384(.A1(new_n476), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g385(.A1(new_n459), .A2(new_n471), .A3(new_n512), .ZN(new_n522));
  NAND2_X1  g386(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g387(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g388(.A(new_n512), .B1(new_n433), .B2(new_n436), .ZN(new_n525));
  INV_X1    g389(.A(new_n512), .ZN(new_n526));
  AOI22_X1  g390(.A1(new_n523), .A2(new_n525), .B1(new_n488), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g391(.A1(new_n524), .A2(new_n527), .ZN(G399));
  NOR2_X1   g392(.A1(new_n400), .A2(G116), .ZN(new_n529));
  NAND2_X1  g393(.A1(new_n143), .A2(new_n181), .ZN(RLL_wire_A_92));
  XNOR2_X1 RLL_XNOR_92 (.A(RLL_wire_A_92), .B(KEYINPUT92), .ZN(new_n530) );
  NAND3_X1  g394(.A1(new_n529), .A2(new_n530), .A3(G1), .ZN(new_n531));
  OAI21_X1  g395(.A(new_n531), .B1(new_n150), .B2(new_n530), .ZN(new_n532));
  XNOR2_X1  g396(.A(new_n532), .B(KEYINPUT28), .ZN(new_n533));
  INV_X1    g397(.A(KEYINPUT31), .ZN(RLL_wire_A_93));
  XOR2_X1 RLL_XOR_93 (.A(RLL_wire_A_93), .B(KEYINPUT93), .Z(new_n534) );
  AND2_X1   g398(.A1(new_n469), .A2(new_n394), .ZN(RLL_wire_A_94));
  XOR2_X1 RLL_XOR_94 (.A(RLL_wire_A_94), .B(KEYINPUT94), .Z(new_n535) );
  AND3_X1   g399(.A1(new_n417), .A2(G179), .A3(new_n422), .ZN(new_n536));
  NAND3_X1  g400(.A1(new_n535), .A2(new_n536), .A3(new_n379), .ZN(new_n537));
  INV_X1    g401(.A(KEYINPUT30), .ZN(RLL_wire_A_95));
  XOR2_X1 RLL_XOR_95 (.A(RLL_wire_A_95), .B(KEYINPUT95), .Z(new_n538) );
  NAND2_X1  g402(.A1(new_n478), .A2(new_n479), .ZN(new_n539));
  AND3_X1   g403(.A1(new_n423), .A2(new_n220), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g404(.A1(new_n367), .A2(new_n376), .B1(new_n469), .B2(new_n373), .ZN(new_n541));
  AOI22_X1  g405(.A1(new_n537), .A2(new_n538), .B1(new_n540), .B2(new_n541), .ZN(RLL_wire_A_96));
  XNOR2_X1 RLL_XNOR_96 (.A(RLL_wire_A_96), .B(KEYINPUT96), .ZN(new_n542) );
  NAND4_X1  g406(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT30), .A4(new_n379), .ZN(new_n543));
  AOI211_X1 g407(.A(new_n534), .B(new_n526), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g408(.A1(new_n537), .A2(new_n538), .ZN(new_n545));
  NAND2_X1  g409(.A1(new_n540), .A2(new_n541), .ZN(new_n546));
  NAND3_X1  g410(.A1(new_n545), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g411(.A(KEYINPUT31), .B1(new_n547), .B2(new_n512), .ZN(new_n548));
  NOR2_X1   g412(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g413(.A1(new_n415), .A2(new_n439), .A3(new_n476), .A4(new_n526), .ZN(new_n550));
  AOI21_X1  g414(.A(new_n518), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g415(.A(new_n526), .B1(new_n497), .B2(new_n490), .ZN(new_n552));
  INV_X1    g416(.A(KEYINPUT29), .ZN(new_n553));
  NAND2_X1  g417(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g418(.A(new_n491), .ZN(new_n555));
  NAND3_X1  g419(.A1(new_n485), .A2(new_n493), .A3(KEYINPUT26), .ZN(new_n556));
  OAI21_X1  g420(.A(new_n495), .B1(new_n414), .B2(new_n384), .ZN(RLL_wire_A_97));
  XOR2_X1 RLL_XOR_97 (.A(RLL_wire_A_97), .B(KEYINPUT97), .Z(new_n557) );
  AOI21_X1  g421(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g422(.A1(new_n472), .A2(new_n433), .A3(new_n436), .ZN(new_n559));
  AND2_X1   g423(.A1(new_n381), .A2(new_n384), .ZN(new_n560));
  NAND4_X1  g424(.A1(new_n559), .A2(new_n560), .A3(new_n485), .A4(new_n475), .ZN(RLL_wire_A_98));
  XOR2_X1 RLL_XOR_98 (.A(RLL_wire_A_98), .B(KEYINPUT98), .Z(new_n561) );
  AOI21_X1  g425(.A(new_n512), .B1(new_n558), .B2(new_n561), .ZN(RLL_wire_A_99));
  XNOR2_X1 RLL_XNOR_99 (.A(RLL_wire_A_99), .B(KEYINPUT99), .ZN(new_n562) );
  NAND2_X1  g426(.A1(new_n562), .A2(KEYINPUT29), .ZN(new_n563));
  AOI21_X1  g427(.A(new_n551), .B1(new_n554), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g428(.A(new_n533), .B1(new_n564), .B2(G1), .ZN(G364));
  NAND2_X1  g429(.A1(new_n517), .A2(new_n518), .ZN(new_n566));
  INV_X1    g430(.A(new_n519), .ZN(new_n567));
  AND2_X1   g431(.A1(new_n147), .A2(G13), .ZN(new_n568));
  NAND2_X1  g432(.A1(new_n568), .A2(G45), .ZN(new_n569));
  NAND3_X1  g433(.A1(new_n530), .A2(new_n569), .A3(G1), .ZN(new_n570));
  NAND3_X1  g434(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  INV_X1    g435(.A(new_n570), .ZN(new_n572));
  NAND2_X1  g436(.A1(new_n192), .A2(new_n143), .ZN(new_n573));
  INV_X1    g437(.A(G355), .ZN(new_n574));
  OAI22_X1  g438(.A1(new_n573), .A2(new_n574), .B1(G116), .B2(new_n143), .ZN(new_n575));
  NAND2_X1  g439(.A1(new_n176), .A2(G45), .ZN(new_n576));
  NAND2_X1  g440(.A1(new_n298), .A2(new_n143), .ZN(new_n577));
  AOI21_X1  g441(.A(new_n577), .B1(new_n182), .B2(new_n151), .ZN(new_n578));
  AOI21_X1  g442(.A(new_n575), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g443(.A1(G13), .A2(G33), .ZN(new_n580));
  INV_X1    g444(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g445(.A1(new_n581), .A2(G20), .ZN(new_n582));
  INV_X1    g446(.A(G169), .ZN(new_n583));
  AOI21_X1  g447(.A(new_n146), .B1(G20), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g448(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g449(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g450(.A(new_n572), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g451(.A1(new_n147), .A2(new_n220), .ZN(new_n588));
  INV_X1    g452(.A(new_n588), .ZN(new_n589));
  NOR3_X1   g453(.A1(new_n589), .A2(new_n336), .A3(G200), .ZN(new_n590));
  INV_X1    g454(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g455(.A1(new_n589), .A2(G190), .A3(G200), .ZN(new_n592));
  INV_X1    g456(.A(new_n592), .ZN(new_n593));
  OAI22_X1  g457(.A1(new_n203), .A2(new_n591), .B1(new_n593), .B2(new_n156), .ZN(RLL_wire_A_100));
  XOR2_X1 RLL_XOR_100 (.A(RLL_wire_A_100), .B(KEYINPUT100), .Z(new_n594) );
  NAND2_X1  g458(.A1(new_n588), .A2(G200), .ZN(RLL_wire_A_101));
  XOR2_X1 RLL_XOR_101 (.A(RLL_wire_A_101), .B(KEYINPUT101), .Z(new_n595) );
  NOR2_X1   g459(.A1(new_n595), .A2(new_n336), .ZN(new_n596));
  AOI21_X1  g460(.A(new_n594), .B1(G50), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g461(.A1(new_n147), .A2(G190), .ZN(new_n598));
  NOR2_X1   g462(.A1(G179), .A2(G200), .ZN(new_n599));
  NAND2_X1  g463(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g464(.A(G159), .ZN(new_n601));
  NOR2_X1   g465(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g466(.A(new_n602), .B(KEYINPUT32), .ZN(new_n603));
  NOR2_X1   g467(.A1(new_n241), .A2(G179), .ZN(new_n604));
  NAND3_X1  g468(.A1(new_n604), .A2(G20), .A3(G190), .ZN(new_n605));
  OAI21_X1  g469(.A(new_n192), .B1(new_n605), .B2(new_n399), .ZN(new_n606));
  NAND2_X1  g470(.A1(new_n604), .A2(new_n598), .ZN(new_n607));
  INV_X1    g471(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g472(.A(new_n606), .B1(G107), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g473(.A1(new_n595), .A2(G190), .ZN(new_n610));
  AOI21_X1  g474(.A(new_n147), .B1(new_n599), .B2(G190), .ZN(new_n611));
  INV_X1    g475(.A(new_n611), .ZN(new_n612));
  AOI22_X1  g476(.A1(new_n610), .A2(G68), .B1(G97), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g477(.A1(new_n597), .A2(new_n603), .A3(new_n609), .A4(new_n613), .ZN(new_n614));
  INV_X1    g478(.A(new_n596), .ZN(new_n615));
  INV_X1    g479(.A(G326), .ZN(new_n616));
  OAI22_X1  g480(.A1(new_n615), .A2(new_n616), .B1(new_n611), .B2(new_n462), .ZN(new_n617));
  AOI21_X1  g481(.A(new_n617), .B1(G311), .B2(new_n592), .ZN(new_n618));
  INV_X1    g482(.A(new_n605), .ZN(new_n619));
  AOI21_X1  g483(.A(new_n192), .B1(new_n619), .B2(G303), .ZN(new_n620));
  INV_X1    g484(.A(new_n600), .ZN(new_n621));
  AOI22_X1  g485(.A1(new_n608), .A2(G283), .B1(new_n621), .B2(G329), .ZN(new_n622));
  XNOR2_X1  g486(.A(KEYINPUT33), .B(G317), .ZN(new_n623));
  AOI22_X1  g487(.A1(G322), .A2(new_n590), .B1(new_n610), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g488(.A1(new_n618), .A2(new_n620), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g489(.A1(new_n614), .A2(new_n625), .ZN(RLL_wire_A_102));
  XNOR2_X1 RLL_XNOR_102 (.A(RLL_wire_A_102), .B(KEYINPUT102), .ZN(new_n626) );
  AOI21_X1  g490(.A(new_n587), .B1(new_n626), .B2(new_n584), .ZN(new_n627));
  INV_X1    g491(.A(new_n582), .ZN(RLL_wire_A_103));
  XOR2_X1 RLL_XOR_103 (.A(RLL_wire_A_103), .B(KEYINPUT103), .Z(new_n628) );
  OAI21_X1  g492(.A(new_n627), .B1(new_n516), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g493(.A1(new_n571), .A2(new_n629), .ZN(new_n630));
  INV_X1    g494(.A(new_n630), .ZN(G396));
  NOR2_X1   g495(.A1(new_n584), .A2(new_n580), .ZN(new_n632));
  INV_X1    g496(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g497(.A(new_n572), .B1(G77), .B2(new_n633), .ZN(new_n634));
  INV_X1    g498(.A(new_n610), .ZN(new_n635));
  INV_X1    g499(.A(G283), .ZN(new_n636));
  OAI22_X1  g500(.A1(new_n593), .A2(new_n392), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g501(.A(new_n637), .B1(G303), .B2(new_n596), .ZN(new_n638));
  AOI21_X1  g502(.A(new_n192), .B1(new_n619), .B2(G107), .ZN(new_n639));
  AOI22_X1  g503(.A1(new_n608), .A2(G87), .B1(new_n621), .B2(G311), .ZN(new_n640));
  AOI22_X1  g504(.A1(new_n590), .A2(G294), .B1(G97), .B2(new_n612), .ZN(new_n641));
  NAND4_X1  g505(.A1(new_n638), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  AOI22_X1  g506(.A1(G137), .A2(new_n596), .B1(new_n610), .B2(G150), .ZN(new_n643));
  INV_X1    g507(.A(G143), .ZN(new_n644));
  OAI221_X1 g508(.A(new_n643), .B1(new_n644), .B2(new_n591), .C1(new_n601), .C2(new_n593), .ZN(new_n645));
  XOR2_X1   g509(.A(new_n645), .B(KEYINPUT34), .Z(new_n646));
  AOI22_X1  g510(.A1(new_n619), .A2(G50), .B1(new_n608), .B2(G68), .ZN(new_n647));
  AOI21_X1  g511(.A(new_n298), .B1(new_n621), .B2(G132), .ZN(new_n648));
  OAI211_X1 g512(.A(new_n647), .B(new_n648), .C1(new_n203), .C2(new_n611), .ZN(new_n649));
  OAI21_X1  g513(.A(new_n642), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g514(.A(new_n634), .B1(new_n650), .B2(new_n584), .ZN(new_n651));
  OR2_X1    g515(.A1(new_n243), .A2(new_n244), .ZN(new_n652));
  NAND2_X1  g516(.A1(new_n239), .A2(new_n512), .ZN(RLL_wire_A_104));
  XOR2_X1 RLL_XOR_104 (.A(RLL_wire_A_104), .B(KEYINPUT104), .Z(new_n653) );
  OAI211_X1 g517(.A(new_n652), .B(new_n653), .C1(new_n228), .C2(new_n242), .ZN(new_n654));
  NAND3_X1  g518(.A1(new_n501), .A2(new_n239), .A3(new_n512), .ZN(new_n655));
  NAND2_X1  g519(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g520(.A(new_n651), .B1(new_n581), .B2(new_n656), .ZN(new_n657));
  INV_X1    g521(.A(new_n656), .ZN(new_n658));
  NAND2_X1  g522(.A1(new_n552), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g523(.A(new_n526), .B(new_n656), .C1(new_n497), .C2(new_n490), .ZN(new_n660));
  NAND3_X1  g524(.A1(new_n659), .A2(new_n551), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g525(.A1(new_n661), .A2(new_n570), .ZN(new_n662));
  AOI21_X1  g526(.A(new_n551), .B1(new_n659), .B2(new_n660), .ZN(new_n663));
  OAI21_X1  g527(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(G384));
  INV_X1    g528(.A(new_n351), .ZN(new_n665));
  OAI211_X1 g529(.A(G116), .B(new_n148), .C1(new_n665), .C2(KEYINPUT35), .ZN(new_n666));
  AOI21_X1  g530(.A(new_n666), .B1(KEYINPUT35), .B2(new_n665), .ZN(new_n667));
  XNOR2_X1  g531(.A(new_n667), .B(KEYINPUT36), .ZN(new_n668));
  OR3_X1    g532(.A1(new_n150), .A2(new_n156), .A3(new_n303), .ZN(new_n669));
  NAND2_X1  g533(.A1(new_n138), .A2(G68), .ZN(new_n670));
  AOI211_X1 g534(.A(new_n188), .B(G13), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  NOR2_X1   g535(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g536(.A1(new_n652), .A2(new_n512), .ZN(new_n673));
  INV_X1    g537(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g538(.A1(new_n660), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g539(.A1(new_n291), .A2(new_n292), .ZN(new_n676));
  NAND2_X1  g540(.A1(new_n292), .A2(new_n512), .ZN(new_n677));
  NAND3_X1  g541(.A1(new_n676), .A2(new_n284), .A3(new_n677), .ZN(new_n678));
  OAI211_X1 g542(.A(new_n292), .B(new_n512), .C1(new_n291), .C2(new_n285), .ZN(new_n679));
  NAND2_X1  g543(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g544(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g545(.A1(new_n302), .A2(new_n307), .ZN(new_n682));
  AOI21_X1  g546(.A(new_n202), .B1(new_n682), .B2(new_n309), .ZN(new_n683));
  AOI21_X1  g547(.A(new_n318), .B1(new_n683), .B2(new_n308), .ZN(new_n684));
  NOR2_X1   g548(.A1(new_n684), .A2(new_n510), .ZN(new_n685));
  OAI21_X1  g549(.A(new_n685), .B1(new_n335), .B2(new_n343), .ZN(new_n686));
  OAI21_X1  g550(.A(new_n339), .B1(new_n684), .B2(new_n331), .ZN(new_n687));
  OAI21_X1  g551(.A(KEYINPUT37), .B1(new_n687), .B2(new_n685), .ZN(new_n688));
  NAND2_X1  g552(.A1(new_n320), .A2(new_n332), .ZN(RLL_wire_A_105));
  XOR2_X1 RLL_XOR_105 (.A(RLL_wire_A_105), .B(KEYINPUT105), .Z(new_n689) );
  INV_X1    g553(.A(new_n510), .ZN(new_n690));
  NAND2_X1  g554(.A1(new_n320), .A2(new_n690), .ZN(new_n691));
  INV_X1    g555(.A(KEYINPUT37), .ZN(new_n692));
  NAND4_X1  g556(.A1(new_n689), .A2(new_n691), .A3(new_n692), .A4(new_n339), .ZN(new_n693));
  NAND2_X1  g557(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g558(.A1(new_n686), .A2(KEYINPUT38), .A3(new_n694), .ZN(RLL_wire_A_106));
  XNOR2_X1 RLL_XNOR_106 (.A(RLL_wire_A_106), .B(KEYINPUT106), .ZN(new_n695) );
  AOI21_X1  g559(.A(KEYINPUT38), .B1(new_n686), .B2(new_n694), .ZN(new_n696));
  NOR2_X1   g560(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI22_X1  g561(.A1(new_n681), .A2(new_n697), .B1(new_n500), .B2(new_n690), .ZN(new_n698));
  NOR2_X1   g562(.A1(new_n676), .A2(new_n512), .ZN(new_n699));
  OAI21_X1  g563(.A(KEYINPUT39), .B1(new_n695), .B2(new_n696), .ZN(new_n700));
  INV_X1    g564(.A(KEYINPUT38), .ZN(new_n701));
  AND3_X1   g565(.A1(new_n316), .A2(new_n319), .A3(new_n338), .ZN(new_n702));
  NOR2_X1   g566(.A1(new_n702), .A2(new_n499), .ZN(new_n703));
  AOI21_X1  g567(.A(new_n692), .B1(new_n703), .B2(new_n691), .ZN(new_n704));
  INV_X1    g568(.A(new_n693), .ZN(new_n705));
  NOR2_X1   g569(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g570(.A1(new_n340), .A2(new_n342), .ZN(new_n707));
  AOI21_X1  g571(.A(new_n691), .B1(new_n500), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g572(.A(new_n701), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g573(.A(KEYINPUT39), .ZN(new_n710));
  NAND3_X1  g574(.A1(new_n686), .A2(KEYINPUT38), .A3(new_n694), .ZN(new_n711));
  NAND3_X1  g575(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g576(.A1(new_n700), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g577(.A(new_n698), .B1(new_n699), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g578(.A1(new_n554), .A2(new_n345), .A3(new_n563), .ZN(new_n715));
  AND2_X1   g579(.A1(new_n715), .A2(new_n505), .ZN(new_n716));
  XNOR2_X1  g580(.A(new_n714), .B(new_n716), .ZN(new_n717));
  INV_X1    g581(.A(KEYINPUT40), .ZN(new_n718));
  NAND2_X1  g582(.A1(new_n547), .A2(new_n512), .ZN(new_n719));
  NAND2_X1  g583(.A1(new_n719), .A2(new_n534), .ZN(new_n720));
  NAND3_X1  g584(.A1(new_n547), .A2(KEYINPUT31), .A3(new_n512), .ZN(new_n721));
  NAND3_X1  g585(.A1(new_n550), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g586(.A1(new_n722), .A2(new_n680), .A3(new_n656), .ZN(new_n723));
  OAI21_X1  g587(.A(new_n718), .B1(new_n697), .B2(new_n723), .ZN(new_n724));
  AND3_X1   g588(.A1(new_n722), .A2(new_n680), .A3(new_n656), .ZN(new_n725));
  NAND2_X1  g589(.A1(new_n709), .A2(new_n711), .ZN(new_n726));
  NAND3_X1  g590(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT40), .ZN(new_n727));
  NAND2_X1  g591(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g592(.A1(new_n345), .A2(new_n722), .ZN(new_n729));
  AOI21_X1  g593(.A(new_n518), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g594(.A(new_n730), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  OAI22_X1  g595(.A1(new_n717), .A2(new_n731), .B1(new_n188), .B2(new_n568), .ZN(new_n732));
  AND2_X1   g596(.A1(new_n717), .A2(new_n731), .ZN(new_n733));
  OAI21_X1  g597(.A(new_n672), .B1(new_n732), .B2(new_n733), .ZN(G367));
  NAND2_X1  g598(.A1(new_n483), .A2(new_n512), .ZN(new_n735));
  OR2_X1    g599(.A1(new_n491), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g600(.A1(new_n485), .A2(new_n735), .ZN(new_n737));
  NAND2_X1  g601(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g602(.A(new_n738), .ZN(new_n739));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n740));
  NAND2_X1  g604(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g605(.A(new_n560), .B1(new_n359), .B2(new_n526), .ZN(new_n742));
  OR3_X1    g606(.A1(new_n492), .A2(new_n359), .A3(new_n526), .ZN(new_n743));
  NAND2_X1  g607(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g608(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g609(.A(new_n384), .B1(new_n745), .B2(new_n472), .ZN(new_n746));
  NAND3_X1  g610(.A1(new_n523), .A2(new_n744), .A3(new_n525), .ZN(new_n747));
  AOI22_X1  g611(.A1(new_n746), .A2(new_n526), .B1(KEYINPUT42), .B2(new_n747), .ZN(new_n748));
  OR2_X1    g612(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g613(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g614(.A1(new_n738), .A2(KEYINPUT43), .ZN(new_n751));
  AOI21_X1  g615(.A(new_n741), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g616(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g617(.A1(new_n524), .A2(new_n745), .ZN(new_n754));
  NAND3_X1  g618(.A1(new_n750), .A2(new_n741), .A3(new_n751), .ZN(new_n755));
  AND3_X1   g619(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g620(.A(new_n754), .B1(new_n753), .B2(new_n755), .ZN(new_n757));
  NOR2_X1   g621(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g622(.A(new_n530), .B(KEYINPUT41), .ZN(new_n759));
  NAND2_X1  g623(.A1(new_n527), .A2(new_n744), .ZN(new_n760));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n761));
  XNOR2_X1  g625(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g626(.A(KEYINPUT44), .ZN(RLL_wire_A_107));
  XOR2_X1 RLL_XOR_107 (.A(RLL_wire_A_107), .B(KEYINPUT107), .Z(new_n763) );
  OR3_X1    g627(.A1(new_n527), .A2(new_n763), .A3(new_n744), .ZN(new_n764));
  OAI21_X1  g628(.A(new_n763), .B1(new_n527), .B2(new_n744), .ZN(new_n765));
  NAND2_X1  g629(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g630(.A1(new_n762), .A2(new_n766), .ZN(RLL_wire_A_108));
  XNOR2_X1 RLL_XNOR_108 (.A(RLL_wire_A_108), .B(KEYINPUT108), .ZN(new_n767) );
  INV_X1    g631(.A(new_n524), .ZN(new_n768));
  NAND2_X1  g632(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g633(.A1(new_n523), .A2(new_n525), .ZN(new_n770));
  NAND2_X1  g634(.A1(new_n523), .A2(new_n525), .ZN(new_n771));
  NAND2_X1  g635(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g636(.A1(new_n567), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g637(.A1(new_n519), .A2(new_n771), .A3(new_n770), .ZN(new_n774));
  NAND3_X1  g638(.A1(new_n773), .A2(new_n564), .A3(new_n774), .ZN(new_n775));
  INV_X1    g639(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g640(.A1(new_n762), .A2(new_n766), .A3(new_n524), .ZN(new_n777));
  NAND3_X1  g641(.A1(new_n769), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g642(.A(new_n759), .B1(new_n778), .B2(new_n564), .ZN(new_n779));
  NAND2_X1  g643(.A1(new_n569), .A2(G1), .ZN(new_n780));
  OAI21_X1  g644(.A(new_n758), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI221_X1 g645(.A(new_n585), .B1(new_n143), .B2(new_n232), .C1(new_n172), .C2(new_n577), .ZN(new_n782));
  NAND2_X1  g646(.A1(new_n782), .A2(new_n572), .ZN(new_n783));
  OAI22_X1  g647(.A1(new_n593), .A2(new_n636), .B1(new_n611), .B2(new_n225), .ZN(new_n784));
  INV_X1    g648(.A(G311), .ZN(new_n785));
  OAI22_X1  g649(.A1(new_n591), .A2(new_n420), .B1(new_n615), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g650(.A1(new_n619), .A2(KEYINPUT46), .A3(G116), .ZN(new_n787));
  INV_X1    g651(.A(KEYINPUT46), .ZN(new_n788));
  OAI21_X1  g652(.A(new_n788), .B1(new_n605), .B2(new_n392), .ZN(new_n789));
  OAI211_X1 g653(.A(new_n787), .B(new_n789), .C1(new_n635), .C2(new_n462), .ZN(new_n790));
  INV_X1    g654(.A(G317), .ZN(new_n791));
  OAI221_X1 g655(.A(new_n298), .B1(new_n600), .B2(new_n791), .C1(new_n348), .C2(new_n607), .ZN(new_n792));
  NOR4_X1   g656(.A1(new_n784), .A2(new_n786), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  AOI22_X1  g657(.A1(new_n590), .A2(G150), .B1(G68), .B2(new_n612), .ZN(new_n794));
  OAI21_X1  g658(.A(new_n794), .B1(new_n644), .B2(new_n615), .ZN(new_n795));
  OAI22_X1  g659(.A1(new_n593), .A2(new_n138), .B1(new_n635), .B2(new_n601), .ZN(new_n796));
  OAI21_X1  g660(.A(new_n192), .B1(new_n607), .B2(new_n156), .ZN(new_n797));
  INV_X1    g661(.A(G137), .ZN(new_n798));
  OAI22_X1  g662(.A1(new_n605), .A2(new_n203), .B1(new_n600), .B2(new_n798), .ZN(new_n799));
  NOR4_X1   g663(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g664(.A1(new_n793), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g665(.A(new_n801), .B(KEYINPUT47), .Z(new_n802));
  AOI21_X1  g666(.A(new_n783), .B1(new_n802), .B2(new_n584), .ZN(new_n803));
  OAI21_X1  g667(.A(new_n803), .B1(new_n628), .B2(new_n738), .ZN(new_n804));
  NAND2_X1  g668(.A1(new_n781), .A2(new_n804), .ZN(G387));
  NAND3_X1  g669(.A1(new_n773), .A2(new_n780), .A3(new_n774), .ZN(new_n806));
  OAI22_X1  g670(.A1(new_n573), .A2(new_n529), .B1(G107), .B2(new_n143), .ZN(new_n807));
  OR2_X1    g671(.A1(new_n169), .A2(new_n182), .ZN(new_n808));
  INV_X1    g672(.A(new_n529), .ZN(new_n809));
  AOI211_X1 g673(.A(G45), .B(new_n809), .C1(G68), .C2(G77), .ZN(new_n810));
  NOR2_X1   g674(.A1(new_n229), .A2(G50), .ZN(new_n811));
  XNOR2_X1  g675(.A(new_n811), .B(KEYINPUT50), .ZN(new_n812));
  AOI21_X1  g676(.A(new_n577), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g677(.A(new_n807), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g678(.A(new_n572), .B1(new_n814), .B2(new_n586), .ZN(new_n815));
  INV_X1    g679(.A(G150), .ZN(new_n816));
  OAI22_X1  g680(.A1(new_n605), .A2(new_n156), .B1(new_n600), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g681(.A(new_n298), .B(new_n817), .C1(G97), .C2(new_n608), .ZN(new_n818));
  NAND2_X1  g682(.A1(new_n596), .A2(G159), .ZN(RLL_wire_A_109));
  XOR2_X1 RLL_XOR_109 (.A(RLL_wire_A_109), .B(KEYINPUT109), .Z(new_n819) );
  AOI22_X1  g683(.A1(new_n590), .A2(G50), .B1(new_n406), .B2(new_n612), .ZN(new_n820));
  AOI22_X1  g684(.A1(G68), .A2(new_n592), .B1(new_n610), .B2(new_n207), .ZN(new_n821));
  NAND4_X1  g685(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  OAI22_X1  g686(.A1(new_n605), .A2(new_n462), .B1(new_n611), .B2(new_n636), .ZN(new_n823));
  OAI22_X1  g687(.A1(new_n420), .A2(new_n593), .B1(new_n591), .B2(new_n791), .ZN(new_n824));
  INV_X1    g688(.A(G322), .ZN(new_n825));
  OAI22_X1  g689(.A1(new_n635), .A2(new_n785), .B1(new_n615), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g690(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g691(.A(new_n823), .B1(new_n827), .B2(KEYINPUT48), .ZN(new_n828));
  OAI21_X1  g692(.A(new_n828), .B1(KEYINPUT48), .B2(new_n827), .ZN(new_n829));
  XOR2_X1   g693(.A(new_n829), .B(KEYINPUT49), .Z(new_n830));
  OAI221_X1 g694(.A(new_n298), .B1(new_n600), .B2(new_n616), .C1(new_n392), .C2(new_n607), .ZN(new_n831));
  OAI21_X1  g695(.A(new_n822), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g696(.A(new_n815), .B1(new_n832), .B2(new_n584), .ZN(RLL_wire_A_110));
  XOR2_X1 RLL_XOR_110 (.A(RLL_wire_A_110), .B(KEYINPUT110), .Z(new_n833) );
  OAI21_X1  g697(.A(new_n833), .B1(new_n523), .B2(new_n628), .ZN(new_n834));
  INV_X1    g698(.A(new_n530), .ZN(new_n835));
  NAND2_X1  g699(.A1(new_n775), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g700(.A(new_n564), .B1(new_n773), .B2(new_n774), .ZN(new_n837));
  OAI211_X1 g701(.A(new_n806), .B(new_n834), .C1(new_n836), .C2(new_n837), .ZN(G393));
  INV_X1    g702(.A(new_n777), .ZN(new_n839));
  AOI21_X1  g703(.A(new_n524), .B1(new_n762), .B2(new_n766), .ZN(new_n840));
  NOR2_X1   g704(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g705(.A1(new_n745), .A2(new_n582), .ZN(RLL_wire_A_111));
  XOR2_X1 RLL_XOR_111 (.A(RLL_wire_A_111), .B(KEYINPUT111), .Z(new_n842) );
  OAI221_X1 g706(.A(new_n585), .B1(new_n348), .B2(new_n143), .C1(new_n179), .C2(new_n577), .ZN(new_n843));
  NAND2_X1  g707(.A1(new_n843), .A2(new_n572), .ZN(new_n844));
  AOI22_X1  g708(.A1(G159), .A2(new_n590), .B1(new_n596), .B2(G150), .ZN(new_n845));
  XOR2_X1   g709(.A(new_n845), .B(KEYINPUT51), .Z(new_n846));
  OAI22_X1  g710(.A1(new_n605), .A2(new_n154), .B1(new_n600), .B2(new_n644), .ZN(new_n847));
  AOI211_X1 g711(.A(new_n298), .B(new_n847), .C1(G87), .C2(new_n608), .ZN(new_n848));
  OAI22_X1  g712(.A1(new_n593), .A2(new_n229), .B1(new_n635), .B2(new_n138), .ZN(new_n849));
  AOI21_X1  g713(.A(new_n849), .B1(G77), .B2(new_n612), .ZN(new_n850));
  NAND3_X1  g714(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  AOI22_X1  g715(.A1(G311), .A2(new_n590), .B1(new_n596), .B2(G317), .ZN(new_n852));
  XOR2_X1   g716(.A(new_n852), .B(KEYINPUT52), .Z(new_n853));
  OAI22_X1  g717(.A1(new_n605), .A2(new_n636), .B1(new_n600), .B2(new_n825), .ZN(new_n854));
  AOI211_X1 g718(.A(new_n192), .B(new_n854), .C1(G107), .C2(new_n608), .ZN(new_n855));
  OAI22_X1  g719(.A1(new_n635), .A2(new_n420), .B1(new_n611), .B2(new_n392), .ZN(new_n856));
  AOI21_X1  g720(.A(new_n856), .B1(G294), .B2(new_n592), .ZN(new_n857));
  NAND3_X1  g721(.A1(new_n853), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g722(.A1(new_n851), .A2(new_n858), .ZN(RLL_wire_A_112));
  XNOR2_X1 RLL_XNOR_112 (.A(RLL_wire_A_112), .B(KEYINPUT112), .ZN(new_n859) );
  AOI21_X1  g723(.A(new_n844), .B1(new_n859), .B2(new_n584), .ZN(new_n860));
  AOI22_X1  g724(.A1(new_n841), .A2(new_n780), .B1(new_n842), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g725(.A(new_n775), .B1(new_n839), .B2(new_n840), .ZN(new_n862));
  NAND3_X1  g726(.A1(new_n862), .A2(new_n778), .A3(new_n835), .ZN(new_n863));
  NAND2_X1  g727(.A1(new_n861), .A2(new_n863), .ZN(G390));
  INV_X1    g728(.A(new_n699), .ZN(new_n865));
  AOI21_X1  g729(.A(new_n673), .B1(new_n562), .B2(new_n656), .ZN(new_n866));
  INV_X1    g730(.A(new_n680), .ZN(new_n867));
  OAI211_X1 g731(.A(new_n726), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(RLL_wire_A_113));
  XOR2_X1 RLL_XOR_113 (.A(RLL_wire_A_113), .B(KEYINPUT113), .Z(new_n868) );
  AOI21_X1  g732(.A(new_n699), .B1(new_n675), .B2(new_n680), .ZN(new_n869));
  OAI21_X1  g733(.A(new_n868), .B1(new_n713), .B2(new_n869), .ZN(new_n870));
  AND4_X1   g734(.A1(G330), .A2(new_n722), .A3(new_n680), .A4(new_n656), .ZN(new_n871));
  NAND2_X1  g735(.A1(new_n870), .A2(new_n871), .ZN(RLL_wire_A_114));
  XOR2_X1 RLL_XOR_114 (.A(RLL_wire_A_114), .B(KEYINPUT114), .Z(new_n872) );
  NAND3_X1  g736(.A1(new_n551), .A2(new_n656), .A3(new_n680), .ZN(new_n873));
  OAI211_X1 g737(.A(new_n868), .B(new_n873), .C1(new_n713), .C2(new_n869), .ZN(new_n874));
  NAND3_X1  g738(.A1(new_n345), .A2(G330), .A3(new_n722), .ZN(new_n875));
  NAND3_X1  g739(.A1(new_n715), .A2(new_n505), .A3(new_n875), .ZN(RLL_wire_A_115));
  XOR2_X1 RLL_XOR_115 (.A(RLL_wire_A_115), .B(KEYINPUT115), .Z(new_n876) );
  AOI21_X1  g740(.A(new_n680), .B1(new_n551), .B2(new_n656), .ZN(new_n877));
  OAI21_X1  g741(.A(new_n675), .B1(new_n877), .B2(new_n871), .ZN(new_n878));
  NAND2_X1  g742(.A1(new_n722), .A2(G330), .ZN(new_n879));
  OAI21_X1  g743(.A(new_n867), .B1(new_n879), .B2(new_n658), .ZN(new_n880));
  NAND3_X1  g744(.A1(new_n880), .A2(new_n866), .A3(new_n873), .ZN(new_n881));
  AOI21_X1  g745(.A(new_n876), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g746(.A1(new_n872), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g747(.A1(new_n883), .A2(new_n835), .ZN(new_n884));
  NAND2_X1  g748(.A1(new_n872), .A2(new_n874), .ZN(new_n885));
  INV_X1    g749(.A(new_n882), .ZN(new_n886));
  NAND2_X1  g750(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g751(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g752(.A1(new_n872), .A2(new_n780), .A3(new_n874), .ZN(new_n889));
  OAI21_X1  g753(.A(new_n572), .B1(new_n207), .B2(new_n633), .ZN(new_n890));
  XNOR2_X1  g754(.A(KEYINPUT54), .B(G143), .ZN(new_n891));
  OAI22_X1  g755(.A1(new_n593), .A2(new_n891), .B1(new_n635), .B2(new_n798), .ZN(new_n892));
  AOI21_X1  g756(.A(new_n892), .B1(G159), .B2(new_n612), .ZN(new_n893));
  OAI21_X1  g757(.A(new_n192), .B1(new_n607), .B2(new_n138), .ZN(new_n894));
  AOI21_X1  g758(.A(new_n894), .B1(G125), .B2(new_n621), .ZN(RLL_wire_A_116));
  XNOR2_X1 RLL_XNOR_116 (.A(RLL_wire_A_116), .B(KEYINPUT116), .ZN(new_n895) );
  AOI22_X1  g759(.A1(G132), .A2(new_n590), .B1(new_n596), .B2(G128), .ZN(new_n896));
  NOR2_X1   g760(.A1(new_n605), .A2(new_n816), .ZN(new_n897));
  XNOR2_X1  g761(.A(new_n897), .B(KEYINPUT53), .ZN(new_n898));
  NAND4_X1  g762(.A1(new_n893), .A2(new_n895), .A3(new_n896), .A4(new_n898), .ZN(RLL_wire_A_117));
  XNOR2_X1 RLL_XNOR_117 (.A(RLL_wire_A_117), .B(KEYINPUT117), .ZN(new_n899) );
  OAI22_X1  g763(.A1(new_n593), .A2(new_n348), .B1(new_n635), .B2(new_n225), .ZN(new_n900));
  AOI21_X1  g764(.A(new_n900), .B1(G283), .B2(new_n596), .ZN(new_n901));
  AOI21_X1  g765(.A(new_n192), .B1(new_n619), .B2(G87), .ZN(new_n902));
  AOI22_X1  g766(.A1(new_n608), .A2(G68), .B1(new_n621), .B2(G294), .ZN(new_n903));
  AOI22_X1  g767(.A1(new_n590), .A2(G116), .B1(G77), .B2(new_n612), .ZN(new_n904));
  NAND4_X1  g768(.A1(new_n901), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g769(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g770(.A(new_n890), .B1(new_n906), .B2(new_n584), .ZN(new_n907));
  OAI21_X1  g771(.A(new_n907), .B1(new_n713), .B2(new_n581), .ZN(new_n908));
  NAND2_X1  g772(.A1(new_n889), .A2(new_n908), .ZN(new_n909));
  INV_X1    g773(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g774(.A1(new_n888), .A2(new_n910), .ZN(G378));
  NOR2_X1   g775(.A1(G33), .A2(G41), .ZN(new_n912));
  AOI211_X1 g776(.A(G50), .B(new_n912), .C1(new_n298), .C2(new_n181), .ZN(new_n913));
  NOR2_X1   g777(.A1(new_n607), .A2(new_n203), .ZN(RLL_wire_A_118));
  XOR2_X1 RLL_XOR_118 (.A(RLL_wire_A_118), .B(KEYINPUT118), .Z(new_n914) );
  OAI211_X1 g778(.A(new_n181), .B(new_n298), .C1(new_n605), .C2(new_n156), .ZN(new_n915));
  AOI211_X1 g779(.A(new_n914), .B(new_n915), .C1(G283), .C2(new_n621), .ZN(new_n916));
  NAND2_X1  g780(.A1(new_n590), .A2(G107), .ZN(new_n917));
  AOI22_X1  g781(.A1(new_n406), .A2(new_n592), .B1(new_n610), .B2(G97), .ZN(new_n918));
  AOI22_X1  g782(.A1(new_n596), .A2(G116), .B1(G68), .B2(new_n612), .ZN(new_n919));
  NAND4_X1  g783(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  INV_X1    g784(.A(KEYINPUT58), .ZN(RLL_wire_A_119));
  XOR2_X1 RLL_XOR_119 (.A(RLL_wire_A_119), .B(KEYINPUT119), .Z(new_n921) );
  AOI21_X1  g785(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g786(.A1(G137), .A2(new_n592), .B1(new_n610), .B2(G132), .ZN(new_n923));
  NOR2_X1   g787(.A1(new_n605), .A2(new_n891), .ZN(new_n924));
  AOI21_X1  g788(.A(new_n924), .B1(new_n590), .B2(G128), .ZN(new_n925));
  AOI22_X1  g789(.A1(new_n596), .A2(G125), .B1(G150), .B2(new_n612), .ZN(new_n926));
  NAND3_X1  g790(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g791(.A(new_n927), .B(KEYINPUT59), .ZN(new_n928));
  INV_X1    g792(.A(G124), .ZN(new_n929));
  OAI221_X1 g793(.A(new_n912), .B1(new_n600), .B2(new_n929), .C1(new_n601), .C2(new_n607), .ZN(RLL_wire_A_120));
  XOR2_X1 RLL_XOR_120 (.A(RLL_wire_A_120), .B(KEYINPUT120), .Z(new_n930) );
  OAI221_X1 g794(.A(new_n922), .B1(new_n921), .B2(new_n920), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g795(.A1(new_n931), .A2(new_n584), .ZN(new_n932));
  AOI21_X1  g796(.A(new_n570), .B1(new_n138), .B2(new_n632), .ZN(new_n933));
  OAI21_X1  g797(.A(new_n504), .B1(new_n221), .B2(new_n219), .ZN(new_n934));
  NOR2_X1   g798(.A1(new_n246), .A2(new_n510), .ZN(new_n935));
  XNOR2_X1  g799(.A(new_n935), .B(KEYINPUT56), .ZN(new_n936));
  XNOR2_X1  g800(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  XNOR2_X1  g801(.A(new_n934), .B(new_n937), .ZN(new_n938));
  INV_X1    g802(.A(new_n938), .ZN(new_n939));
  OAI211_X1 g803(.A(new_n932), .B(new_n933), .C1(new_n939), .C2(new_n581), .ZN(new_n940));
  INV_X1    g804(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g805(.A1(new_n724), .A2(G330), .A3(new_n727), .ZN(new_n942));
  NAND2_X1  g806(.A1(new_n942), .A2(new_n938), .ZN(new_n943));
  NAND4_X1  g807(.A1(new_n724), .A2(G330), .A3(new_n727), .A4(new_n939), .ZN(new_n944));
  NAND2_X1  g808(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g809(.A(new_n714), .ZN(new_n946));
  NAND2_X1  g810(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g811(.A1(new_n714), .A2(new_n943), .A3(new_n944), .ZN(new_n948));
  NAND2_X1  g812(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g813(.A(new_n941), .B1(new_n949), .B2(new_n780), .ZN(new_n950));
  INV_X1    g814(.A(new_n876), .ZN(new_n951));
  NAND2_X1  g815(.A1(new_n883), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g816(.A1(new_n714), .A2(new_n943), .A3(new_n944), .ZN(new_n953));
  AOI21_X1  g817(.A(new_n714), .B1(new_n944), .B2(new_n943), .ZN(new_n954));
  OAI211_X1 g818(.A(new_n952), .B(KEYINPUT57), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g819(.A1(new_n955), .A2(new_n835), .ZN(new_n956));
  AOI21_X1  g820(.A(KEYINPUT57), .B1(new_n949), .B2(new_n952), .ZN(new_n957));
  OAI21_X1  g821(.A(new_n950), .B1(new_n956), .B2(new_n957), .ZN(G375));
  INV_X1    g822(.A(new_n759), .ZN(RLL_wire_A_121));
  XNOR2_X1 RLL_XNOR_121 (.A(RLL_wire_A_121), .B(KEYINPUT121), .ZN(new_n959) );
  NAND3_X1  g823(.A1(new_n878), .A2(new_n881), .A3(new_n876), .ZN(RLL_wire_A_122));
  XNOR2_X1 RLL_XNOR_122 (.A(RLL_wire_A_122), .B(KEYINPUT122), .ZN(new_n960) );
  NAND3_X1  g824(.A1(new_n886), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g825(.A(new_n780), .ZN(new_n962));
  AOI21_X1  g826(.A(new_n962), .B1(new_n878), .B2(new_n881), .ZN(RLL_wire_A_123));
  XOR2_X1 RLL_XOR_123 (.A(RLL_wire_A_123), .B(KEYINPUT123), .Z(new_n963) );
  NAND2_X1  g827(.A1(new_n867), .A2(new_n580), .ZN(new_n964));
  OAI21_X1  g828(.A(new_n572), .B1(G68), .B2(new_n633), .ZN(new_n965));
  OAI22_X1  g829(.A1(new_n593), .A2(new_n225), .B1(new_n635), .B2(new_n392), .ZN(new_n966));
  AOI21_X1  g830(.A(new_n966), .B1(G294), .B2(new_n596), .ZN(new_n967));
  AOI21_X1  g831(.A(new_n192), .B1(new_n608), .B2(G77), .ZN(new_n968));
  AOI22_X1  g832(.A1(new_n619), .A2(G97), .B1(new_n621), .B2(G303), .ZN(new_n969));
  AOI22_X1  g833(.A1(new_n590), .A2(G283), .B1(new_n406), .B2(new_n612), .ZN(new_n970));
  NAND4_X1  g834(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g835(.A1(new_n596), .A2(G132), .ZN(new_n972));
  OAI221_X1 g836(.A(new_n972), .B1(new_n635), .B2(new_n891), .C1(new_n798), .C2(new_n591), .ZN(new_n973));
  AOI22_X1  g837(.A1(new_n592), .A2(G150), .B1(G50), .B2(new_n612), .ZN(new_n974));
  NOR2_X1   g838(.A1(new_n914), .A2(new_n298), .ZN(new_n975));
  AOI22_X1  g839(.A1(new_n619), .A2(G159), .B1(new_n621), .B2(G128), .ZN(new_n976));
  NAND3_X1  g840(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g841(.A(new_n971), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g842(.A(new_n965), .B1(new_n978), .B2(new_n584), .ZN(RLL_wire_A_124));
  XOR2_X1 RLL_XOR_124 (.A(RLL_wire_A_124), .B(KEYINPUT124), .Z(new_n979) );
  AOI21_X1  g843(.A(new_n963), .B1(new_n964), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g844(.A1(new_n961), .A2(new_n980), .ZN(G381));
  OR3_X1    g845(.A1(G393), .A2(G396), .A3(G384), .ZN(RLL_wire_A_125));
  XOR2_X1 RLL_XOR_125 (.A(RLL_wire_A_125), .B(KEYINPUT125), .Z(new_n982) );
  NOR4_X1   g846(.A1(G387), .A2(G390), .A3(G381), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g847(.A(new_n909), .B1(new_n884), .B2(new_n887), .ZN(new_n984));
  INV_X1    g848(.A(G375), .ZN(new_n985));
  NAND3_X1  g849(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(G407));
  NAND2_X1  g850(.A1(new_n511), .A2(G213), .ZN(new_n987));
  INV_X1    g851(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g852(.A1(new_n985), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g853(.A1(G407), .A2(G213), .A3(new_n989), .ZN(G409));
  OAI211_X1 g854(.A(G378), .B(new_n950), .C1(new_n956), .C2(new_n957), .ZN(new_n991));
  AND3_X1   g855(.A1(new_n949), .A2(new_n959), .A3(new_n952), .ZN(new_n992));
  NOR2_X1   g856(.A1(new_n953), .A2(new_n954), .ZN(new_n993));
  OAI21_X1  g857(.A(new_n940), .B1(new_n993), .B2(new_n962), .ZN(new_n994));
  OAI21_X1  g858(.A(new_n984), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g859(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  INV_X1    g860(.A(KEYINPUT60), .ZN(new_n997));
  OAI21_X1  g861(.A(new_n960), .B1(new_n882), .B2(new_n997), .ZN(new_n998));
  NAND4_X1  g862(.A1(new_n878), .A2(new_n881), .A3(new_n876), .A4(KEYINPUT60), .ZN(new_n999));
  NAND3_X1  g863(.A1(new_n998), .A2(new_n835), .A3(new_n999), .ZN(new_n1000));
  AND3_X1   g864(.A1(new_n1000), .A2(G384), .A3(new_n980), .ZN(new_n1001));
  AOI21_X1  g865(.A(G384), .B1(new_n1000), .B2(new_n980), .ZN(new_n1002));
  NOR2_X1   g866(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g867(.A1(new_n996), .A2(new_n987), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g868(.A(KEYINPUT63), .ZN(new_n1005));
  NAND2_X1  g869(.A1(new_n1004), .A2(new_n1005), .ZN(RLL_wire_A_126));
  XNOR2_X1 RLL_XNOR_126 (.A(RLL_wire_A_126), .B(KEYINPUT126), .ZN(new_n1006) );
  NAND2_X1  g870(.A1(new_n996), .A2(new_n987), .ZN(new_n1007));
  INV_X1    g871(.A(G2897), .ZN(new_n1008));
  OAI21_X1  g872(.A(new_n1003), .B1(new_n1008), .B2(new_n987), .ZN(new_n1009));
  OAI211_X1 g873(.A(G2897), .B(new_n988), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1010));
  NAND2_X1  g874(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g875(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g876(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g877(.A(G393), .B(G396), .ZN(new_n1014));
  INV_X1    g878(.A(new_n1014), .ZN(new_n1015));
  AND3_X1   g879(.A1(new_n781), .A2(new_n804), .A3(G390), .ZN(new_n1016));
  AOI21_X1  g880(.A(G390), .B1(new_n781), .B2(new_n804), .ZN(new_n1017));
  OAI21_X1  g881(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g882(.A(G390), .ZN(new_n1019));
  NAND2_X1  g883(.A1(G387), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g884(.A1(new_n781), .A2(new_n804), .A3(G390), .ZN(new_n1021));
  NAND3_X1  g885(.A1(new_n1020), .A2(new_n1021), .A3(new_n1014), .ZN(new_n1022));
  AOI21_X1  g886(.A(KEYINPUT61), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g887(.A(new_n988), .B1(new_n991), .B2(new_n995), .ZN(new_n1024));
  NAND3_X1  g888(.A1(new_n1024), .A2(KEYINPUT63), .A3(new_n1003), .ZN(new_n1025));
  NAND4_X1  g889(.A1(new_n1006), .A2(new_n1013), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g890(.A(KEYINPUT61), .ZN(RLL_wire_A_127));
  XOR2_X1 RLL_XOR_127 (.A(RLL_wire_A_127), .B(KEYINPUT127), .Z(new_n1027) );
  OAI21_X1  g891(.A(new_n1027), .B1(new_n1024), .B2(new_n1011), .ZN(new_n1028));
  INV_X1    g892(.A(KEYINPUT62), .ZN(new_n1029));
  NAND2_X1  g893(.A1(new_n1004), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g894(.A1(new_n1024), .A2(KEYINPUT62), .A3(new_n1003), .ZN(new_n1031));
  AOI21_X1  g895(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g896(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1033));
  INV_X1    g897(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g898(.A(new_n1026), .B1(new_n1032), .B2(new_n1034), .ZN(G405));
  NAND2_X1  g899(.A1(G375), .A2(new_n984), .ZN(new_n1036));
  NAND2_X1  g900(.A1(new_n1036), .A2(new_n991), .ZN(new_n1037));
  NAND2_X1  g901(.A1(new_n1037), .A2(new_n1003), .ZN(new_n1038));
  OAI211_X1 g902(.A(new_n1036), .B(new_n991), .C1(new_n1002), .C2(new_n1001), .ZN(new_n1039));
  AND3_X1   g903(.A1(new_n1033), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g904(.A(new_n1033), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1041));
  NOR2_X1   g905(.A1(new_n1040), .A2(new_n1041), .ZN(G402));

endmodule
