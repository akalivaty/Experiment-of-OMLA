

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577;

  XNOR2_X1 U320 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n390) );
  XNOR2_X1 U321 ( .A(n394), .B(KEYINPUT47), .ZN(n395) );
  XNOR2_X1 U322 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U323 ( .A(G99GAT), .B(G85GAT), .Z(n343) );
  XOR2_X1 U324 ( .A(KEYINPUT48), .B(n399), .Z(n544) );
  NOR2_X1 U325 ( .A1(n572), .A2(n492), .ZN(n493) );
  XNOR2_X1 U326 ( .A(n338), .B(n303), .ZN(n304) );
  XOR2_X1 U327 ( .A(n445), .B(n444), .Z(n288) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U329 ( .A(n430), .B(KEYINPUT95), .Z(n290) );
  XNOR2_X1 U330 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n429) );
  XOR2_X1 U331 ( .A(G50GAT), .B(G162GAT), .Z(n440) );
  XNOR2_X1 U332 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U333 ( .A(n391), .B(n390), .ZN(n393) );
  XNOR2_X1 U334 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U335 ( .A(n295), .B(n289), .ZN(n296) );
  XNOR2_X1 U336 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U337 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U338 ( .A(n359), .B(n358), .ZN(n388) );
  NOR2_X1 U339 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U340 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U341 ( .A(n305), .B(n304), .ZN(n360) );
  XNOR2_X1 U342 ( .A(n452), .B(n451), .ZN(n469) );
  NOR2_X1 U343 ( .A1(n528), .A2(n454), .ZN(n560) );
  XOR2_X1 U344 ( .A(n322), .B(n426), .Z(n528) );
  XNOR2_X1 U345 ( .A(n496), .B(n495), .ZN(n504) );
  XNOR2_X1 U346 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n455) );
  XNOR2_X1 U347 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U348 ( .A(n343), .B(n440), .Z(n292) );
  XNOR2_X1 U349 ( .A(G134GAT), .B(G218GAT), .ZN(n291) );
  XNOR2_X1 U350 ( .A(n292), .B(n291), .ZN(n297) );
  XOR2_X1 U351 ( .A(KEYINPUT10), .B(KEYINPUT80), .Z(n294) );
  XNOR2_X1 U352 ( .A(G106GAT), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U353 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U354 ( .A(n298), .B(KEYINPUT9), .Z(n305) );
  XOR2_X1 U355 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n300) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G29GAT), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U358 ( .A(KEYINPUT71), .B(n301), .Z(n338) );
  XNOR2_X1 U359 ( .A(G36GAT), .B(G190GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n302), .B(KEYINPUT81), .ZN(n407) );
  XNOR2_X1 U361 ( .A(n407), .B(KEYINPUT11), .ZN(n303) );
  INV_X1 U362 ( .A(n360), .ZN(n540) );
  XOR2_X1 U363 ( .A(G120GAT), .B(G71GAT), .Z(n347) );
  XOR2_X1 U364 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n307) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n307), .B(n306), .ZN(n410) );
  XOR2_X1 U367 ( .A(n347), .B(n410), .Z(n309) );
  XNOR2_X1 U368 ( .A(G190GAT), .B(G99GAT), .ZN(n308) );
  XNOR2_X1 U369 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U370 ( .A(KEYINPUT91), .B(G176GAT), .Z(n311) );
  NAND2_X1 U371 ( .A1(G227GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U373 ( .A(n313), .B(n312), .Z(n318) );
  XOR2_X1 U374 ( .A(KEYINPUT20), .B(G183GAT), .Z(n315) );
  XNOR2_X1 U375 ( .A(G43GAT), .B(G15GAT), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n316), .B(KEYINPUT92), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U379 ( .A(KEYINPUT90), .B(G134GAT), .Z(n320) );
  XNOR2_X1 U380 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U382 ( .A(G113GAT), .B(n321), .Z(n426) );
  XOR2_X1 U383 ( .A(KEYINPUT66), .B(KEYINPUT69), .Z(n324) );
  XNOR2_X1 U384 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U386 ( .A(G50GAT), .B(G36GAT), .Z(n326) );
  XOR2_X1 U387 ( .A(G141GAT), .B(G22GAT), .Z(n441) );
  XOR2_X1 U388 ( .A(G15GAT), .B(G1GAT), .Z(n361) );
  XNOR2_X1 U389 ( .A(n441), .B(n361), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U391 ( .A(n328), .B(n327), .Z(n330) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U394 ( .A(G8GAT), .B(G113GAT), .Z(n332) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G197GAT), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U397 ( .A(n334), .B(n333), .Z(n340) );
  XOR2_X1 U398 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n336) );
  XNOR2_X1 U399 ( .A(KEYINPUT68), .B(KEYINPUT72), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U402 ( .A(n340), .B(n339), .Z(n530) );
  INV_X1 U403 ( .A(n530), .ZN(n564) );
  XOR2_X1 U404 ( .A(KEYINPUT32), .B(KEYINPUT78), .Z(n342) );
  XNOR2_X1 U405 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U407 ( .A(n344), .B(n343), .Z(n351) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n345), .B(G148GAT), .ZN(n448) );
  XNOR2_X1 U410 ( .A(n448), .B(KEYINPUT76), .ZN(n349) );
  AND2_X1 U411 ( .A1(G230GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n359) );
  XNOR2_X1 U413 ( .A(G176GAT), .B(G92GAT), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n352), .B(G64GAT), .ZN(n409) );
  XNOR2_X1 U415 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n353), .B(KEYINPUT73), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n409), .B(n364), .ZN(n357) );
  XOR2_X1 U418 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n355) );
  XNOR2_X1 U419 ( .A(KEYINPUT77), .B(KEYINPUT74), .ZN(n354) );
  XOR2_X1 U420 ( .A(n355), .B(n354), .Z(n356) );
  XNOR2_X1 U421 ( .A(KEYINPUT36), .B(n360), .ZN(n574) );
  XOR2_X1 U422 ( .A(G8GAT), .B(G183GAT), .Z(n404) );
  XOR2_X1 U423 ( .A(n404), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U424 ( .A(n361), .B(G155GAT), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U426 ( .A(n364), .B(KEYINPUT15), .Z(n366) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U429 ( .A(n368), .B(n367), .Z(n370) );
  XNOR2_X1 U430 ( .A(G22GAT), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U431 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U432 ( .A(KEYINPUT87), .B(G64GAT), .Z(n372) );
  XNOR2_X1 U433 ( .A(G127GAT), .B(G71GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U435 ( .A(n374), .B(n373), .Z(n382) );
  XOR2_X1 U436 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n376) );
  XNOR2_X1 U437 ( .A(KEYINPUT83), .B(KEYINPUT85), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U439 ( .A(KEYINPUT14), .B(KEYINPUT88), .Z(n378) );
  XNOR2_X1 U440 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U443 ( .A(n382), .B(n381), .Z(n536) );
  INV_X1 U444 ( .A(n536), .ZN(n572) );
  NAND2_X1 U445 ( .A1(n574), .A2(n572), .ZN(n384) );
  XOR2_X1 U446 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  NOR2_X1 U448 ( .A1(n388), .A2(n385), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n386), .B(KEYINPUT119), .ZN(n387) );
  NOR2_X1 U450 ( .A1(n564), .A2(n387), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n388), .B(KEYINPUT64), .ZN(n389) );
  XNOR2_X1 U452 ( .A(KEYINPUT41), .B(n389), .ZN(n457) );
  OR2_X1 U453 ( .A1(n457), .A2(n530), .ZN(n391) );
  NOR2_X1 U454 ( .A1(n360), .A2(n572), .ZN(n392) );
  NAND2_X1 U455 ( .A1(n393), .A2(n392), .ZN(n396) );
  XOR2_X1 U456 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n394) );
  XNOR2_X1 U457 ( .A(G211GAT), .B(G218GAT), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n400), .B(KEYINPUT94), .ZN(n401) );
  XOR2_X1 U459 ( .A(n401), .B(KEYINPUT21), .Z(n403) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(G204GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n450) );
  XOR2_X1 U462 ( .A(KEYINPUT102), .B(n404), .Z(n406) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U465 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U468 ( .A(n450), .B(n413), .Z(n518) );
  INV_X1 U469 ( .A(n518), .ZN(n414) );
  NAND2_X1 U470 ( .A1(n544), .A2(n414), .ZN(n416) );
  XOR2_X1 U471 ( .A(KEYINPUT124), .B(KEYINPUT54), .Z(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n439) );
  XOR2_X1 U473 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n418) );
  XNOR2_X1 U474 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U476 ( .A(G148GAT), .B(G120GAT), .Z(n420) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(G141GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n438) );
  XOR2_X1 U480 ( .A(G85GAT), .B(G57GAT), .Z(n424) );
  XNOR2_X1 U481 ( .A(G162GAT), .B(KEYINPUT101), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U483 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U484 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n436) );
  XOR2_X1 U486 ( .A(KEYINPUT4), .B(KEYINPUT100), .Z(n433) );
  XNOR2_X1 U487 ( .A(n429), .B(G155GAT), .ZN(n430) );
  XNOR2_X1 U488 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n290), .B(n431), .ZN(n445) );
  XNOR2_X1 U490 ( .A(n445), .B(KEYINPUT99), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U492 ( .A(G1GAT), .B(n434), .Z(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n546) );
  NAND2_X1 U495 ( .A1(n439), .A2(n546), .ZN(n562) );
  XOR2_X1 U496 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n443) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  NAND2_X1 U499 ( .A1(G228GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n288), .B(n446), .ZN(n447) );
  XOR2_X1 U501 ( .A(n447), .B(KEYINPUT23), .Z(n452) );
  XNOR2_X1 U502 ( .A(n448), .B(KEYINPUT93), .ZN(n449) );
  NOR2_X1 U503 ( .A1(n562), .A2(n469), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n360), .A2(n560), .ZN(n456) );
  INV_X1 U506 ( .A(n457), .ZN(n548) );
  NAND2_X1 U507 ( .A1(n560), .A2(n548), .ZN(n460) );
  XOR2_X1 U508 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  XNOR2_X1 U509 ( .A(n458), .B(G176GAT), .ZN(n459) );
  XNOR2_X1 U510 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  NOR2_X1 U511 ( .A1(n388), .A2(n530), .ZN(n461) );
  XOR2_X1 U512 ( .A(KEYINPUT79), .B(n461), .Z(n494) );
  XOR2_X1 U513 ( .A(KEYINPUT27), .B(n518), .Z(n466) );
  XOR2_X1 U514 ( .A(KEYINPUT28), .B(n469), .Z(n523) );
  INV_X1 U515 ( .A(n546), .ZN(n462) );
  AND2_X1 U516 ( .A1(n523), .A2(n462), .ZN(n463) );
  NAND2_X1 U517 ( .A1(n466), .A2(n463), .ZN(n527) );
  XNOR2_X1 U518 ( .A(KEYINPUT103), .B(n527), .ZN(n464) );
  NAND2_X1 U519 ( .A1(n464), .A2(n528), .ZN(n475) );
  NAND2_X1 U520 ( .A1(n469), .A2(n528), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT26), .ZN(n563) );
  INV_X1 U522 ( .A(n466), .ZN(n467) );
  NOR2_X1 U523 ( .A1(n563), .A2(n467), .ZN(n543) );
  XOR2_X1 U524 ( .A(n543), .B(KEYINPUT104), .Z(n472) );
  NOR2_X1 U525 ( .A1(n528), .A2(n518), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U527 ( .A(KEYINPUT25), .B(n470), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n473), .A2(n546), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n491) );
  NAND2_X1 U531 ( .A1(n572), .A2(n540), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT89), .B(n476), .Z(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  AND2_X1 U534 ( .A1(n491), .A2(n478), .ZN(n506) );
  NAND2_X1 U535 ( .A1(n494), .A2(n506), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT105), .B(n479), .Z(n488) );
  NOR2_X1 U537 ( .A1(n546), .A2(n488), .ZN(n481) );
  XNOR2_X1 U538 ( .A(KEYINPUT34), .B(KEYINPUT106), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U540 ( .A(G1GAT), .B(n482), .Z(G1324GAT) );
  NOR2_X1 U541 ( .A1(n518), .A2(n488), .ZN(n484) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT107), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  NOR2_X1 U544 ( .A1(n528), .A2(n488), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT35), .B(KEYINPUT108), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n523), .A2(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT109), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1327GAT) );
  XNOR2_X1 U551 ( .A(KEYINPUT110), .B(KEYINPUT38), .ZN(n496) );
  NAND2_X1 U552 ( .A1(n574), .A2(n491), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n493), .Z(n516) );
  NAND2_X1 U554 ( .A1(n516), .A2(n494), .ZN(n495) );
  NOR2_X1 U555 ( .A1(n546), .A2(n504), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n518), .A2(n504), .ZN(n499) );
  XOR2_X1 U559 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n501) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT112), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n528), .A2(n504), .ZN(n502) );
  XOR2_X1 U564 ( .A(n503), .B(n502), .Z(G1330GAT) );
  NOR2_X1 U565 ( .A1(n523), .A2(n504), .ZN(n505) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n505), .Z(G1331GAT) );
  NOR2_X1 U567 ( .A1(n564), .A2(n457), .ZN(n515) );
  NAND2_X1 U568 ( .A1(n506), .A2(n515), .ZN(n511) );
  NOR2_X1 U569 ( .A1(n546), .A2(n511), .ZN(n507) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n507), .Z(n508) );
  XNOR2_X1 U571 ( .A(KEYINPUT42), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n518), .A2(n511), .ZN(n509) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n528), .A2(n511), .ZN(n510) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n510), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U579 ( .A(G78GAT), .B(n514), .Z(G1335GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n522) );
  NOR2_X1 U581 ( .A1(n546), .A2(n522), .ZN(n517) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n522), .ZN(n519) );
  XOR2_X1 U584 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U585 ( .A1(n528), .A2(n522), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT114), .B(n520), .Z(n521) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT115), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U593 ( .A1(n544), .A2(n529), .ZN(n539) );
  NOR2_X1 U594 ( .A1(n530), .A2(n539), .ZN(n531) );
  XOR2_X1 U595 ( .A(G113GAT), .B(n531), .Z(G1340GAT) );
  NOR2_X1 U596 ( .A1(n539), .A2(n457), .ZN(n535) );
  XOR2_X1 U597 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n533) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U601 ( .A1(n536), .A2(n539), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(n537), .Z(n538) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n555), .A2(n564), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n552) );
  XOR2_X1 U612 ( .A(KEYINPUT52), .B(KEYINPUT122), .Z(n550) );
  NAND2_X1 U613 ( .A1(n555), .A2(n548), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(G155GAT), .B(KEYINPUT123), .Z(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n572), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n360), .A2(n555), .ZN(n556) );
  XNOR2_X1 U620 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n560), .A2(n564), .ZN(n558) );
  INV_X1 U622 ( .A(KEYINPUT125), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n572), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n575) );
  NAND2_X1 U628 ( .A1(n575), .A2(n564), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n566) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n575), .A2(n388), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n571), .Z(G1353GAT) );
  NAND2_X1 U637 ( .A1(n575), .A2(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT62), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(n577), .ZN(G1355GAT) );
endmodule

