//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(G355));
  NOR2_X1   g0006(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT66), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND4_X1  g0014(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n207), .B1(new_n210), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n216), .B(new_n217), .Z(new_n218));
  NOR2_X1   g0018(.A1(new_n210), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT0), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n218), .B(new_n221), .C1(new_n224), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G50), .B(G68), .Z(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n222), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n202), .A2(new_n223), .ZN(new_n248));
  XOR2_X1   g0048(.A(KEYINPUT8), .B(G58), .Z(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n223), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n223), .A2(new_n253), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n250), .A2(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n247), .B1(new_n248), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n247), .B1(new_n257), .B2(G20), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(G50), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(KEYINPUT9), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT9), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n269), .B1(new_n203), .B2(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n222), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n276), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n280), .B2(G226), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G190), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n264), .A2(new_n266), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(G200), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(KEYINPUT70), .C2(KEYINPUT10), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT10), .B1(new_n285), .B2(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n286), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT68), .B(G179), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n282), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n293), .B(new_n262), .C1(G169), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n258), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n203), .ZN(new_n297));
  INV_X1    g0097(.A(new_n260), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n203), .ZN(new_n299));
  INV_X1    g0099(.A(new_n247), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n249), .A2(new_n301), .B1(G20), .B2(G77), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT15), .B(G87), .Z(new_n303));
  NAND3_X1  g0103(.A1(new_n303), .A2(new_n223), .A3(G33), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n300), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n278), .B1(new_n280), .B2(G244), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n267), .A2(G232), .A3(new_n268), .ZN(new_n310));
  INV_X1    g0110(.A(G107), .ZN(new_n311));
  INV_X1    g0111(.A(G238), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n310), .B1(new_n311), .B2(new_n267), .C1(new_n270), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n274), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n309), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n307), .B1(new_n316), .B2(G200), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n283), .B2(new_n316), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n306), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n291), .B2(new_n316), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  AND4_X1   g0122(.A1(new_n287), .A2(new_n290), .A3(new_n295), .A4(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n249), .A2(new_n296), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n298), .B2(new_n249), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n267), .A2(G226), .A3(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT3), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G33), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n328), .A2(new_n330), .A3(G223), .A4(new_n268), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n327), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n274), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n278), .B1(new_n280), .B2(G232), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n334), .A2(new_n283), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(G200), .B1(new_n334), .B2(new_n335), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT75), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n267), .A2(new_n341), .A3(G20), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n328), .A2(new_n330), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT7), .B1(new_n343), .B2(new_n223), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G58), .A2(G68), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n223), .B1(new_n227), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G159), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n254), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT74), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(G58), .A2(G68), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G58), .A2(G68), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n301), .A2(G159), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n345), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n300), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n345), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n340), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n341), .B1(new_n267), .B2(G20), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n343), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n226), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n359), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  AND4_X1   g0169(.A1(new_n340), .A2(new_n369), .A3(new_n247), .A4(new_n361), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n326), .B(new_n339), .C1(new_n362), .C2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT17), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n326), .B1(new_n362), .B2(new_n370), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n319), .B1(new_n334), .B2(new_n335), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n334), .A2(new_n335), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n291), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(KEYINPUT18), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n366), .A2(new_n367), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(G68), .B1(new_n350), .B2(new_n356), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n247), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n382));
  INV_X1    g0182(.A(new_n361), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT75), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n369), .A2(new_n340), .A3(new_n361), .A4(new_n247), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n325), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n379), .B1(new_n386), .B2(new_n376), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n378), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n372), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G41), .ZN(new_n391));
  OAI211_X1 g0191(.A(G1), .B(G13), .C1(new_n253), .C2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(G238), .A3(new_n276), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n279), .A2(G274), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT72), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n328), .A2(new_n330), .A3(G232), .A4(G1698), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n328), .A2(new_n330), .A3(G226), .A4(new_n268), .ZN(new_n401));
  INV_X1    g0201(.A(G97), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n400), .B(new_n401), .C1(new_n253), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT71), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(new_n274), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n403), .B2(new_n274), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT13), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT13), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n399), .B(new_n409), .C1(new_n405), .C2(new_n406), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(G190), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n296), .A2(new_n226), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT12), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n226), .A2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(G50), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n414), .B1(new_n251), .B2(new_n203), .C1(new_n415), .C2(new_n254), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(KEYINPUT11), .A3(new_n247), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n413), .B(new_n417), .C1(new_n226), .C2(new_n298), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT11), .B1(new_n416), .B2(new_n247), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G200), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n408), .B2(new_n410), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n403), .A2(new_n274), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT71), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n403), .A2(new_n404), .A3(new_n274), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n409), .B1(new_n428), .B2(new_n399), .ZN(new_n429));
  INV_X1    g0229(.A(new_n410), .ZN(new_n430));
  OAI21_X1  g0230(.A(G169), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n319), .B1(new_n408), .B2(new_n410), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n408), .A2(G179), .A3(new_n410), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n420), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n424), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n439), .A2(KEYINPUT73), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(KEYINPUT73), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n323), .B(new_n390), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT79), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n391), .A2(KEYINPUT5), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n257), .A2(G45), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G41), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(KEYINPUT79), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n277), .B1(KEYINPUT5), .B2(new_n391), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n447), .A2(new_n452), .A3(new_n453), .A4(new_n392), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n391), .A2(KEYINPUT5), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n449), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(G264), .A3(new_n392), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n267), .A2(G250), .A3(new_n268), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n267), .A2(G257), .A3(G1698), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G294), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n274), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n319), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(G179), .B2(new_n464), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n328), .A2(new_n330), .A3(new_n223), .A4(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT22), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n267), .A2(new_n469), .A3(new_n223), .A4(G87), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G116), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT23), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n223), .B2(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n311), .A2(KEYINPUT23), .A3(G20), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n472), .B1(new_n471), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n247), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT84), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(new_n247), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n258), .A2(G107), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT25), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n487), .A2(KEYINPUT85), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(KEYINPUT85), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(KEYINPUT25), .C2(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n257), .A2(G33), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n300), .A2(new_n258), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G107), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n466), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n258), .A2(G116), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G116), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n246), .A2(new_n222), .B1(G20), .B2(new_n500), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n223), .C1(G33), .C2(new_n402), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(KEYINPUT20), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT83), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(new_n504), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n505), .A2(new_n506), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT79), .B1(new_n449), .B2(new_n451), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n455), .B(G274), .C1(new_n273), .C2(new_n222), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n456), .A2(G270), .A3(new_n392), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n517), .A2(new_n452), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n328), .A2(new_n330), .A3(G257), .A4(new_n268), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n328), .A2(new_n330), .A3(G264), .A4(G1698), .ZN(new_n522));
  INV_X1    g0322(.A(G303), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n267), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n274), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n456), .A2(KEYINPUT82), .A3(G270), .A4(new_n392), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n514), .A2(KEYINPUT21), .A3(G169), .A4(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT21), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(G169), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n513), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n520), .A2(G179), .A3(new_n525), .A4(new_n526), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n513), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n497), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n527), .A2(new_n283), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n527), .A2(G200), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n536), .A2(new_n513), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n495), .B1(new_n482), .B2(new_n484), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n464), .A2(new_n283), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(G200), .B2(new_n464), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n446), .A2(G250), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n274), .A2(new_n543), .B1(new_n277), .B2(new_n446), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n328), .A2(new_n330), .A3(G238), .A4(new_n268), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n328), .A2(new_n330), .A3(G244), .A4(G1698), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n473), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n547), .B2(new_n274), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n291), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n319), .B2(new_n548), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n267), .A2(new_n223), .A3(G68), .ZN(new_n551));
  NAND3_X1  g0351(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n223), .ZN(new_n553));
  INV_X1    g0353(.A(G87), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n402), .A3(new_n311), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n251), .B2(new_n402), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n551), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n303), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n559), .A2(new_n247), .B1(new_n296), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n492), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n550), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n328), .A2(new_n330), .A3(G244), .A4(new_n268), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n328), .A2(new_n330), .A3(G250), .A4(G1698), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT78), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n267), .A2(KEYINPUT78), .A3(G250), .A4(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n503), .B1(new_n564), .B2(new_n565), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n274), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n291), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n456), .A2(G257), .A3(new_n392), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n573), .A2(new_n454), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n454), .A3(new_n575), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n319), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n311), .B1(new_n366), .B2(new_n367), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n402), .A2(new_n311), .A3(KEYINPUT6), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT6), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G97), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n311), .A2(KEYINPUT76), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT76), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G107), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n580), .A2(new_n582), .B1(new_n583), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g0387(.A(G20), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n254), .A2(new_n203), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT77), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n579), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n588), .A2(KEYINPUT77), .A3(new_n590), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n300), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n296), .A2(new_n402), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n492), .B2(new_n402), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n576), .B(new_n578), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT81), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n547), .A2(new_n274), .ZN(new_n600));
  INV_X1    g0400(.A(new_n544), .ZN(new_n601));
  AND4_X1   g0401(.A1(KEYINPUT80), .A2(new_n600), .A3(G190), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT80), .B1(new_n548), .B2(G190), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n600), .A2(G190), .A3(new_n601), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT80), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n548), .A2(KEYINPUT80), .A3(G190), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(KEYINPUT81), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n493), .A2(G87), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n561), .B(new_n610), .C1(new_n422), .C2(new_n548), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n604), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n581), .A2(G97), .A3(G107), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n402), .A2(KEYINPUT6), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n584), .A2(G107), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n311), .A2(KEYINPUT76), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n614), .A2(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n223), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n592), .B1(new_n620), .B2(new_n589), .ZN(new_n621));
  INV_X1    g0421(.A(new_n579), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n594), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n597), .B1(new_n623), .B2(new_n247), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n573), .A2(G190), .A3(new_n454), .A4(new_n575), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n577), .A2(G200), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n563), .A2(new_n598), .A3(new_n613), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n443), .A2(new_n535), .A3(new_n542), .A4(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n295), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n290), .A2(new_n287), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT90), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n290), .A2(KEYINPUT90), .A3(new_n287), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n437), .A2(new_n438), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n424), .B2(new_n321), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n372), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT89), .B1(new_n378), .B2(new_n387), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n378), .A2(new_n387), .A3(KEYINPUT89), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n631), .B1(new_n636), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n623), .A2(new_n247), .ZN(new_n644));
  INV_X1    g0444(.A(new_n597), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(new_n319), .B2(new_n577), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(new_n613), .A3(new_n563), .A4(new_n576), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT88), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT86), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n548), .A2(new_n319), .ZN(new_n651));
  AOI211_X1 g0451(.A(new_n574), .B(new_n544), .C1(new_n274), .C2(new_n547), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n549), .B(KEYINPUT86), .C1(new_n319), .C2(new_n548), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n562), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT87), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n611), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n548), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G200), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(KEYINPUT87), .A3(new_n561), .A4(new_n610), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n607), .A2(new_n608), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n648), .B1(new_n664), .B2(new_n598), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n611), .B1(new_n662), .B2(new_n599), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n666), .A2(new_n609), .B1(new_n550), .B2(new_n562), .ZN(new_n667));
  INV_X1    g0467(.A(new_n578), .ZN(new_n668));
  INV_X1    g0468(.A(new_n576), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n668), .A2(new_n624), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n667), .A2(new_n670), .A3(new_n671), .A4(KEYINPUT26), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n649), .A2(new_n665), .A3(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n598), .B(new_n627), .C1(new_n497), .C2(new_n534), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n656), .A2(new_n663), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n539), .A2(new_n541), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n656), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n643), .B1(new_n442), .B2(new_n679), .ZN(G369));
  NAND2_X1  g0480(.A1(new_n485), .A2(new_n496), .ZN(new_n681));
  INV_X1    g0481(.A(new_n466), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G13), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G20), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n257), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n691), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n676), .B1(new_n539), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n691), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n514), .A3(new_n691), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n534), .A2(new_n538), .B1(new_n513), .B2(new_n693), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT91), .Z(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n695), .A2(new_n697), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n692), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n219), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  NOR4_X1   g0510(.A1(new_n710), .A2(new_n257), .A3(G116), .A4(new_n555), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n229), .B2(new_n710), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT28), .Z(new_n713));
  AOI21_X1  g0513(.A(new_n648), .B1(new_n675), .B2(new_n670), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n693), .B1(new_n716), .B2(new_n678), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n718));
  INV_X1    g0518(.A(new_n656), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n598), .A2(new_n627), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n683), .B2(new_n696), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n664), .B1(new_n539), .B2(new_n541), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n649), .A2(new_n665), .A3(new_n672), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n691), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n718), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n291), .B1(new_n458), .B2(new_n463), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n577), .A2(new_n527), .A3(new_n659), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n573), .A2(new_n575), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n458), .A2(new_n463), .A3(new_n548), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n731), .A2(new_n532), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n730), .B1(new_n733), .B2(KEYINPUT30), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n731), .A2(new_n532), .A3(new_n732), .A4(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT31), .B(new_n691), .C1(new_n734), .C2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n691), .B1(new_n734), .B2(new_n736), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n628), .A2(new_n535), .A3(new_n542), .A4(new_n693), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n738), .A3(new_n741), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n746), .A2(G330), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n728), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n713), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n222), .B1(G20), .B2(new_n319), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n709), .A2(new_n267), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT94), .Z(new_n757));
  NAND2_X1  g0557(.A1(new_n229), .A2(new_n448), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n758), .C1(new_n448), .C2(new_n241), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n709), .A2(new_n343), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n760), .A2(G355), .B1(new_n500), .B2(new_n709), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n755), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n753), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n223), .A2(G179), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G329), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n422), .A2(G190), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n764), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n343), .B1(new_n766), .B2(new_n767), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n283), .A2(new_n422), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n764), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n574), .A2(new_n223), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n772), .ZN(new_n778));
  INV_X1    g0578(.A(G326), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n776), .A2(new_n523), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n283), .A2(G179), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n223), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n771), .B(new_n780), .C1(G294), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n777), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n785), .A2(new_n283), .A3(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n777), .A2(new_n769), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n786), .A2(G322), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n777), .A2(new_n765), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n784), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n776), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G87), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n795), .B1(new_n226), .B2(new_n787), .C1(new_n203), .C2(new_n792), .ZN(new_n796));
  INV_X1    g0596(.A(new_n786), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n797), .A2(new_n225), .B1(new_n415), .B2(new_n778), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n267), .B1(new_n770), .B2(new_n311), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT95), .B(G159), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n766), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT32), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n804), .B1(new_n803), .B2(new_n802), .C1(new_n402), .C2(new_n782), .ZN(new_n805));
  OR3_X1    g0605(.A1(new_n796), .A2(new_n798), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n763), .B1(new_n793), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n710), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n257), .B1(new_n685), .B2(G45), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT93), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n762), .A2(new_n807), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n752), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n701), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n702), .A2(new_n812), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n701), .A2(G330), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT97), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n307), .A2(new_n691), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n322), .A2(KEYINPUT99), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n318), .A2(new_n321), .A3(new_n820), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT99), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n693), .B(new_n825), .C1(new_n673), .C2(new_n678), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n321), .A2(new_n693), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n821), .A2(new_n827), .A3(new_n824), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n725), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n747), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n811), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  INV_X1    g0632(.A(new_n792), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G150), .A2(new_n788), .B1(new_n833), .B2(new_n800), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n778), .C1(new_n836), .C2(new_n797), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  INV_X1    g0638(.A(new_n766), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n343), .B1(new_n839), .B2(G132), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n226), .B2(new_n770), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G58), .B2(new_n783), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n838), .B(new_n842), .C1(new_n415), .C2(new_n776), .ZN(new_n843));
  INV_X1    g0643(.A(G294), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n797), .A2(new_n844), .B1(new_n500), .B2(new_n792), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G283), .B2(new_n788), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n343), .B1(new_n766), .B2(new_n791), .C1(new_n554), .C2(new_n770), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G97), .B2(new_n783), .ZN(new_n848));
  INV_X1    g0648(.A(new_n778), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n794), .A2(G107), .B1(new_n849), .B2(G303), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n763), .B1(new_n843), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n753), .A2(new_n750), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT98), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n812), .B(new_n852), .C1(new_n203), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n751), .B2(new_n828), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n832), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G384));
  NAND2_X1  g0659(.A1(new_n346), .A2(G77), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n228), .A2(new_n860), .B1(G50), .B2(new_n226), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(G1), .A3(new_n684), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n586), .A2(new_n587), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(G116), .B(new_n224), .C1(new_n864), .C2(KEYINPUT35), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT100), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n865), .A2(new_n866), .B1(KEYINPUT35), .B2(new_n864), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  XNOR2_X1  g0668(.A(KEYINPUT101), .B(KEYINPUT36), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n744), .A2(new_n742), .A3(new_n737), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT103), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n360), .A2(new_n361), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n326), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n377), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n371), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n689), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n874), .B1(new_n371), .B2(new_n877), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n386), .A2(new_n376), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT37), .B1(new_n884), .B2(KEYINPUT104), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n371), .B1(new_n386), .B2(new_n689), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT104), .B1(new_n373), .B2(new_n377), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n885), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n880), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n389), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n372), .B1(new_n641), .B2(new_n640), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n386), .A2(new_n689), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n886), .B2(new_n884), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n895), .A2(new_n896), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n898), .B2(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n872), .A2(new_n828), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n436), .B1(new_n433), .B2(new_n434), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n431), .A2(KEYINPUT14), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n438), .B(new_n691), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT102), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n437), .A2(KEYINPUT102), .A3(new_n438), .A4(new_n691), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n438), .A2(new_n691), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n905), .A2(new_n906), .B1(new_n439), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n873), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n439), .A2(new_n907), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n913), .A2(new_n873), .A3(new_n828), .A4(new_n872), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n325), .B(new_n338), .C1(new_n384), .C2(new_n385), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n376), .B1(new_n326), .B2(new_n875), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT103), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n880), .A3(new_n878), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n886), .A2(new_n888), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n919), .A2(KEYINPUT37), .B1(new_n920), .B2(new_n885), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n880), .B1(new_n372), .B2(new_n388), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n914), .B1(new_n894), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n443), .B(new_n872), .C1(new_n910), .C2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(G330), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n899), .A2(new_n909), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT40), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n923), .A2(new_n894), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n873), .A3(new_n909), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n926), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n872), .A2(G330), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n442), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n925), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n728), .A2(new_n443), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n643), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n921), .A2(new_n915), .A3(new_n922), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n891), .B2(new_n893), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT39), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT39), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n941), .B(new_n894), .C1(new_n898), .C2(KEYINPUT38), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n437), .A2(new_n438), .A3(new_n693), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n321), .A2(new_n691), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n908), .B1(new_n826), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n929), .A2(new_n949), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n641), .A2(new_n640), .A3(new_n879), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n937), .A2(new_n953), .B1(new_n257), .B2(new_n685), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n937), .A2(new_n953), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n871), .B1(new_n954), .B2(new_n955), .ZN(G367));
  NAND2_X1  g0756(.A1(new_n561), .A2(new_n610), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n691), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n656), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n675), .A2(new_n958), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(KEYINPUT105), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT105), .B2(new_n960), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(new_n814), .ZN(new_n963));
  INV_X1    g0763(.A(new_n757), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n754), .B1(new_n219), .B2(new_n560), .C1(new_n964), .C2(new_n237), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n811), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n786), .A2(G150), .B1(new_n794), .B2(G58), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G50), .A2(new_n833), .B1(new_n849), .B2(G143), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n788), .A2(new_n800), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n267), .B1(new_n766), .B2(new_n835), .C1(new_n203), .C2(new_n770), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G68), .B2(new_n783), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n786), .A2(G303), .B1(G311), .B2(new_n849), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n343), .B1(new_n766), .B2(new_n974), .C1(new_n402), .C2(new_n770), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G107), .B2(new_n783), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G283), .A2(new_n833), .B1(new_n788), .B2(G294), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n776), .A2(new_n500), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT46), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n972), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT108), .Z(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT47), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n763), .B1(new_n982), .B2(KEYINPUT47), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n966), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n963), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n809), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n624), .A2(new_n693), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n720), .A2(new_n988), .B1(new_n598), .B2(new_n693), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n707), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT45), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n707), .A2(new_n989), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n705), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n991), .A2(new_n704), .A3(new_n993), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n706), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n703), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n702), .B2(new_n698), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n748), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n748), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n710), .B(KEYINPUT41), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n987), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n706), .A2(new_n721), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT42), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n989), .B(KEYINPUT107), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n497), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n691), .B1(new_n1012), .B2(new_n598), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1007), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT106), .Z(new_n1016));
  XNOR2_X1  g0816(.A(new_n1014), .B(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n705), .A2(new_n1010), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1017), .B(new_n1018), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n986), .B1(new_n1006), .B2(new_n1020), .ZN(G387));
  NOR2_X1   g0821(.A1(new_n1002), .A2(new_n808), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n748), .B2(new_n1000), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1000), .A2(new_n987), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n757), .B1(new_n448), .B2(new_n234), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n555), .A2(G116), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n760), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n250), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT50), .B1(new_n250), .B2(G50), .ZN(new_n1030));
  AOI21_X1  g0830(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1029), .A2(new_n1026), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1028), .A2(new_n1032), .B1(new_n311), .B2(new_n709), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n811), .B1(new_n1033), .B2(new_n755), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n778), .A2(new_n348), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT109), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n267), .B1(new_n766), .B2(new_n252), .C1(new_n402), .C2(new_n770), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n303), .B2(new_n783), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G68), .A2(new_n833), .B1(new_n788), .B2(new_n249), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n786), .A2(G50), .B1(new_n794), .B2(G77), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n267), .B1(new_n839), .B2(G326), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G303), .A2(new_n833), .B1(new_n788), .B2(G311), .ZN(new_n1043));
  INV_X1    g0843(.A(G322), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n778), .C1(new_n974), .C2(new_n797), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT48), .Z(new_n1046));
  OAI22_X1  g0846(.A1(new_n776), .A2(new_n844), .B1(new_n768), .B2(new_n782), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1042), .B1(new_n500), .B2(new_n770), .C1(new_n1048), .C2(KEYINPUT49), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1048), .A2(KEYINPUT49), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1041), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1034), .B1(new_n1051), .B2(new_n753), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n695), .B2(new_n814), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1023), .A2(new_n1024), .A3(new_n1053), .ZN(G393));
  NAND2_X1  g0854(.A1(new_n997), .A2(new_n987), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n757), .A2(new_n244), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n754), .C1(new_n402), .C2(new_n219), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n267), .B1(new_n766), .B2(new_n836), .C1(new_n554), .C2(new_n770), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n794), .A2(G68), .B1(new_n788), .B2(G50), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n250), .B2(new_n792), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(G77), .C2(new_n783), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n786), .A2(G159), .B1(G150), .B2(new_n849), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT51), .Z(new_n1063));
  OAI221_X1 g0863(.A(new_n343), .B1(new_n766), .B2(new_n1044), .C1(new_n311), .C2(new_n770), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G294), .A2(new_n833), .B1(new_n788), .B2(G303), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n768), .B2(new_n776), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(G116), .C2(new_n783), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n786), .A2(G311), .B1(G317), .B2(new_n849), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n1061), .A2(new_n1063), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n811), .B(new_n1057), .C1(new_n1070), .C2(new_n763), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT110), .Z(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1011), .B2(new_n814), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1055), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n995), .A2(new_n1001), .A3(new_n996), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1003), .A2(new_n710), .A3(new_n1075), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT111), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(KEYINPUT111), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G390));
  INV_X1    g0880(.A(new_n643), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n442), .B1(new_n718), .B2(new_n727), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1081), .A2(new_n1082), .A3(new_n933), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n947), .B1(new_n725), .B2(new_n825), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n746), .A2(G330), .A3(new_n828), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n908), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1086), .A2(KEYINPUT113), .B1(new_n909), .B2(G330), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT113), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1088), .A3(new_n908), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1084), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n747), .A2(new_n828), .A3(new_n913), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n714), .A2(new_n715), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n691), .B1(new_n723), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n947), .B1(new_n1093), .B2(new_n825), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n908), .B1(new_n900), .B2(new_n926), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1083), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n944), .B1(new_n1084), .B2(new_n908), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n940), .A3(new_n942), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n944), .B(KEYINPUT112), .Z(new_n1100));
  OAI211_X1 g0900(.A(new_n899), .B(new_n1100), .C1(new_n908), .C2(new_n1094), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1099), .A2(new_n1101), .A3(new_n1091), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n909), .A2(G330), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1097), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n442), .A2(new_n932), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n935), .A2(new_n643), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1086), .A2(KEYINPUT113), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n1103), .A3(new_n1089), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1084), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1096), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1103), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1099), .A2(new_n1101), .A3(new_n1091), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1113), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1105), .A2(new_n1118), .A3(new_n710), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n940), .A2(new_n942), .A3(new_n750), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n811), .B1(new_n249), .B2(new_n854), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n770), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G68), .A2(new_n1123), .B1(new_n839), .B2(G294), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n203), .B2(new_n782), .C1(new_n797), .C2(new_n500), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n778), .A2(new_n768), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n402), .A2(new_n792), .B1(new_n787), .B2(new_n311), .ZN(new_n1127));
  OR3_X1    g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n795), .A2(new_n343), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT114), .Z(new_n1130));
  NAND2_X1  g0930(.A1(new_n794), .A2(G150), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n786), .A2(G132), .B1(G128), .B2(new_n849), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n343), .B1(new_n839), .B2(G125), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n415), .B2(new_n770), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G159), .B2(new_n783), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT54), .B(G143), .Z(new_n1137));
  AOI22_X1  g0937(.A1(G137), .A2(new_n788), .B1(new_n833), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1128), .A2(new_n1130), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1122), .B1(new_n1140), .B2(new_n753), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1120), .A2(new_n987), .B1(new_n1121), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1119), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT115), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1119), .A2(new_n1142), .A3(KEYINPUT115), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(G378));
  NAND2_X1  g0947(.A1(new_n1118), .A2(new_n1083), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n634), .A2(new_n295), .A3(new_n635), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n263), .A2(new_n689), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1154), .B1(new_n1157), .B2(new_n1151), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT117), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n931), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(G330), .C1(new_n910), .C2(new_n924), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n944), .B1(new_n940), .B2(new_n942), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n950), .A2(new_n951), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1161), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n931), .A2(new_n953), .A3(new_n1160), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1170));
  OAI21_X1  g0970(.A(G330), .B1(new_n910), .B2(new_n924), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(KEYINPUT117), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1169), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1148), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1148), .A2(new_n1168), .A3(new_n1174), .A4(KEYINPUT57), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n710), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1168), .A2(new_n1174), .A3(new_n987), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n811), .B1(G50), .B2(new_n854), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n786), .A2(G107), .B1(G97), .B2(new_n788), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n560), .B2(new_n792), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1123), .A2(G58), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n267), .A2(G41), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n226), .B2(new_n782), .C1(new_n768), .C2(new_n766), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n776), .A2(new_n203), .B1(new_n778), .B2(new_n500), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1183), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT58), .Z(new_n1190));
  NOR2_X1   g0990(.A1(G33), .A2(G41), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT116), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1185), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n415), .B2(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n786), .A2(G128), .B1(G137), .B2(new_n833), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n794), .A2(new_n1137), .B1(new_n849), .B2(G125), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n788), .A2(G132), .B1(G150), .B2(new_n783), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  INV_X1    g1000(.A(G124), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n801), .A2(new_n770), .B1(new_n766), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1199), .B2(KEYINPUT59), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1192), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1190), .B1(new_n1195), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1181), .B1(new_n1205), .B2(new_n753), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1159), .B2(new_n751), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1180), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1179), .A2(new_n1208), .ZN(G375));
  AOI21_X1  g1009(.A(new_n812), .B1(new_n226), .B2(new_n855), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n839), .A2(G128), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1184), .A2(new_n1211), .A3(new_n267), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G150), .A2(new_n833), .B1(new_n788), .B2(new_n1137), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n348), .B2(new_n776), .C1(new_n835), .C2(new_n797), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1212), .B(new_n1214), .C1(G50), .C2(new_n783), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n849), .A2(G132), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT121), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n797), .A2(new_n768), .B1(new_n402), .B2(new_n776), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n343), .B1(new_n770), .B2(new_n203), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT120), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n783), .A2(new_n303), .B1(new_n839), .B2(G303), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n778), .B2(new_n844), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1218), .A2(new_n1220), .A3(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n311), .A2(new_n792), .B1(new_n787), .B2(new_n500), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT119), .Z(new_n1225));
  AOI22_X1  g1025(.A1(new_n1215), .A2(new_n1217), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1210), .B1(new_n763), .B2(new_n1226), .C1(new_n913), .C2(new_n751), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1096), .B1(new_n1110), .B2(new_n1109), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n809), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(KEYINPUT118), .A3(new_n1107), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT118), .B1(new_n1228), .B2(new_n1107), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1097), .A2(new_n1005), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1230), .B1(new_n1234), .B2(new_n1235), .ZN(G381));
  NAND2_X1  g1036(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n809), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1238), .A2(new_n1019), .B1(new_n963), .B2(new_n985), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1079), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G375), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1143), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OR3_X1    g1044(.A1(new_n1241), .A2(G381), .A3(new_n1244), .ZN(G407));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G343), .C2(new_n1244), .ZN(G409));
  XOR2_X1   g1046(.A(G393), .B(G396), .Z(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G387), .B2(KEYINPUT125), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G387), .A2(new_n1247), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(G390), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1250), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1079), .B1(new_n1252), .B2(new_n1248), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G213), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(G343), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1179), .A2(G378), .A3(new_n1208), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1005), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1180), .B(new_n1207), .C1(new_n1175), .C2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1243), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1256), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1097), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1111), .A2(new_n1112), .A3(new_n1107), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n710), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1264), .A2(KEYINPUT123), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT118), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1265), .A2(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1272), .A2(new_n1231), .B1(new_n1097), .B2(new_n1262), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1270), .B1(new_n1273), .B2(new_n1267), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1269), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G384), .B1(new_n1275), .B2(new_n1230), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n858), .B(new_n1229), .C1(new_n1269), .C2(new_n1274), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1261), .A2(KEYINPUT63), .A3(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1254), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1256), .A2(G2897), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1261), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT124), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1256), .ZN(new_n1288));
  AND4_X1   g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1278), .A4(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1261), .B2(new_n1278), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1285), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1280), .A2(new_n1281), .A3(new_n1284), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1284), .A2(new_n1281), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1261), .A2(KEYINPUT62), .A3(new_n1278), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1294), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(KEYINPUT126), .B(new_n1295), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1293), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1292), .B1(new_n1300), .B2(new_n1254), .ZN(G405));
  NOR2_X1   g1101(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1254), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1254), .A2(new_n1302), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1257), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1243), .B2(G375), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1303), .A2(new_n1308), .A3(new_n1307), .A4(new_n1304), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(G402));
endmodule


