//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  AOI211_X1 g0002(.A(G50), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT66), .Z(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT67), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(KEYINPUT67), .B1(new_n211), .B2(new_n212), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n207), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n201), .A2(new_n202), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n210), .A2(new_n219), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT68), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT71), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G232), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G107), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n253), .B(new_n254), .C1(new_n255), .C2(new_n251), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n248), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n261), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n262), .B1(G244), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n258), .A2(new_n271), .A3(new_n267), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT70), .ZN(new_n274));
  INV_X1    g0074(.A(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT8), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT8), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n279), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT15), .B(G87), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n224), .A2(G33), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n223), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n274), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n286), .A2(new_n274), .A3(new_n288), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n288), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n260), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n295), .A2(new_n297), .B1(new_n296), .B2(new_n294), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n273), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n286), .A2(new_n274), .A3(new_n288), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n300), .B2(new_n289), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n268), .A2(G200), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n258), .A2(G190), .A3(new_n267), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n246), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n251), .A2(G222), .A3(new_n252), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n251), .A2(G223), .A3(G1698), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n307), .B(new_n308), .C1(new_n296), .C2(new_n251), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n257), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n262), .B1(G226), .B2(new_n266), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(G179), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n224), .B1(new_n220), .B2(new_n221), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n280), .A2(G150), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n285), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n288), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n221), .B1(new_n260), .B2(G20), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n295), .A2(new_n321), .B1(new_n221), .B2(new_n294), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n313), .A2(new_n315), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n320), .A2(new_n322), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n312), .A2(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n323), .A2(KEYINPUT9), .B1(new_n314), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT10), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n312), .A2(G190), .B1(new_n326), .B2(new_n327), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n323), .A2(KEYINPUT9), .B1(new_n314), .B2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT10), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n324), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n292), .A2(new_n298), .A3(new_n303), .A4(new_n302), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n270), .A2(new_n272), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n301), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT71), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n306), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G58), .A2(G68), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n201), .A2(new_n202), .A3(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT76), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n249), .A2(new_n224), .A3(new_n250), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT7), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n224), .A4(new_n250), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n345), .B1(new_n350), .B2(G68), .ZN(new_n351));
  INV_X1    g0151(.A(G68), .ZN(new_n352));
  AOI211_X1 g0152(.A(KEYINPUT76), .B(new_n352), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  OAI211_X1 g0153(.A(KEYINPUT16), .B(new_n344), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n287), .A2(new_n223), .ZN(new_n355));
  AND2_X1   g0155(.A1(KEYINPUT3), .A2(G33), .ZN(new_n356));
  NOR2_X1   g0156(.A1(KEYINPUT3), .A2(G33), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT7), .B1(new_n358), .B2(new_n224), .ZN(new_n359));
  INV_X1    g0159(.A(new_n349), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n344), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n355), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n354), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT78), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n355), .A2(new_n293), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n260), .A2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n279), .A2(new_n368), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n367), .A2(new_n369), .B1(new_n293), .B2(new_n279), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT77), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n252), .A2(G226), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n251), .B(new_n374), .C1(G223), .C2(G1698), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n264), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n264), .A2(G274), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n230), .A2(new_n265), .B1(new_n378), .B2(new_n261), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n325), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n375), .A2(new_n376), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n257), .ZN(new_n382));
  INV_X1    g0182(.A(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n380), .B1(new_n384), .B2(G190), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n365), .A2(new_n366), .A3(new_n373), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n365), .A2(new_n373), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n377), .A2(new_n379), .A3(new_n271), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(G169), .B2(new_n384), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n372), .B1(new_n354), .B2(new_n364), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT18), .B1(new_n395), .B2(new_n392), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n366), .A3(KEYINPUT17), .A4(new_n385), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n388), .A2(new_n394), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n341), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G97), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(G226), .B(new_n252), .C1(new_n356), .C2(new_n357), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT72), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT72), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n251), .A2(new_n405), .A3(G226), .A4(new_n252), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n264), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n262), .B1(G238), .B2(new_n266), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT13), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT13), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n400), .A2(new_n401), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n406), .B2(new_n404), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n412), .B(new_n409), .C1(new_n414), .C2(new_n264), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(new_n415), .A3(G190), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT73), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT73), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n411), .A2(new_n415), .A3(new_n418), .A4(G190), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n224), .A2(G33), .A3(G77), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n352), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n355), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g0223(.A(new_n423), .B(KEYINPUT11), .Z(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT74), .B1(new_n293), .B2(G68), .ZN(new_n425));
  XOR2_X1   g0225(.A(new_n425), .B(KEYINPUT12), .Z(new_n426));
  NAND3_X1  g0226(.A1(new_n295), .A2(G68), .A3(new_n368), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n411), .A2(new_n415), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(G200), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n420), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n411), .A2(new_n415), .A3(G179), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n411), .A2(new_n415), .A3(KEYINPUT75), .A4(G179), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n429), .A2(G169), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT14), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n429), .A2(new_n439), .A3(G169), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n431), .B1(new_n428), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n399), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n260), .A2(G45), .ZN(new_n445));
  OR2_X1    g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  NAND2_X1  g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(new_n257), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n257), .A2(new_n259), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n449), .A2(G270), .B1(new_n450), .B2(new_n448), .ZN(new_n451));
  OAI211_X1 g0251(.A(G264), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n452));
  OAI211_X1 g0252(.A(G257), .B(new_n252), .C1(new_n356), .C2(new_n357), .ZN(new_n453));
  XOR2_X1   g0253(.A(KEYINPUT81), .B(G303), .Z(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(new_n251), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n257), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(G179), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n287), .A2(new_n223), .B1(G20), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n224), .C1(G33), .C2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n459), .A2(KEYINPUT20), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT20), .B1(new_n459), .B2(new_n462), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n294), .A2(new_n458), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n260), .A2(G33), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n355), .A2(new_n293), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(new_n458), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n457), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT82), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n269), .B1(new_n451), .B2(new_n456), .ZN(new_n473));
  OAI221_X1 g0273(.A(new_n466), .B1(new_n468), .B2(new_n458), .C1(new_n463), .C2(new_n464), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n451), .A2(new_n456), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(new_n474), .A3(G169), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT21), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n474), .B1(new_n478), .B2(G200), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n329), .B2(new_n478), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n477), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT83), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT4), .A2(G244), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n252), .B(new_n486), .C1(new_n356), .C2(new_n357), .ZN(new_n487));
  INV_X1    g0287(.A(G244), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n249), .B2(new_n250), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n460), .C1(new_n489), .C2(KEYINPUT4), .ZN(new_n490));
  OAI21_X1  g0290(.A(G250), .B1(new_n356), .B2(new_n357), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n252), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n257), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n449), .A2(G257), .B1(new_n450), .B2(new_n448), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n493), .A2(KEYINPUT79), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT79), .B1(new_n493), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n269), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n493), .A2(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n280), .A2(G77), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n500), .A2(new_n461), .A3(G107), .ZN(new_n501));
  XNOR2_X1  g0301(.A(G97), .B(G107), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n499), .B1(new_n503), .B2(new_n224), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n255), .B1(new_n348), .B2(new_n349), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n288), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  MUX2_X1   g0306(.A(new_n293), .B(new_n468), .S(G97), .Z(new_n507));
  AOI22_X1  g0307(.A1(new_n498), .A2(new_n271), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n497), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n493), .A2(new_n494), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n493), .A2(KEYINPUT79), .A3(new_n494), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(G190), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n506), .A2(new_n507), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n325), .B1(new_n493), .B2(new_n494), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G45), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G1), .ZN(new_n520));
  INV_X1    g0320(.A(new_n447), .ZN(new_n521));
  NOR2_X1   g0321(.A1(KEYINPUT5), .A2(G41), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G264), .A3(new_n264), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT85), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n523), .A2(new_n526), .A3(G264), .A4(new_n264), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n450), .A2(new_n448), .ZN(new_n529));
  OAI211_X1 g0329(.A(G257), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G250), .B(new_n252), .C1(new_n356), .C2(new_n357), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT84), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n251), .A2(KEYINPUT84), .A3(G250), .A4(new_n252), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n528), .B(new_n529), .C1(new_n264), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n257), .B1(new_n540), .B2(new_n532), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n541), .A2(G190), .A3(new_n529), .A4(new_n528), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n224), .B(G87), .C1(new_n356), .C2(new_n357), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT22), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n251), .A2(new_n545), .A3(new_n224), .A4(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(G20), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT23), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n224), .B2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n255), .A2(KEYINPUT23), .A3(G20), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n547), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n548), .B1(new_n547), .B2(new_n554), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n288), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT25), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n293), .B2(G107), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n293), .A2(new_n559), .A3(G107), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n255), .A2(new_n468), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n539), .A2(new_n542), .A3(new_n558), .A4(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G244), .B(G1698), .C1(new_n356), .C2(new_n357), .ZN(new_n566));
  OAI211_X1 g0366(.A(G238), .B(new_n252), .C1(new_n356), .C2(new_n357), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n549), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n257), .ZN(new_n569));
  INV_X1    g0369(.A(G250), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n520), .A2(KEYINPUT80), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(G274), .B1(KEYINPUT80), .B2(G250), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n445), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n264), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(G169), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n569), .A2(new_n574), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(new_n271), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n224), .B1(new_n401), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n461), .A3(new_n255), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n224), .B(G68), .C1(new_n356), .C2(new_n357), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n578), .B1(new_n285), .B2(new_n461), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n288), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n282), .A2(new_n283), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT15), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G87), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n588), .A2(new_n590), .A3(new_n283), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n294), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n586), .B(new_n592), .C1(new_n284), .C2(new_n468), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n325), .B1(new_n569), .B2(new_n574), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n295), .A2(G87), .A3(new_n467), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n586), .A2(new_n595), .A3(new_n592), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n576), .A2(G190), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n577), .A2(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n509), .A2(new_n518), .A3(new_n565), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n538), .A2(new_n269), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n541), .A2(new_n271), .A3(new_n529), .A4(new_n528), .ZN(new_n602));
  INV_X1    g0402(.A(new_n557), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n355), .B1(new_n603), .B2(new_n555), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n601), .B(new_n602), .C1(new_n604), .C2(new_n563), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n444), .A2(new_n485), .A3(new_n607), .ZN(G372));
  NAND2_X1  g0408(.A1(new_n441), .A2(new_n428), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n431), .B2(new_n339), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n388), .A3(new_n397), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n396), .A3(new_n394), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n331), .A2(new_n335), .ZN(new_n613));
  XOR2_X1   g0413(.A(new_n613), .B(KEYINPUT86), .Z(new_n614));
  AOI21_X1  g0414(.A(new_n324), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n569), .A2(new_n574), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n269), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(new_n593), .C1(G179), .C2(new_n616), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n605), .A2(new_n477), .A3(new_n481), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n597), .A2(new_n598), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n497), .A2(new_n508), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  OAI221_X1 g0424(.A(new_n618), .B1(new_n619), .B2(new_n600), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n444), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n615), .A2(new_n626), .ZN(G369));
  NAND3_X1  g0427(.A1(new_n260), .A2(new_n224), .A3(G13), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(G213), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G343), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n470), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT87), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT88), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n485), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n637), .B2(new_n485), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n477), .A2(new_n481), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n636), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G330), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n633), .B1(new_n604), .B2(new_n563), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n606), .B1(new_n565), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n606), .B2(new_n634), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n640), .A2(new_n634), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n605), .B2(new_n633), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n208), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n581), .A2(G116), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G1), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n222), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n657), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT28), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT30), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n541), .A2(new_n576), .A3(new_n528), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n495), .A2(new_n496), .A3(new_n457), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n663), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n664), .B(KEYINPUT89), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(KEYINPUT30), .A3(new_n667), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n576), .A2(G179), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n478), .A3(new_n538), .A4(new_n510), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n674), .A2(KEYINPUT31), .A3(new_n633), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT31), .B1(new_n674), .B2(new_n633), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n485), .A2(new_n607), .A3(new_n634), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n643), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n625), .A2(new_n634), .A3(new_n680), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n625), .A2(new_n634), .B1(KEYINPUT90), .B2(KEYINPUT29), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n662), .B1(new_n684), .B2(G1), .ZN(G364));
  AND2_X1   g0485(.A1(new_n224), .A2(G13), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n260), .B1(new_n686), .B2(G45), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n657), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT91), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(G13), .A2(G33), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G20), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n223), .B1(G20), .B2(new_n269), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n208), .A2(G355), .A3(new_n251), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n655), .A2(new_n251), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(G45), .B2(new_n660), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n244), .A2(G45), .ZN(new_n699));
  OAI221_X1 g0499(.A(new_n696), .B1(G116), .B2(new_n208), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n690), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n694), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n224), .A2(G179), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n329), .A3(G200), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n255), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n358), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(G190), .A3(G200), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G87), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n224), .A2(new_n271), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G200), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n329), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n706), .B(new_n709), .C1(new_n221), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(G190), .A2(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n703), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G159), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT32), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n710), .B(KEYINPUT92), .Z(new_n720));
  NOR3_X1   g0520(.A1(new_n720), .A2(new_n329), .A3(G200), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n719), .B1(new_n722), .B2(new_n275), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n720), .A2(G190), .A3(G200), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n714), .B(new_n723), .C1(G77), .C2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n271), .A2(new_n325), .A3(G190), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G97), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n711), .A2(G190), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n730), .B2(new_n352), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT93), .ZN(new_n732));
  INV_X1    g0532(.A(G326), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n713), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g0534(.A1(KEYINPUT33), .A2(G317), .ZN(new_n735));
  NAND2_X1  g0535(.A1(KEYINPUT33), .A2(G317), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n730), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n734), .B(new_n737), .C1(G294), .C2(new_n727), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n721), .A2(G322), .ZN(new_n739));
  INV_X1    g0539(.A(new_n704), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n251), .B1(new_n740), .B2(G283), .ZN(new_n741));
  INV_X1    g0541(.A(new_n716), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n708), .A2(G303), .B1(new_n742), .B2(G329), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(G311), .B2(new_n724), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n725), .A2(new_n732), .B1(new_n738), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n642), .ZN(new_n747));
  INV_X1    g0547(.A(new_n693), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n701), .B1(new_n702), .B2(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n688), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n644), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n747), .A2(G330), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(G396));
  NOR2_X1   g0554(.A1(new_n694), .A2(new_n691), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n689), .B1(G77), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n721), .A2(G143), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G137), .A2(new_n712), .B1(new_n729), .B2(G150), .ZN(new_n759));
  INV_X1    g0559(.A(new_n724), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(new_n717), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT34), .Z(new_n762));
  NAND2_X1  g0562(.A1(new_n740), .A2(G68), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n221), .B2(new_n707), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n358), .B(new_n764), .C1(G132), .C2(new_n742), .ZN(new_n765));
  INV_X1    g0565(.A(new_n727), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n275), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n712), .A2(G303), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n768), .B(new_n728), .C1(new_n730), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n707), .A2(new_n255), .B1(new_n716), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n251), .B(new_n772), .C1(G87), .C2(new_n740), .ZN(new_n773));
  INV_X1    g0573(.A(G294), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n773), .B1(new_n760), .B2(new_n458), .C1(new_n774), .C2(new_n722), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n762), .A2(new_n767), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n757), .B1(new_n776), .B2(new_n694), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n339), .A2(new_n633), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n301), .A2(new_n633), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n337), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(new_n339), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n777), .B1(new_n692), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n625), .A2(new_n634), .ZN(new_n783));
  INV_X1    g0583(.A(new_n781), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n618), .B1(new_n619), .B2(new_n600), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n621), .B(KEYINPUT26), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n781), .B(new_n634), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT94), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n785), .B(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n679), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n688), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n782), .B1(new_n793), .B2(new_n794), .ZN(G384));
  INV_X1    g0595(.A(new_n503), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT35), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT35), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n797), .A2(G116), .A3(new_n225), .A4(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT36), .Z(new_n800));
  NAND3_X1  g0600(.A1(new_n222), .A2(G77), .A3(new_n342), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n221), .A2(G68), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n260), .B(G13), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n631), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n394), .B2(new_n396), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n778), .B(KEYINPUT95), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n788), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n420), .A2(new_n430), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n428), .A2(new_n633), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n609), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n428), .B(new_n633), .C1(new_n431), .C2(new_n441), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT96), .ZN(new_n815));
  INV_X1    g0615(.A(new_n344), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n361), .A2(KEYINPUT76), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n350), .A2(new_n345), .A3(G68), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n288), .B1(new_n819), .B2(KEYINPUT16), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT97), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n344), .B1(new_n351), .B2(new_n353), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n363), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n824), .A2(KEYINPUT97), .A3(new_n288), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n822), .A2(new_n354), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n370), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n631), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n398), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(KEYINPUT98), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT98), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n398), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n393), .A2(new_n805), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n826), .B2(new_n827), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n395), .A2(new_n385), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT37), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n395), .A2(new_n392), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n389), .A2(KEYINPUT99), .A3(new_n805), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT99), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n395), .B2(new_n631), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n838), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n830), .A2(new_n832), .B1(new_n836), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT100), .B1(new_n845), .B2(KEYINPUT38), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n354), .B1(new_n820), .B2(new_n821), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT97), .B1(new_n824), .B2(new_n288), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n827), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n833), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n835), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n844), .B1(new_n851), .B2(new_n843), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n831), .B1(new_n828), .B2(new_n398), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n828), .A2(new_n398), .A3(new_n831), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT100), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n852), .B(KEYINPUT38), .C1(new_n853), .C2(new_n854), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n846), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n806), .B1(new_n815), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n398), .A2(new_n841), .A3(new_n839), .ZN(new_n863));
  INV_X1    g0663(.A(new_n844), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n843), .B1(new_n838), .B2(new_n842), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n857), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n441), .A2(new_n428), .A3(new_n634), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT101), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n861), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT102), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n683), .A2(new_n875), .A3(new_n444), .ZN(new_n876));
  NAND2_X1  g0676(.A1(KEYINPUT90), .A2(KEYINPUT29), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n783), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n625), .A2(new_n634), .A3(new_n680), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n444), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT102), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(new_n615), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n874), .B(new_n883), .Z(new_n884));
  NAND2_X1  g0684(.A1(new_n674), .A2(new_n633), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT31), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n674), .A2(KEYINPUT31), .A3(new_n633), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n678), .A3(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n889), .A2(new_n781), .A3(new_n813), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n860), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n868), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT40), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n443), .B1(new_n677), .B2(new_n678), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n643), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n897), .B2(new_n896), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n884), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n260), .B2(new_n686), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n884), .A2(new_n899), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n804), .B1(new_n901), .B2(new_n902), .ZN(G367));
  XOR2_X1   g0703(.A(new_n687), .B(KEYINPUT108), .Z(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n684), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT107), .B1(new_n647), .B2(new_n650), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n644), .B(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n908), .A2(new_n651), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n651), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT44), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n515), .A2(new_n633), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n509), .A2(new_n518), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n497), .A2(new_n508), .A3(new_n633), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n912), .B1(new_n653), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n916), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n652), .A2(KEYINPUT44), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n653), .A2(KEYINPUT45), .A3(new_n916), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT45), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n652), .B2(new_n918), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n917), .A2(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n644), .A2(KEYINPUT106), .A3(new_n647), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n923), .B(new_n924), .Z(new_n925));
  AOI21_X1  g0725(.A(new_n906), .B1(new_n911), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n656), .B(new_n927), .Z(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n905), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n651), .A2(new_n918), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT42), .Z(new_n932));
  INV_X1    g0732(.A(new_n518), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n509), .B1(new_n933), .B2(new_n605), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n634), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT104), .ZN(new_n936));
  INV_X1    g0736(.A(new_n618), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n596), .A2(new_n633), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT103), .Z(new_n939));
  MUX2_X1   g0739(.A(new_n599), .B(new_n937), .S(new_n939), .Z(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n935), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n936), .B1(new_n935), .B2(new_n941), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n940), .B(KEYINPUT43), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n942), .A2(new_n943), .B1(new_n935), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n648), .A2(new_n918), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n930), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n697), .ZN(new_n949));
  OAI221_X1 g0749(.A(new_n695), .B1(new_n208), .B2(new_n284), .C1(new_n949), .C2(new_n236), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n689), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(G317), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n358), .B1(new_n716), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n707), .A2(new_n458), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n713), .A2(new_n771), .B1(KEYINPUT46), .B2(new_n954), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n953), .B(new_n955), .C1(G97), .C2(new_n740), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n769), .B2(new_n760), .C1(new_n454), .C2(new_n722), .ZN(new_n957));
  AOI22_X1  g0757(.A1(KEYINPUT46), .A2(new_n954), .B1(new_n729), .B2(G294), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n255), .B2(new_n766), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n766), .A2(new_n352), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n721), .B2(G150), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n724), .A2(G50), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n358), .B1(new_n708), .B2(G58), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n740), .A2(G77), .B1(new_n742), .B2(G137), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G143), .A2(new_n712), .B1(new_n729), .B2(G159), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n957), .A2(new_n959), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT47), .Z(new_n969));
  OAI221_X1 g0769(.A(new_n951), .B1(new_n748), .B2(new_n940), .C1(new_n969), .C2(new_n702), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n948), .A2(new_n970), .ZN(G387));
  OAI21_X1  g0771(.A(new_n695), .B1(new_n208), .B2(new_n255), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n358), .A2(G45), .ZN(new_n973));
  INV_X1    g0773(.A(new_n658), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n318), .A2(G50), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n519), .B1(new_n352), .B2(new_n296), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n975), .B2(new_n976), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n251), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n233), .A2(new_n973), .B1(new_n974), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n972), .B1(new_n981), .B2(new_n208), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n690), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT112), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n724), .A2(G68), .B1(new_n279), .B2(new_n729), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT113), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n251), .B1(new_n704), .B2(new_n461), .ZN(new_n987));
  INV_X1    g0787(.A(G150), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n707), .A2(new_n296), .B1(new_n716), .B2(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(G159), .C2(new_n712), .ZN(new_n990));
  INV_X1    g0790(.A(new_n284), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n727), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n721), .A2(G50), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n986), .A2(new_n990), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n454), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G317), .A2(new_n721), .B1(new_n724), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(G322), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n730), .A2(new_n771), .B1(new_n713), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT48), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n708), .A2(G294), .B1(G283), .B2(new_n727), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(KEYINPUT49), .A3(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n358), .B1(new_n716), .B2(new_n733), .C1(new_n458), .C2(new_n704), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT115), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT49), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n994), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n984), .B1(new_n694), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n647), .B2(new_n748), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT116), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n909), .A2(new_n906), .A3(new_n910), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n656), .B(KEYINPUT117), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n911), .A2(new_n904), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1015), .B(new_n1020), .C1(new_n1022), .C2(new_n1023), .ZN(G393));
  OR2_X1    g0824(.A1(new_n923), .A2(new_n648), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n923), .A2(new_n648), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1017), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1019), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n1016), .B2(new_n925), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT118), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n905), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n1027), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n695), .B1(new_n208), .B2(new_n461), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n241), .B2(new_n697), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n690), .A2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n729), .A2(new_n995), .B1(new_n727), .B2(G116), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n760), .B2(new_n774), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT119), .Z(new_n1040));
  OAI22_X1  g0840(.A1(new_n707), .A2(new_n769), .B1(new_n716), .B2(new_n997), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1040), .A2(new_n251), .A3(new_n705), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n721), .A2(G311), .B1(G317), .B2(new_n712), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  AOI22_X1  g0844(.A1(new_n721), .A2(G159), .B1(G150), .B2(new_n712), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT51), .Z(new_n1046));
  NAND2_X1  g0846(.A1(new_n727), .A2(G77), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n730), .B2(new_n221), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n708), .A2(G68), .B1(new_n742), .B2(G143), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1049), .B(new_n251), .C1(new_n580), .C2(new_n704), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(new_n279), .C2(new_n724), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1042), .A2(new_n1044), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1037), .B1(new_n748), .B2(new_n916), .C1(new_n1052), .C2(new_n702), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1034), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1031), .A2(new_n1054), .ZN(G390));
  NAND2_X1  g0855(.A1(new_n679), .A2(new_n444), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n875), .B1(new_n683), .B2(new_n444), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n681), .A2(new_n682), .A3(new_n443), .A4(KEYINPUT102), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n615), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT122), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n813), .B1(new_n679), .B2(new_n781), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n889), .A2(G330), .A3(new_n781), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n813), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n808), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n679), .A2(new_n781), .A3(new_n813), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n788), .A4(new_n807), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT122), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n882), .A2(new_n1070), .A3(new_n615), .A4(new_n1056), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1060), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1066), .A2(KEYINPUT121), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT121), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1064), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT120), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n814), .B2(new_n873), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n788), .A2(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1078), .A2(KEYINPUT120), .A3(new_n872), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n862), .A2(new_n1080), .A3(new_n869), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n868), .A2(new_n873), .A3(new_n814), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1073), .B(new_n1075), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AND4_X1   g0883(.A1(new_n1074), .A2(new_n1081), .A3(new_n1064), .A4(new_n1082), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1072), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1073), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1075), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1081), .A2(new_n1074), .A3(new_n1064), .A4(new_n1082), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1060), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1085), .A2(new_n1019), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1047), .B1(new_n722), .B2(new_n458), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT124), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n742), .A2(G294), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n709), .A2(new_n763), .A3(new_n358), .A4(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n730), .A2(new_n255), .B1(new_n713), .B2(new_n769), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(G97), .C2(new_n724), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n707), .A2(KEYINPUT53), .A3(new_n988), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT53), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n708), .B2(G150), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1100), .B(new_n1102), .C1(G128), .C2(new_n712), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT123), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n724), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(G132), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n722), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(G125), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n251), .B1(new_n716), .B2(new_n1109), .C1(new_n221), .C2(new_n704), .ZN(new_n1110));
  INV_X1    g0910(.A(G137), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n730), .A2(new_n1111), .B1(new_n766), .B2(new_n717), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1095), .A2(new_n1099), .B1(new_n1103), .B2(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n689), .B1(new_n279), .B2(new_n756), .C1(new_n1114), .C2(new_n702), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n870), .B2(new_n691), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n904), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1093), .A2(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(new_n324), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n614), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n327), .A3(new_n805), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n614), .B(new_n1120), .C1(new_n323), .C2(new_n631), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n692), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n251), .A2(G41), .ZN(new_n1131));
  AOI211_X1 g0931(.A(G50), .B(new_n1131), .C1(new_n248), .C2(new_n263), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n296), .B2(new_n707), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n740), .A2(G58), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n769), .B2(new_n716), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(new_n724), .C2(new_n991), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n730), .A2(new_n461), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n960), .B(new_n1137), .C1(G116), .C2(new_n712), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1136), .B(new_n1138), .C1(new_n255), .C2(new_n722), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT58), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1132), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n713), .A2(new_n1109), .B1(new_n766), .B2(new_n988), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n721), .A2(G128), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1105), .A2(new_n708), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n760), .C2(new_n1111), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1142), .B(new_n1145), .C1(G132), .C2(new_n729), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n740), .A2(G159), .ZN(new_n1149));
  AOI211_X1 g0949(.A(G33), .B(G41), .C1(new_n742), .C2(G124), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1141), .B1(new_n1140), .B2(new_n1139), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n694), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n750), .C1(G50), .C2(new_n756), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1130), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n896), .A2(G330), .A3(new_n1129), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1129), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n892), .A2(new_n860), .B1(new_n894), .B2(KEYINPUT40), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n643), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n874), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n870), .A2(new_n873), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1163), .A2(new_n1157), .A3(new_n1160), .A4(new_n861), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1156), .B1(new_n1165), .B2(new_n904), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1091), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1060), .A2(new_n1071), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT125), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT125), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1168), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1085), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1172), .A3(new_n1165), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1169), .A2(new_n1172), .A3(KEYINPUT57), .A4(new_n1165), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1019), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1166), .B1(new_n1175), .B2(new_n1177), .ZN(G375));
  INV_X1    g0978(.A(new_n1069), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1168), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n928), .A3(new_n1091), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1069), .A2(new_n904), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n689), .B1(G68), .B2(new_n756), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n992), .B1(new_n760), .B2(new_n255), .C1(new_n769), .C2(new_n722), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G116), .A2(new_n729), .B1(new_n712), .B2(G294), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n251), .B1(new_n740), .B2(G77), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n708), .A2(G97), .B1(new_n742), .B2(G303), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n712), .A2(G132), .B1(new_n727), .B2(G50), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n708), .A2(G159), .B1(new_n742), .B2(G128), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n251), .A4(new_n1134), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n724), .A2(G150), .B1(new_n729), .B2(new_n1105), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n1111), .B2(new_n722), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1184), .A2(new_n1188), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1183), .B1(new_n694), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n813), .B2(new_n692), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1182), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1181), .A2(new_n1198), .ZN(G381));
  NAND2_X1  g0999(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1019), .A3(new_n1176), .ZN(new_n1201));
  INV_X1    g1001(.A(G378), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(new_n1166), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n948), .A2(new_n970), .A3(new_n1031), .A4(new_n1054), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1021), .B(KEYINPUT110), .ZN(new_n1205));
  INV_X1    g1005(.A(G396), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1015), .A4(new_n1020), .ZN(new_n1207));
  INV_X1    g1007(.A(G384), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1181), .A2(new_n1208), .A3(new_n1198), .ZN(new_n1209));
  OR4_X1    g1009(.A1(new_n1203), .A2(new_n1204), .A3(new_n1207), .A4(new_n1209), .ZN(G407));
  INV_X1    g1010(.A(new_n1203), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n632), .A2(G213), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(G407), .A2(G213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT126), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(G407), .A2(KEYINPUT126), .A3(G213), .A4(new_n1214), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(G409));
  NAND2_X1  g1019(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1180), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1179), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1019), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT127), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1029), .B1(new_n1220), .B2(new_n1180), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT127), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1226), .A3(new_n1222), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G384), .B1(new_n1228), .B2(new_n1198), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1208), .B(new_n1197), .C1(new_n1224), .C2(new_n1227), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1166), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(G378), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1169), .A2(new_n1172), .A3(new_n928), .A4(new_n1165), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1213), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1176), .A2(new_n1019), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1232), .B1(new_n1236), .B2(new_n1200), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1231), .B(new_n1235), .C1(new_n1237), .C2(new_n1202), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT62), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  OAI211_X1 g1040(.A(G2897), .B(new_n1213), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1227), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1226), .B1(new_n1225), .B2(new_n1222), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1198), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1208), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1228), .A2(G384), .A3(new_n1198), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1213), .A2(G2897), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1202), .B1(new_n1201), .B2(new_n1166), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1212), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1241), .B(new_n1248), .C1(new_n1249), .C2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G375), .A2(G378), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1231), .A4(new_n1235), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1239), .A2(new_n1240), .A3(new_n1252), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1207), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(G390), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1204), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1204), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1256), .A2(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1247), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1253), .A2(new_n1235), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1238), .A2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1231), .A4(new_n1235), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n1271), .A3(new_n1262), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1264), .A2(new_n1273), .ZN(G405));
  OAI21_X1  g1074(.A(new_n1231), .B1(new_n1211), .B2(new_n1249), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1253), .B(new_n1203), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(new_n1262), .ZN(G402));
endmodule


