//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  OR3_X1    g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  OR2_X1    g002(.A1(G125), .A2(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(G125), .A2(G140), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n188), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(KEYINPUT72), .ZN(new_n196));
  OAI211_X1 g010(.A(G146), .B(new_n188), .C1(new_n191), .C2(new_n192), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G119), .B(G128), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT24), .B(G110), .Z(new_n201));
  AOI22_X1  g015(.A1(new_n196), .A2(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G128), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n206), .C1(G119), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G110), .ZN(new_n209));
  XOR2_X1   g023(.A(new_n209), .B(KEYINPUT70), .Z(new_n210));
  NAND2_X1  g024(.A1(new_n202), .A2(new_n210), .ZN(new_n211));
  OAI22_X1  g025(.A1(new_n208), .A2(G110), .B1(new_n200), .B2(new_n201), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n189), .B2(new_n190), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(new_n197), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n217), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n211), .A2(new_n220), .A3(new_n215), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT25), .B1(new_n224), .B2(G902), .ZN(new_n225));
  INV_X1    g039(.A(G217), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(G234), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n222), .A2(new_n229), .A3(new_n227), .A4(new_n223), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n228), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n222), .A2(new_n227), .A3(new_n232), .A4(new_n223), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(G472), .A2(G902), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  INV_X1    g050(.A(G116), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(G119), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n203), .A2(KEYINPUT67), .A3(G116), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n238), .B(new_n239), .C1(G116), .C2(new_n203), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n240), .B(new_n241), .Z(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT11), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(G137), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(G137), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(new_n244), .C1(new_n245), .C2(G137), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT11), .A3(G134), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n247), .A2(new_n248), .A3(new_n250), .A4(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(G131), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT64), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(KEYINPUT64), .A3(G146), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n258), .A2(new_n259), .B1(G143), .B2(new_n194), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT0), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(new_n207), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n207), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n194), .A2(G143), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n265), .A2(new_n256), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n263), .A2(new_n264), .B1(new_n266), .B2(new_n262), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n254), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n269), .A3(G128), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n207), .B1(new_n265), .B2(KEYINPUT1), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n260), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n248), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n245), .A2(G137), .ZN(new_n274));
  OAI21_X1  g088(.A(G131), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n272), .B(new_n275), .C1(G131), .C2(new_n253), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT30), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n254), .A2(new_n267), .A3(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n280), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n243), .B(new_n279), .C1(new_n283), .C2(KEYINPUT30), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n268), .A2(new_n242), .A3(new_n276), .ZN(new_n286));
  INV_X1    g100(.A(G237), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT68), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G237), .ZN(new_n290));
  AOI21_X1  g104(.A(G953), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G210), .ZN(new_n292));
  INV_X1    g106(.A(G101), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n294), .B(new_n295), .Z(new_n296));
  NAND4_X1  g110(.A1(new_n284), .A2(new_n285), .A3(new_n286), .A4(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n286), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT28), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n286), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n299), .B(new_n301), .C1(new_n283), .C2(new_n242), .ZN(new_n302));
  INV_X1    g116(.A(new_n296), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT30), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n277), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n280), .A2(new_n276), .A3(new_n282), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n298), .B1(new_n309), .B2(new_n243), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n285), .B1(new_n310), .B2(new_n296), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n235), .B1(new_n305), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT32), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT32), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n314), .B(new_n235), .C1(new_n305), .C2(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n301), .ZN(new_n317));
  OR3_X1    g131(.A1(new_n278), .A2(KEYINPUT69), .A3(new_n242), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT69), .B1(new_n278), .B2(new_n242), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n286), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n317), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n303), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n302), .A2(new_n303), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n322), .B1(new_n310), .B2(new_n296), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G472), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n234), .B1(new_n316), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n330));
  INV_X1    g144(.A(G104), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G107), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR4_X1   g148(.A1(new_n331), .A2(KEYINPUT74), .A3(KEYINPUT3), .A4(G107), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(G107), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n336), .A2(KEYINPUT75), .A3(new_n293), .A4(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G107), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n339), .A3(G104), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT3), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n333), .A2(new_n330), .A3(new_n339), .A4(G104), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n341), .A2(new_n293), .A3(new_n337), .A4(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n337), .A3(new_n342), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G101), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n338), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n349), .A3(G101), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n351), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n243), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n337), .B(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n339), .A2(KEYINPUT77), .A3(G104), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT77), .B1(new_n339), .B2(G104), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n293), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n338), .B2(new_n345), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT5), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n203), .A3(G116), .ZN(new_n364));
  OAI211_X1 g178(.A(G113), .B(new_n364), .C1(new_n240), .C2(new_n363), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n240), .A2(new_n241), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n355), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(G110), .B(G122), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n355), .A2(new_n368), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n370), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(KEYINPUT6), .A3(new_n374), .ZN(new_n375));
  OR3_X1    g189(.A1(new_n369), .A2(KEYINPUT6), .A3(new_n371), .ZN(new_n376));
  MUX2_X1   g190(.A(new_n272), .B(new_n267), .S(G125), .Z(new_n377));
  NAND2_X1  g191(.A1(new_n218), .A2(G224), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(KEYINPUT7), .A3(new_n378), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT85), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n362), .B(new_n367), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n370), .B(KEYINPUT8), .Z(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n378), .A2(KEYINPUT7), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(new_n385), .A3(new_n387), .A4(new_n372), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n380), .A2(new_n388), .A3(new_n227), .ZN(new_n389));
  OAI21_X1  g203(.A(G210), .B1(G237), .B2(G902), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n390), .A2(KEYINPUT86), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n391), .ZN(new_n393));
  OAI21_X1  g207(.A(G214), .B1(G237), .B2(G902), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n394), .B(KEYINPUT84), .Z(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G116), .B(G122), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n339), .ZN(new_n401));
  XNOR2_X1  g215(.A(G128), .B(G143), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n245), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(KEYINPUT13), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n207), .A2(KEYINPUT13), .A3(G143), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(G134), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT91), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n400), .A2(new_n339), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT92), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n402), .B(new_n245), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n237), .A2(KEYINPUT14), .A3(G122), .ZN(new_n413));
  INV_X1    g227(.A(new_n400), .ZN(new_n414));
  OAI211_X1 g228(.A(G107), .B(new_n413), .C1(new_n414), .C2(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT9), .B(G234), .Z(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(G217), .A3(new_n218), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT93), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n420), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n227), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT94), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT94), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n426), .A3(new_n227), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n399), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n398), .B1(new_n424), .B2(KEYINPUT94), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(G234), .A2(G237), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n431), .A2(G952), .A3(new_n218), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n431), .A2(G902), .A3(G953), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT21), .B(G898), .Z(new_n436));
  OAI21_X1  g250(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G475), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n255), .A2(KEYINPUT87), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n291), .A2(G214), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n291), .B2(G214), .ZN(new_n441));
  OAI211_X1 g255(.A(KEYINPUT18), .B(G131), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n191), .A2(G146), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n214), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n189), .A2(new_n190), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(new_n194), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT88), .B1(new_n447), .B2(new_n213), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n291), .A2(G214), .ZN(new_n450));
  INV_X1    g264(.A(new_n439), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT18), .A2(G131), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n291), .A2(G214), .A3(new_n439), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n442), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT89), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n442), .A2(new_n449), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n331), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT17), .B(G131), .C1(new_n440), .C2(new_n441), .ZN(new_n463));
  OAI21_X1  g277(.A(G131), .B1(new_n440), .B2(new_n441), .ZN(new_n464));
  INV_X1    g278(.A(G131), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n452), .A2(new_n465), .A3(new_n454), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT17), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n196), .A2(new_n463), .A3(new_n468), .A4(new_n199), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n460), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n197), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n191), .B1(new_n472), .B2(KEYINPUT19), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n191), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n475), .B2(new_n194), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n464), .A2(new_n466), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n462), .B1(new_n460), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n438), .B(new_n227), .C1(new_n470), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n462), .B1(new_n460), .B2(new_n469), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n227), .B1(new_n470), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G475), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n460), .A2(new_n469), .A3(new_n462), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n457), .A2(new_n459), .B1(new_n477), .B2(new_n476), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n462), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n488), .A2(KEYINPUT20), .A3(new_n438), .A4(new_n227), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n482), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n430), .A2(new_n437), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n396), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT10), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n357), .A2(new_n360), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G101), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n270), .B1(new_n266), .B2(new_n271), .ZN(new_n497));
  INV_X1    g311(.A(new_n345), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n343), .A2(new_n344), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n496), .B(new_n497), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT79), .B1(new_n362), .B2(new_n497), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n494), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT82), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n272), .A2(KEYINPUT10), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n354), .A2(new_n267), .B1(new_n362), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n254), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n507), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(KEYINPUT82), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n509), .A3(new_n507), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT80), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT80), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n504), .A2(new_n514), .A3(new_n509), .A4(new_n507), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n508), .A2(new_n511), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G110), .B(G140), .ZN(new_n517));
  INV_X1    g331(.A(G227), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(G953), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n517), .B(new_n519), .Z(new_n520));
  OAI21_X1  g334(.A(KEYINPUT83), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n515), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n502), .A2(new_n503), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n362), .A2(new_n272), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n254), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n254), .B(new_n526), .C1(new_n523), .C2(new_n524), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n522), .A2(new_n520), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n507), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n500), .A2(new_n501), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n362), .A2(KEYINPUT79), .A3(new_n497), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT10), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT82), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n508), .A3(new_n254), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n522), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT83), .ZN(new_n539));
  INV_X1    g353(.A(new_n520), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n521), .A2(new_n531), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G469), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n227), .ZN(new_n544));
  NAND2_X1  g358(.A1(G469), .A2(G902), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n522), .A2(new_n529), .A3(new_n530), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n540), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n516), .A2(new_n520), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(G469), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n418), .A2(new_n227), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G221), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n552), .B(KEYINPUT73), .Z(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n329), .A2(new_n493), .A3(new_n550), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(G101), .ZN(G3));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n305), .A2(new_n311), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(new_n227), .ZN(new_n559));
  INV_X1    g373(.A(new_n312), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n559), .A2(new_n560), .A3(new_n234), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n550), .A2(new_n561), .A3(new_n554), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT95), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n550), .A2(new_n561), .A3(new_n564), .A4(new_n554), .ZN(new_n565));
  INV_X1    g379(.A(new_n394), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n380), .A2(new_n388), .A3(new_n227), .A4(new_n390), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n390), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n389), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(KEYINPUT96), .A3(new_n567), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n570), .B2(new_n573), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n563), .A2(new_n565), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT98), .B(G478), .Z(new_n579));
  NAND2_X1  g393(.A1(new_n424), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n581));
  INV_X1    g395(.A(new_n422), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n417), .A2(new_n420), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n421), .A2(KEYINPUT33), .A3(new_n422), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n397), .A2(G902), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n491), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n437), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n578), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT34), .B(G104), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  INV_X1    g409(.A(new_n437), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n430), .A2(new_n596), .A3(new_n490), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT99), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n578), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n339), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT100), .B(KEYINPUT35), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G9));
  NOR2_X1   g416(.A1(new_n221), .A2(KEYINPUT36), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n216), .B(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n227), .A3(new_n232), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n231), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n493), .A2(new_n550), .A3(new_n554), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n305), .A2(new_n311), .ZN(new_n608));
  OAI21_X1  g422(.A(G472), .B1(new_n608), .B2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n312), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT37), .B(G110), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  AND2_X1   g427(.A1(new_n550), .A2(new_n554), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n606), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n575), .A2(new_n576), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n316), .A2(new_n328), .ZN(new_n617));
  INV_X1    g431(.A(G900), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n432), .B1(new_n434), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n490), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n430), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n615), .A2(new_n616), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n207), .ZN(G30));
  XOR2_X1   g439(.A(new_n619), .B(KEYINPUT39), .Z(new_n626));
  NAND2_X1  g440(.A1(new_n614), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT40), .Z(new_n628));
  NAND2_X1  g442(.A1(new_n392), .A2(new_n393), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n606), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n227), .B1(new_n320), .B2(new_n296), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n310), .A2(new_n303), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n316), .A2(new_n635), .ZN(new_n636));
  NOR4_X1   g450(.A1(new_n636), .A2(new_n491), .A3(new_n430), .A4(new_n566), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n628), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G143), .ZN(G45));
  NAND2_X1  g453(.A1(new_n617), .A2(new_n606), .ZN(new_n640));
  INV_X1    g454(.A(new_n619), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n490), .A2(new_n588), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n490), .A2(new_n588), .A3(KEYINPUT102), .A4(new_n641), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n614), .A3(new_n577), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G146), .ZN(G48));
  NAND2_X1  g463(.A1(new_n542), .A2(new_n227), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G469), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n554), .A3(new_n544), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n651), .A2(KEYINPUT103), .A3(new_n554), .A4(new_n544), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n654), .A2(new_n577), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n329), .A3(new_n592), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT41), .B(G113), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G15));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n656), .A2(new_n660), .A3(new_n329), .A4(new_n598), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n654), .A2(new_n329), .A3(new_n577), .A4(new_n655), .ZN(new_n662));
  INV_X1    g476(.A(new_n598), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT104), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G116), .ZN(G18));
  INV_X1    g480(.A(new_n492), .ZN(new_n667));
  INV_X1    g481(.A(new_n640), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n656), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G119), .ZN(G21));
  NOR2_X1   g484(.A1(new_n430), .A2(new_n491), .ZN(new_n671));
  INV_X1    g485(.A(new_n234), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n297), .B1(new_n321), .B2(new_n296), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n235), .B1(new_n673), .B2(new_n311), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n672), .A2(new_n609), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n437), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n656), .A2(new_n671), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G122), .ZN(G24));
  NAND3_X1  g493(.A1(new_n609), .A2(new_n674), .A3(new_n606), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n646), .A2(KEYINPUT105), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n644), .A2(new_n682), .A3(new_n645), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n680), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n654), .A2(new_n577), .A3(new_n655), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n187), .ZN(G27));
  NAND2_X1  g504(.A1(new_n547), .A2(KEYINPUT107), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n546), .A2(new_n692), .A3(new_n540), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(G469), .A3(new_n548), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n544), .A2(new_n545), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n566), .B1(new_n392), .B2(new_n393), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n695), .A2(new_n554), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n681), .A2(new_n683), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n697), .A2(KEYINPUT42), .A3(new_n329), .A4(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n329), .A2(new_n695), .A3(new_n554), .A4(new_n696), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n681), .A2(new_n683), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G131), .ZN(G33));
  NAND3_X1  g519(.A1(new_n697), .A2(new_n329), .A3(new_n622), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G134), .ZN(G36));
  NAND2_X1  g521(.A1(new_n547), .A2(new_n548), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n691), .A2(new_n548), .A3(new_n693), .ZN(new_n711));
  OAI211_X1 g525(.A(G469), .B(new_n710), .C1(new_n711), .C2(new_n709), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT46), .A3(new_n545), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(KEYINPUT108), .A3(new_n544), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT108), .B1(new_n713), .B2(new_n544), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT46), .B1(new_n712), .B2(new_n545), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n553), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n626), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n719), .A2(KEYINPUT109), .ZN(new_n720));
  INV_X1    g534(.A(new_n696), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n491), .A2(new_n588), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT43), .Z(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n610), .A3(new_n606), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n719), .A2(KEYINPUT109), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n720), .A2(new_n726), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G137), .ZN(G39));
  OR2_X1    g544(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n646), .B(new_n721), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n617), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n234), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  AND2_X1   g550(.A1(new_n661), .A2(new_n664), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n657), .A2(new_n669), .A3(new_n678), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n592), .A3(KEYINPUT111), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n744));
  INV_X1    g558(.A(new_n429), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n425), .A2(new_n427), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n399), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT112), .B1(new_n428), .B2(new_n429), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n490), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n742), .A2(new_n749), .A3(new_n437), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n396), .B2(new_n591), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n743), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n563), .A2(new_n565), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n555), .B1(new_n607), .B2(new_n610), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n741), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n755), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n563), .A2(new_n565), .A3(new_n753), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(KEYINPUT113), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n697), .A2(new_n684), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n734), .A2(new_n721), .A3(new_n621), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n747), .A2(new_n748), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n614), .A3(new_n606), .A4(new_n763), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n704), .A2(new_n706), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n739), .A2(new_n740), .A3(new_n760), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n654), .A2(new_n577), .A3(new_n671), .A4(new_n655), .ZN(new_n767));
  OAI22_X1  g581(.A1(new_n591), .A2(new_n662), .B1(new_n767), .B2(new_n676), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n654), .A2(new_n655), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n769), .A2(new_n616), .A3(new_n492), .A4(new_n640), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n760), .A2(new_n771), .A3(new_n765), .A4(new_n665), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT114), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n774));
  OR3_X1    g588(.A1(new_n615), .A2(new_n616), .A3(new_n623), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n775), .B(new_n648), .C1(new_n687), .C2(new_n688), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n636), .A2(new_n606), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n554), .A3(new_n641), .A4(new_n695), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n577), .A2(new_n671), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n774), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n656), .A2(KEYINPUT106), .A3(new_n684), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n685), .A2(new_n686), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n624), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n780), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(KEYINPUT52), .A3(new_n648), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n766), .A2(new_n773), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n789), .B1(new_n781), .B2(new_n786), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n766), .A3(new_n773), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT54), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT115), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n796));
  INV_X1    g610(.A(new_n772), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n791), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n790), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n793), .A2(new_n800), .A3(KEYINPUT54), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n651), .A2(new_n544), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n731), .B(new_n732), .C1(new_n554), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n723), .A2(new_n432), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(new_n675), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n805), .A2(new_n696), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n769), .A2(new_n721), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n807), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(new_n680), .ZN(new_n814));
  NOR2_X1   g628(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n769), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n808), .A3(new_n566), .A4(new_n631), .ZN(new_n817));
  NAND2_X1  g631(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n672), .A2(new_n812), .A3(new_n432), .A4(new_n636), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n491), .A3(new_n589), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n809), .A2(new_n814), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n811), .B(new_n822), .Z(new_n823));
  AND2_X1   g637(.A1(new_n808), .A2(new_n656), .ZN(new_n824));
  INV_X1    g638(.A(new_n329), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n813), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(KEYINPUT48), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n218), .A2(G952), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n820), .B2(new_n590), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n830), .B(new_n832), .C1(KEYINPUT48), .C2(new_n829), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n802), .A2(new_n823), .A3(new_n824), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(G952), .A2(G953), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n804), .A2(KEYINPUT49), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n631), .ZN(new_n837));
  INV_X1    g651(.A(new_n722), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n672), .A2(new_n838), .A3(new_n395), .A4(new_n554), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT110), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n804), .A2(KEYINPUT49), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n636), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n834), .A2(new_n835), .B1(new_n837), .B2(new_n842), .ZN(G75));
  NAND2_X1  g657(.A1(new_n375), .A2(new_n376), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n379), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n788), .A2(new_n789), .B1(new_n797), .B2(new_n791), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n227), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT120), .B1(new_n848), .B2(G210), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n850));
  XNOR2_X1  g664(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n849), .B2(new_n850), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n218), .A2(G952), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n848), .A2(G210), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n850), .ZN(new_n859));
  INV_X1    g673(.A(new_n851), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n845), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n854), .A2(new_n856), .A3(new_n863), .ZN(G51));
  INV_X1    g678(.A(new_n542), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n799), .A2(KEYINPUT121), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n790), .A2(new_n798), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT54), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n847), .A2(new_n869), .A3(new_n796), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n545), .B(KEYINPUT57), .Z(new_n872));
  AOI21_X1  g686(.A(new_n865), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n847), .A2(new_n227), .A3(new_n712), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n856), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT122), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n856), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(G54));
  NAND3_X1  g693(.A1(new_n848), .A2(KEYINPUT58), .A3(G475), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(new_n488), .Z(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n855), .ZN(G60));
  AND2_X1   g696(.A1(new_n584), .A2(new_n585), .ZN(new_n883));
  XNOR2_X1  g697(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n397), .A2(new_n227), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n802), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n871), .A2(new_n883), .A3(new_n886), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n887), .A2(new_n888), .A3(new_n855), .ZN(G63));
  XNOR2_X1  g703(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(G217), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT60), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n867), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n867), .A2(KEYINPUT124), .A3(new_n893), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n224), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n856), .ZN(new_n899));
  INV_X1    g713(.A(new_n604), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n896), .B2(new_n897), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n891), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n901), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n856), .A3(new_n898), .A4(new_n890), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(G66));
  AOI21_X1  g719(.A(new_n218), .B1(new_n436), .B2(G224), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n739), .A2(new_n760), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n218), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n844), .B1(G898), .B2(new_n218), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n908), .B(new_n909), .Z(G69));
  XNOR2_X1  g724(.A(new_n309), .B(new_n475), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n735), .A2(new_n729), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n779), .A2(new_n825), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n720), .A2(new_n727), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n704), .A2(new_n706), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n776), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n913), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n912), .B1(new_n918), .B2(new_n218), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(G900), .B2(new_n218), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n329), .B1(new_n590), .B2(new_n749), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n627), .A2(new_n721), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n638), .A2(new_n648), .A3(new_n784), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT62), .Z(new_n924));
  NAND3_X1  g738(.A1(new_n913), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n218), .A3(new_n912), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(G953), .B1(new_n518), .B2(new_n618), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n928), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n920), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(G72));
  NAND2_X1  g746(.A1(G472), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT63), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n925), .B2(new_n907), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n855), .B1(new_n937), .B2(new_n634), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n918), .B2(new_n907), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n310), .A3(new_n303), .ZN(new_n940));
  INV_X1    g754(.A(new_n634), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n310), .A2(new_n303), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n793), .A2(new_n941), .A3(new_n936), .A4(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(G57));
endmodule


