//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  OR2_X1    g000(.A1(KEYINPUT66), .A2(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT66), .A2(G128), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G119), .A3(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  AOI21_X1  g008(.A(KEYINPUT23), .B1(new_n190), .B2(G119), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(new_n191), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .A4(new_n188), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI22_X1  g012(.A1(new_n193), .A2(new_n194), .B1(new_n198), .B2(G110), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(KEYINPUT16), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(new_n208), .B2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n199), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n198), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT78), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n212), .A2(G110), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n193), .A2(new_n194), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n200), .A3(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n201), .A2(new_n203), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(new_n216), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(new_n204), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n221));
  AOI21_X1  g035(.A(G146), .B1(new_n221), .B2(new_n217), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n215), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n210), .B1(new_n214), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT80), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n204), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n208), .A2(G146), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n226), .A2(new_n227), .B1(new_n193), .B2(new_n194), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n212), .A2(G110), .A3(new_n213), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n228), .A2(new_n229), .B1(new_n199), .B2(new_n209), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G953), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(G221), .A3(G234), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT79), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G137), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n225), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n230), .A2(new_n231), .A3(new_n237), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G217), .ZN(new_n243));
  INV_X1    g057(.A(G902), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(G234), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G902), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(new_n244), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n241), .A2(KEYINPUT25), .A3(new_n244), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n248), .B1(new_n253), .B2(new_n245), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  OR2_X1    g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n204), .A2(G143), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n256), .B(new_n257), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n258), .B2(G146), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n204), .A2(KEYINPUT64), .A3(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(G146), .ZN(new_n265));
  INV_X1    g079(.A(new_n256), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n263), .A2(new_n264), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n271));
  INV_X1    g085(.A(G134), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(G137), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(G137), .ZN(new_n274));
  INV_X1    g088(.A(G137), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT11), .A3(G134), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G131), .ZN(new_n278));
  INV_X1    g092(.A(G131), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n273), .A2(new_n276), .A3(new_n279), .A4(new_n274), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n261), .A2(KEYINPUT70), .A3(new_n267), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n270), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n275), .A2(G134), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n272), .A2(G137), .ZN(new_n285));
  OAI21_X1  g099(.A(G131), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n288));
  NOR2_X1   g102(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(G128), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(G143), .B(G146), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n204), .A2(G143), .ZN(new_n295));
  AND2_X1   g109(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(new_n289), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n187), .A2(new_n188), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n287), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n283), .A2(KEYINPUT30), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT30), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n268), .B1(new_n280), .B2(new_n278), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n280), .A2(new_n286), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n297), .A2(new_n298), .ZN(new_n305));
  INV_X1    g119(.A(new_n294), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n296), .A2(new_n289), .A3(new_n190), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n308), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n304), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n302), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G116), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G119), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT68), .B1(new_n314), .B2(G116), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n312), .A3(G119), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT2), .A2(G113), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n321));
  INV_X1    g135(.A(G113), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n319), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n318), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n318), .B2(new_n325), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n301), .A2(new_n311), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT71), .B(new_n326), .C1(new_n328), .C2(new_n329), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n333), .A2(new_n300), .A3(new_n283), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G101), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(KEYINPUT72), .A2(G237), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT72), .A2(G237), .ZN(new_n340));
  AOI21_X1  g154(.A(G953), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G210), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n341), .B2(G210), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n345), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n343), .A3(new_n337), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n336), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n307), .A2(new_n309), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n261), .A2(new_n267), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n355), .A2(new_n287), .B1(new_n356), .B2(new_n281), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n318), .A2(new_n325), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n318), .A2(new_n325), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n318), .A2(new_n325), .A3(new_n327), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n357), .A2(new_n362), .A3(KEYINPUT75), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n356), .A2(new_n281), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n300), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n366), .B2(new_n330), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n354), .B1(new_n368), .B2(new_n335), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n347), .B2(new_n350), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n346), .A2(new_n349), .A3(KEYINPUT74), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n335), .A2(new_n354), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n353), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n335), .A2(new_n354), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n333), .A2(new_n334), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n283), .A2(new_n300), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n335), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n379), .B1(KEYINPUT28), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n351), .A2(KEYINPUT29), .ZN(new_n385));
  AOI21_X1  g199(.A(G902), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n353), .B(KEYINPUT77), .C1(new_n369), .C2(new_n375), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n378), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(G472), .A2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n373), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n369), .B2(new_n379), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n331), .A2(new_n335), .A3(new_n351), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT31), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT73), .B(KEYINPUT31), .Z(new_n395));
  NAND4_X1  g209(.A1(new_n331), .A2(new_n335), .A3(new_n351), .A4(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n390), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n388), .A2(G472), .B1(KEYINPUT32), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT75), .B1(new_n357), .B2(new_n362), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n366), .A2(new_n364), .A3(new_n330), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n335), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT28), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n373), .B1(new_n403), .B2(new_n374), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n394), .A2(new_n396), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n389), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT76), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n409));
  OAI211_X1 g223(.A(KEYINPUT76), .B(new_n389), .C1(new_n404), .C2(new_n405), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n255), .B1(new_n399), .B2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(KEYINPUT72), .A2(G237), .ZN(new_n413));
  NOR2_X1   g227(.A1(KEYINPUT72), .A2(G237), .ZN(new_n414));
  OAI211_X1 g228(.A(G214), .B(new_n233), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n258), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT72), .B(G237), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(G143), .A3(G214), .A4(new_n233), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G131), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT17), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n416), .A2(new_n418), .A3(new_n279), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n220), .A2(new_n222), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n423), .B(new_n424), .C1(new_n421), .C2(new_n420), .ZN(new_n425));
  XNOR2_X1  g239(.A(G113), .B(G122), .ZN(new_n426));
  INV_X1    g240(.A(G104), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(KEYINPUT18), .A2(G131), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n416), .A2(new_n418), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT90), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n416), .A2(new_n418), .A3(new_n432), .A4(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  INV_X1    g249(.A(new_n429), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n204), .B1(new_n201), .B2(new_n203), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n207), .A2(new_n204), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT89), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n205), .B2(new_n437), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n419), .A2(new_n436), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n434), .A2(new_n435), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n435), .B1(new_n434), .B2(new_n443), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n425), .B(new_n428), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n420), .A2(new_n422), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n207), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT93), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n218), .A2(KEYINPUT19), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT93), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n452), .A3(new_n207), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n450), .A2(new_n204), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n227), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n434), .A2(new_n443), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT91), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n434), .A2(new_n435), .A3(new_n443), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n446), .B1(new_n460), .B2(new_n428), .ZN(new_n461));
  NOR3_X1   g275(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(G475), .A2(G902), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n446), .B(KEYINPUT94), .C1(new_n460), .C2(new_n428), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n463), .B1(new_n468), .B2(KEYINPUT20), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n425), .B1(new_n444), .B2(new_n445), .ZN(new_n470));
  INV_X1    g284(.A(new_n428), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n472), .B2(new_n446), .ZN(new_n473));
  INV_X1    g287(.A(G475), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G122), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(G116), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(G116), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G107), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n258), .A2(G128), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT13), .Z(new_n484));
  NAND3_X1  g298(.A1(new_n187), .A2(G143), .A3(new_n188), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G134), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n483), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n482), .B(new_n487), .C1(G134), .C2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n272), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n478), .A2(KEYINPUT14), .ZN(new_n491));
  OR3_X1    g305(.A1(new_n476), .A2(KEYINPUT14), .A3(G116), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT95), .A4(new_n479), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n493), .B(G107), .C1(KEYINPUT95), .C2(new_n492), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n480), .A2(new_n481), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n489), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT9), .B(G234), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n498), .A2(new_n243), .A3(G953), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n497), .A2(new_n500), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n244), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G478), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI221_X1 g320(.A(new_n244), .B1(KEYINPUT15), .B2(new_n504), .C1(new_n501), .C2(new_n502), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n233), .A2(G952), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(G234), .B2(G237), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT21), .B(G898), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n510), .B(KEYINPUT96), .Z(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI211_X1 g326(.A(new_n244), .B(new_n233), .C1(G234), .C2(G237), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n506), .A2(new_n507), .A3(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n469), .A2(new_n475), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G214), .B1(G237), .B2(G902), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n518), .B(KEYINPUT84), .Z(new_n519));
  NAND2_X1  g333(.A1(new_n360), .A2(new_n361), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n481), .A2(G104), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n427), .A2(G107), .ZN(new_n522));
  OAI21_X1  g336(.A(G101), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT3), .B1(new_n427), .B2(G107), .ZN(new_n524));
  AOI21_X1  g338(.A(G101), .B1(new_n427), .B2(G107), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT3), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n481), .A3(G104), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT82), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT82), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n318), .A2(KEYINPUT5), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT5), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n322), .B1(new_n313), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n520), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n528), .A2(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n427), .A2(G107), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n524), .A2(new_n527), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G101), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n543), .B1(new_n544), .B2(new_n542), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n330), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT85), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT6), .ZN(new_n549));
  XNOR2_X1  g363(.A(G110), .B(G122), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n360), .A2(new_n361), .B1(new_n534), .B2(new_n536), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n553), .A2(new_n533), .B1(new_n330), .B2(new_n545), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n549), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT85), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n549), .B1(new_n554), .B2(new_n550), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n547), .A2(new_n551), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n307), .A2(new_n309), .A3(new_n202), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n202), .B1(new_n261), .B2(new_n267), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(KEYINPUT86), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n233), .A2(G224), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n567), .B(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n557), .A2(new_n560), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n537), .B1(new_n328), .B2(new_n329), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n529), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n538), .A2(new_n573), .A3(KEYINPUT87), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n550), .B(KEYINPUT8), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n573), .B2(KEYINPUT87), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT88), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n573), .A2(KEYINPUT87), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n579), .A2(new_n574), .A3(new_n580), .A4(new_n576), .ZN(new_n581));
  INV_X1    g395(.A(new_n566), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n569), .A2(KEYINPUT7), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n562), .A2(new_n564), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n561), .ZN(new_n585));
  OAI211_X1 g399(.A(KEYINPUT7), .B(new_n569), .C1(new_n565), .C2(new_n566), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n585), .A2(new_n586), .B1(new_n554), .B2(new_n550), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n578), .A2(new_n581), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n571), .A2(new_n588), .A3(new_n244), .ZN(new_n589));
  OAI21_X1  g403(.A(G210), .B1(G237), .B2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n571), .A2(new_n588), .A3(new_n244), .A4(new_n590), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n519), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n307), .B2(new_n309), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n533), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(KEYINPUT4), .A2(new_n528), .B1(new_n541), .B2(G101), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n541), .A2(KEYINPUT4), .A3(G101), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n270), .B(new_n282), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n523), .A2(new_n528), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT1), .ZN(new_n602));
  OAI21_X1  g416(.A(G128), .B1(new_n259), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n288), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n601), .B1(new_n604), .B2(new_n293), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n595), .ZN(new_n606));
  INV_X1    g420(.A(new_n281), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n597), .A2(new_n600), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n531), .A2(new_n309), .A3(new_n307), .A4(new_n532), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n605), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT12), .B1(new_n610), .B2(new_n281), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT12), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n612), .B(new_n607), .C1(new_n609), .C2(new_n605), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n608), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(G110), .B(G140), .ZN(new_n615));
  INV_X1    g429(.A(G227), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(G953), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n615), .B(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n533), .A2(new_n596), .B1(new_n605), .B2(new_n595), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n600), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n281), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n614), .A2(new_n618), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G469), .B1(new_n624), .B2(G902), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT83), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n607), .B1(new_n621), .B2(new_n600), .ZN(new_n627));
  AND4_X1   g441(.A1(new_n607), .A2(new_n597), .A3(new_n600), .A4(new_n606), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n618), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n608), .B(new_n619), .C1(new_n611), .C2(new_n613), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(G469), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n626), .A2(new_n631), .A3(new_n632), .A4(new_n244), .ZN(new_n633));
  AOI21_X1  g447(.A(G902), .B1(new_n629), .B2(new_n630), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n626), .B1(new_n634), .B2(new_n632), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n625), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G221), .B1(new_n498), .B2(G902), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT81), .Z(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n594), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n412), .A2(new_n517), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G101), .ZN(G3));
  NOR2_X1   g456(.A1(new_n504), .A2(new_n244), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n503), .B2(G478), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n497), .B(new_n499), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT33), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n645), .B1(new_n647), .B2(G478), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n469), .B2(new_n475), .ZN(new_n649));
  INV_X1    g463(.A(new_n519), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n552), .A2(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n651));
  AOI21_X1  g465(.A(G902), .B1(new_n651), .B2(new_n570), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n590), .B1(new_n652), .B2(new_n588), .ZN(new_n653));
  INV_X1    g467(.A(new_n593), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n515), .B(new_n650), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n254), .A2(new_n636), .A3(new_n639), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n244), .B1(new_n404), .B2(new_n405), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(G472), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n408), .A2(new_n659), .A3(new_n410), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT98), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NAND3_X1  g480(.A1(new_n465), .A2(new_n467), .A3(new_n462), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n465), .A2(KEYINPUT99), .A3(new_n467), .A4(new_n462), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n669), .A2(new_n670), .B1(KEYINPUT20), .B2(new_n468), .ZN(new_n671));
  INV_X1    g485(.A(new_n475), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n506), .A2(new_n507), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n671), .A2(new_n655), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n661), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  INV_X1    g492(.A(new_n660), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT25), .B1(new_n241), .B2(new_n244), .ZN(new_n680));
  AOI211_X1 g494(.A(new_n250), .B(G902), .C1(new_n239), .C2(new_n240), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n245), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n237), .A2(KEYINPUT36), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n224), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n246), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n640), .A2(new_n517), .A3(new_n679), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  XNOR2_X1  g503(.A(new_n509), .B(KEYINPUT100), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n692), .B2(new_n513), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n671), .A2(new_n674), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n686), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n399), .B2(new_n411), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(new_n696), .A3(new_n640), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  NAND2_X1  g512(.A1(new_n620), .A2(new_n623), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n610), .A2(new_n281), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n612), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n610), .A2(KEYINPUT12), .A3(new_n281), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n628), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n699), .B1(new_n703), .B2(new_n619), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n632), .B1(new_n704), .B2(new_n244), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n631), .A2(new_n632), .A3(new_n244), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT83), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n634), .A2(new_n626), .A3(new_n632), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n693), .B(KEYINPUT39), .Z(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n709), .A2(new_n638), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT40), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n469), .A2(new_n475), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n592), .A2(new_n593), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT38), .ZN(new_n719));
  INV_X1    g533(.A(new_n673), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n686), .A2(new_n720), .A3(new_n519), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n398), .A2(KEYINPUT32), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n391), .A2(KEYINPUT101), .A3(new_n383), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n393), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT101), .B1(new_n391), .B2(new_n383), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n244), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G472), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n411), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  AND4_X1   g542(.A1(new_n717), .A2(new_n719), .A3(new_n721), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n715), .A2(new_n716), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G143), .ZN(G45));
  INV_X1    g545(.A(new_n693), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n648), .B(new_n732), .C1(new_n469), .C2(new_n475), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n696), .A2(new_n734), .A3(new_n640), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  OR2_X1    g550(.A1(new_n634), .A2(new_n632), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n639), .B(new_n737), .C1(new_n633), .C2(new_n635), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT103), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n707), .A2(new_n708), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n639), .A4(new_n737), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n656), .A3(new_n412), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND3_X1  g560(.A1(new_n675), .A2(new_n743), .A3(new_n412), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT104), .B(G116), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G18));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n388), .A2(G472), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n411), .A2(new_n751), .A3(new_n722), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n517), .A3(new_n686), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n739), .A2(new_n594), .A3(new_n742), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n739), .A2(new_n594), .A3(new_n742), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(KEYINPUT105), .A3(new_n517), .A4(new_n696), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n314), .ZN(G21));
  NOR2_X1   g573(.A1(new_n384), .A2(new_n373), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n389), .B1(new_n760), .B2(new_n405), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n254), .A2(new_n515), .A3(new_n659), .A4(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n673), .B1(new_n469), .B2(new_n475), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n756), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n686), .A2(new_n659), .A3(new_n761), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n717), .A2(new_n768), .A3(new_n648), .A4(new_n732), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n769), .B2(new_n754), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n686), .A2(new_n659), .A3(new_n761), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n733), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n756), .A2(new_n772), .A3(KEYINPUT106), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT107), .B(G125), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G27));
  INV_X1    g590(.A(new_n412), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n592), .A2(new_n650), .A3(new_n593), .ZN(new_n778));
  NAND2_X1  g592(.A1(G469), .A2(G902), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT108), .Z(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n704), .B2(new_n632), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n707), .B2(new_n708), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n778), .A2(new_n783), .A3(new_n784), .A4(new_n638), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n782), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n638), .B1(new_n740), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n592), .A2(new_n650), .A3(new_n593), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT109), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n777), .B1(new_n786), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n733), .A2(KEYINPUT42), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n406), .A2(new_n409), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n255), .B1(new_n399), .B2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n734), .B(new_n795), .C1(new_n785), .C2(new_n790), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n792), .A2(new_n793), .B1(new_n796), .B2(KEYINPUT42), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G131), .ZN(G33));
  OAI211_X1 g612(.A(new_n412), .B(new_n694), .C1(new_n785), .C2(new_n790), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  NOR2_X1   g614(.A1(new_n469), .A2(new_n475), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n648), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT43), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n679), .A2(new_n695), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT44), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n807));
  OAI21_X1  g621(.A(G469), .B1(new_n624), .B2(KEYINPUT45), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n624), .A2(KEYINPUT45), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n808), .B2(new_n809), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n781), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT46), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n813), .A2(new_n814), .B1(new_n708), .B2(new_n707), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n638), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n711), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n804), .A2(KEYINPUT44), .A3(new_n805), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(new_n789), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n804), .A2(new_n805), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT44), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(KEYINPUT111), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n807), .A2(new_n819), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G137), .ZN(G39));
  INV_X1    g640(.A(new_n752), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n778), .A2(new_n254), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n734), .A3(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n817), .A2(KEYINPUT47), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n817), .A2(KEYINPUT47), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(new_n200), .ZN(G42));
  AND3_X1   g647(.A1(new_n648), .A2(new_n639), .A3(new_n650), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n740), .A2(new_n737), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n834), .B(new_n254), .C1(KEYINPUT49), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(KEYINPUT49), .B2(new_n835), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n719), .A2(new_n717), .A3(new_n728), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n747), .A2(new_n744), .A3(new_n765), .A4(new_n687), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT112), .B1(new_n801), .B2(new_n673), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n469), .A2(new_n720), .A3(new_n842), .A4(new_n475), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n655), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n661), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n641), .B(new_n662), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n758), .A2(new_n840), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n669), .A2(new_n670), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n468), .A2(KEYINPUT20), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n720), .A2(new_n672), .A3(new_n732), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT113), .B1(new_n671), .B2(new_n852), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n778), .A2(new_n709), .A3(new_n638), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(new_n696), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n772), .B1(new_n785), .B2(new_n790), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n799), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n799), .A2(new_n858), .A3(new_n859), .A4(KEYINPUT114), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n848), .A2(new_n864), .A3(new_n797), .ZN(new_n865));
  INV_X1    g679(.A(new_n763), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n682), .A2(new_n685), .A3(new_n732), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n783), .A2(new_n867), .A3(new_n638), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(new_n868), .A3(new_n728), .A4(new_n594), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n697), .A2(new_n735), .A3(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n870), .A2(new_n774), .A3(KEYINPUT52), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT52), .B1(new_n870), .B2(new_n774), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT53), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n840), .A2(new_n847), .ZN(new_n875));
  INV_X1    g689(.A(new_n758), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n875), .A2(new_n876), .A3(new_n797), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n770), .A2(new_n773), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n697), .A2(new_n735), .A3(new_n869), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n870), .A2(new_n774), .A3(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n877), .A2(new_n883), .A3(new_n884), .A4(new_n864), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n884), .A2(KEYINPUT115), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n865), .A2(KEYINPUT115), .A3(new_n884), .A4(new_n883), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT54), .B1(new_n874), .B2(new_n885), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n254), .A2(new_n659), .A3(new_n761), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n804), .A2(new_n691), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT50), .ZN(new_n898));
  INV_X1    g712(.A(new_n719), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n519), .A3(new_n743), .ZN(new_n900));
  OR3_X1    g714(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n898), .B1(new_n897), .B2(new_n900), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n897), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n830), .A2(new_n831), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n835), .A2(new_n639), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n789), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n691), .A2(new_n804), .A3(new_n743), .A4(new_n789), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n743), .A2(new_n789), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n254), .A2(new_n509), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n728), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n717), .A2(new_n648), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n908), .A2(new_n768), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n903), .A2(new_n907), .A3(KEYINPUT51), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n903), .A2(new_n907), .A3(new_n913), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n904), .A2(new_n756), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n508), .B(KEYINPUT117), .ZN(new_n919));
  INV_X1    g733(.A(new_n649), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n919), .B1(new_n911), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(KEYINPUT118), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT118), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n908), .A2(KEYINPUT48), .A3(new_n795), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT48), .B1(new_n908), .B2(new_n795), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AND4_X1   g740(.A1(new_n914), .A2(new_n917), .A3(new_n922), .A4(new_n926), .ZN(new_n927));
  AND4_X1   g741(.A1(new_n891), .A2(new_n894), .A3(new_n895), .A4(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(G952), .A2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n839), .B1(new_n928), .B2(new_n929), .ZN(G75));
  NOR2_X1   g744(.A1(new_n233), .A2(G952), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n651), .B(new_n570), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n874), .A2(new_n885), .A3(G210), .A4(G902), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n874), .A2(G902), .A3(new_n885), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT119), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n874), .A2(new_n885), .A3(new_n939), .A4(G902), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n938), .A2(new_n591), .A3(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n933), .A2(new_n935), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n931), .B(new_n936), .C1(new_n941), .C2(new_n942), .ZN(G51));
  XNOR2_X1  g757(.A(new_n780), .B(KEYINPUT57), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n874), .A2(KEYINPUT54), .A3(new_n885), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n892), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT120), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(new_n944), .C1(new_n945), .C2(new_n892), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n631), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n938), .A2(new_n940), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n810), .A2(new_n812), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n931), .B1(new_n950), .B2(new_n953), .ZN(G54));
  INV_X1    g768(.A(KEYINPUT121), .ZN(new_n955));
  INV_X1    g769(.A(new_n465), .ZN(new_n956));
  INV_X1    g770(.A(new_n467), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(KEYINPUT58), .A2(G475), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n951), .A2(new_n955), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n938), .A2(new_n940), .A3(new_n959), .ZN(new_n961));
  INV_X1    g775(.A(new_n958), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT121), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n931), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(G60));
  INV_X1    g779(.A(new_n647), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n643), .B(KEYINPUT59), .Z(new_n967));
  OAI211_X1 g781(.A(new_n966), .B(new_n967), .C1(new_n945), .C2(new_n892), .ZN(new_n968));
  INV_X1    g782(.A(new_n931), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n892), .B(new_n893), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n889), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n967), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n973), .B2(new_n647), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n874), .A2(new_n885), .A3(new_n684), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n969), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT61), .B1(new_n979), .B2(KEYINPUT122), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n242), .B1(new_n886), .B2(new_n976), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(new_n969), .A3(new_n978), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G66));
  AOI21_X1  g797(.A(new_n233), .B1(new_n511), .B2(G224), .ZN(new_n984));
  INV_X1    g798(.A(new_n848), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n233), .ZN(new_n986));
  INV_X1    g800(.A(G898), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n651), .B1(new_n987), .B2(G953), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n986), .B(new_n988), .ZN(G69));
  NAND2_X1  g803(.A1(new_n301), .A2(new_n311), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT123), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n990), .B(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n774), .A2(new_n697), .A3(new_n735), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT124), .Z(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n730), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  INV_X1    g811(.A(new_n832), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n844), .A2(new_n649), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n999), .A2(new_n412), .A3(new_n710), .A4(new_n857), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n825), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n995), .A2(new_n1002), .A3(new_n730), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n997), .A2(new_n1001), .A3(new_n233), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n993), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n616), .A2(G900), .A3(G953), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT125), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n866), .A2(new_n594), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n819), .A2(new_n795), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n1011), .A2(new_n797), .A3(new_n799), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n825), .A3(new_n998), .ZN(new_n1013));
  INV_X1    g827(.A(new_n995), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n825), .A2(new_n998), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1016), .A2(KEYINPUT125), .A3(new_n995), .A4(new_n1012), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1007), .B1(new_n1018), .B2(G953), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1006), .B1(new_n1019), .B2(new_n993), .ZN(G72));
  NAND3_X1  g834(.A1(new_n352), .A2(new_n331), .A3(new_n335), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1015), .A2(new_n1017), .A3(new_n848), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT126), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1021), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n336), .A2(new_n351), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n997), .A2(new_n1001), .A3(new_n848), .A4(new_n1003), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(new_n1025), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n336), .A2(new_n352), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT127), .Z(new_n1031));
  INV_X1    g845(.A(new_n393), .ZN(new_n1032));
  OR2_X1    g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n1033), .A2(new_n1024), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n889), .A2(new_n890), .A3(new_n1034), .ZN(new_n1035));
  NOR4_X1   g849(.A1(new_n1026), .A2(new_n1029), .A3(new_n931), .A4(new_n1035), .ZN(G57));
endmodule


