//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G110), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n191), .B2(G128), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(new_n197), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT24), .B(G110), .ZN(new_n201));
  INV_X1    g015(.A(new_n198), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(new_n192), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT16), .ZN(new_n209));
  OR3_X1    g023(.A1(new_n207), .A2(KEYINPUT16), .A3(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G146), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n206), .A2(new_n208), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT22), .B(G137), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n216), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G119), .ZN(new_n221));
  INV_X1    g035(.A(new_n195), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(new_n193), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n199), .A2(new_n198), .ZN(new_n224));
  OAI21_X1  g038(.A(G110), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT70), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G110), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n202), .A2(new_n192), .ZN(new_n231));
  INV_X1    g045(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n211), .ZN(new_n234));
  AOI21_X1  g048(.A(G146), .B1(new_n209), .B2(new_n210), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n215), .B(new_n219), .C1(new_n230), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n211), .A2(new_n214), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n200), .B2(new_n203), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n225), .A2(KEYINPUT70), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n228), .B1(new_n227), .B2(G110), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n235), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n243), .A2(new_n211), .B1(new_n231), .B2(new_n232), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n239), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n219), .B(KEYINPUT71), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT72), .B(new_n237), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n229), .A3(new_n226), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(new_n249), .A3(new_n215), .A4(new_n219), .ZN(new_n250));
  AOI211_X1 g064(.A(new_n190), .B(G902), .C1(new_n247), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n237), .A2(KEYINPUT72), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n246), .B1(new_n248), .B2(new_n215), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n250), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT25), .B1(new_n254), .B2(new_n188), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n189), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n189), .A2(G902), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT66), .ZN(new_n265));
  XOR2_X1   g079(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n266));
  INV_X1    g080(.A(KEYINPUT11), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G137), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G131), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n269), .A2(new_n271), .A3(new_n275), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n213), .A2(G143), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G146), .ZN(new_n280));
  AND2_X1   g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G143), .B(G146), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G128), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n277), .A2(KEYINPUT65), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(G128), .B1(new_n278), .B2(new_n280), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n279), .A2(KEYINPUT1), .A3(G146), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n283), .A2(new_n292), .A3(G128), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n268), .A2(G137), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n270), .A2(G134), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n276), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n285), .B1(new_n276), .B2(new_n274), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(KEYINPUT65), .ZN(new_n302));
  XNOR2_X1  g116(.A(G116), .B(G119), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT2), .B(G113), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n300), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n276), .A2(new_n297), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT64), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT64), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n276), .A2(new_n297), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n294), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n277), .A2(new_n286), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n305), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n266), .B1(new_n307), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n299), .A2(new_n313), .A3(new_n305), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n265), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n301), .A2(KEYINPUT65), .B1(new_n298), .B2(new_n294), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n312), .A2(new_n320), .A3(new_n313), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n306), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n305), .A3(new_n323), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n264), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT30), .B1(new_n300), .B2(new_n302), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n325), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n307), .B1(new_n333), .B2(new_n306), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT31), .A3(new_n264), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n319), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(G472), .A2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT32), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n319), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT31), .B1(new_n334), .B2(new_n264), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n305), .B1(new_n332), .B2(new_n325), .ZN(new_n342));
  INV_X1    g156(.A(new_n264), .ZN(new_n343));
  NOR4_X1   g157(.A1(new_n342), .A2(new_n330), .A3(new_n307), .A4(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n340), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n337), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n306), .B1(new_n300), .B2(new_n302), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n328), .A3(KEYINPUT68), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n351), .B(new_n306), .C1(new_n300), .C2(new_n302), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(KEYINPUT28), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT29), .A3(new_n318), .A4(new_n264), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n315), .A2(new_n318), .A3(new_n265), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n334), .A2(new_n264), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n188), .B(new_n354), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G472), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n259), .B1(new_n348), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G469), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(new_n364), .B2(G107), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G104), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n364), .A2(G107), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G101), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(KEYINPUT4), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(new_n285), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n370), .A2(G101), .ZN(new_n374));
  AOI21_X1  g188(.A(G101), .B1(new_n364), .B2(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n365), .A2(new_n375), .A3(new_n368), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT4), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n374), .A2(new_n377), .A3(KEYINPUT73), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT73), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n376), .A2(KEYINPUT4), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n371), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n373), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n277), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n288), .B2(new_n290), .ZN(new_n385));
  OAI211_X1 g199(.A(KEYINPUT75), .B(new_n289), .C1(new_n283), .C2(G128), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n293), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n365), .A2(new_n375), .A3(new_n368), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT74), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(new_n367), .B2(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n367), .A2(G104), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n364), .A2(KEYINPUT74), .A3(G107), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n388), .B1(G101), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT10), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(G101), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n398), .A2(KEYINPUT76), .A3(new_n376), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT76), .B1(new_n398), .B2(new_n376), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT10), .B(new_n294), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n382), .A2(new_n383), .A3(new_n397), .A4(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G140), .ZN(new_n403));
  INV_X1    g217(.A(G227), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G953), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n409));
  INV_X1    g223(.A(G101), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT74), .B1(new_n364), .B2(G107), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n364), .A2(G107), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n410), .B1(new_n413), .B2(new_n392), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n409), .B1(new_n414), .B2(new_n388), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n283), .A2(new_n292), .A3(G128), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n289), .B1(new_n283), .B2(G128), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n398), .A2(KEYINPUT76), .A3(new_n376), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n415), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n395), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT12), .A3(new_n277), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n277), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT12), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n408), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n382), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n397), .A2(new_n401), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n277), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n407), .B1(new_n429), .B2(new_n402), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n363), .B(new_n188), .C1(new_n426), .C2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT12), .B1(new_n421), .B2(new_n277), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n424), .B(new_n383), .C1(new_n420), .C2(new_n395), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n402), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n406), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n402), .A2(new_n407), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n429), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(G469), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n363), .A2(new_n188), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n431), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT9), .B(G234), .ZN(new_n443));
  OAI21_X1  g257(.A(G221), .B1(new_n443), .B2(G902), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT77), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n207), .B1(new_n416), .B2(new_n417), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n282), .B(G125), .C1(new_n283), .C2(new_n284), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G224), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n451), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G122), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT78), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT2), .B(G113), .Z(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n303), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n191), .A2(G116), .ZN(new_n460));
  INV_X1    g274(.A(G116), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G119), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(new_n304), .ZN(new_n464));
  OAI22_X1  g278(.A1(KEYINPUT4), .A2(new_n371), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT73), .B1(new_n374), .B2(new_n377), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n380), .A2(new_n379), .A3(new_n371), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G113), .B1(new_n460), .B2(KEYINPUT5), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n464), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n415), .B2(new_n419), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n457), .B1(new_n468), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n456), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n468), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT6), .B(new_n457), .C1(new_n468), .C2(new_n475), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n455), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n456), .B(KEYINPUT8), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n469), .A2(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n471), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n469), .A2(KEYINPUT79), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n473), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n415), .B2(new_n419), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n394), .B1(new_n473), .B2(new_n472), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n483), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n372), .A2(new_n305), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n378), .B2(new_n381), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n473), .B(new_n472), .C1(new_n399), .C2(new_n400), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(new_n456), .ZN(new_n494));
  INV_X1    g308(.A(new_n453), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT80), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n449), .A2(new_n450), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(KEYINPUT7), .A3(new_n495), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(KEYINPUT7), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n449), .A2(new_n450), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n490), .A2(new_n494), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n188), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n448), .B1(new_n482), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n492), .A2(new_n493), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n494), .A2(KEYINPUT6), .B1(new_n504), .B2(new_n457), .ZN(new_n505));
  INV_X1    g319(.A(new_n481), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n454), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n498), .A2(new_n500), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n478), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n509), .B2(new_n490), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n510), .A3(new_n447), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n503), .A2(KEYINPUT81), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G214), .B1(G237), .B2(G902), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n447), .B1(new_n507), .B2(new_n510), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT81), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n518));
  NOR2_X1   g332(.A1(G475), .A2(G902), .ZN(new_n519));
  INV_X1    g333(.A(G237), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n217), .A3(G214), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n279), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n275), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT82), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n526));
  INV_X1    g340(.A(new_n523), .ZN(new_n527));
  AOI21_X1  g341(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n528));
  OAI21_X1  g342(.A(G131), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT82), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n522), .A2(new_n530), .A3(new_n275), .A4(new_n523), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n525), .A2(new_n526), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n234), .A2(new_n235), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n529), .A2(new_n526), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G113), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(new_n364), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n206), .A2(new_n208), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G146), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n214), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT18), .B(G131), .C1(new_n527), .C2(new_n528), .ZN(new_n541));
  NAND2_X1  g355(.A1(KEYINPUT18), .A2(G131), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n522), .A2(new_n523), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n535), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n525), .A2(new_n529), .A3(new_n531), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT19), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT19), .B1(new_n206), .B2(new_n208), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n213), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n211), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n537), .B1(new_n551), .B2(new_n544), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n519), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n544), .ZN(new_n554));
  INV_X1    g368(.A(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT83), .B1(new_n556), .B2(new_n545), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n557), .B2(KEYINPUT20), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n545), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT20), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(KEYINPUT83), .A3(new_n560), .A4(new_n519), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n537), .B1(new_n535), .B2(new_n544), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n188), .B1(new_n546), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT84), .B(G475), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n279), .A2(KEYINPUT13), .A3(G128), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT86), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n279), .A2(G128), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT13), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT86), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n573), .A2(new_n279), .A3(KEYINPUT13), .A4(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n220), .A2(G143), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n569), .A2(new_n572), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G134), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n575), .A3(new_n268), .ZN(new_n578));
  INV_X1    g392(.A(G122), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT85), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT85), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G122), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G116), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n461), .A2(G122), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n367), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n461), .B1(new_n580), .B2(new_n582), .ZN(new_n587));
  INV_X1    g401(.A(new_n585), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n587), .A2(G107), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n577), .B(new_n578), .C1(new_n586), .C2(new_n589), .ZN(new_n590));
  OR3_X1    g404(.A1(new_n579), .A2(KEYINPUT14), .A3(G116), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n585), .A2(KEYINPUT14), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G107), .B1(new_n593), .B2(new_n587), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n584), .A2(new_n367), .A3(new_n585), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n570), .A2(new_n575), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G134), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n578), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n443), .A2(new_n187), .A3(G953), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n590), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n590), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n188), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT87), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n590), .A2(new_n599), .ZN(new_n606));
  INV_X1    g420(.A(new_n600), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n590), .A2(new_n599), .A3(new_n600), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(KEYINPUT87), .A3(new_n188), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G478), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(KEYINPUT15), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n217), .A2(G952), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(G234), .B2(G237), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n188), .B(new_n217), .C1(G234), .C2(G237), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT21), .B(G898), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n614), .B1(new_n603), .B2(new_n604), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n615), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n518), .B1(new_n567), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n614), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n605), .B2(new_n611), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n627), .A2(new_n620), .A3(new_n622), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n558), .A2(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT88), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT77), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n442), .A2(new_n632), .A3(new_n444), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n446), .A2(new_n517), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n362), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n410), .ZN(G3));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n345), .B2(new_n188), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n336), .A2(new_n338), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n638), .A2(new_n639), .A3(new_n259), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n640), .A2(new_n446), .A3(new_n633), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n603), .A2(new_n613), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT33), .B1(new_n608), .B2(new_n609), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n643), .A2(KEYINPUT89), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(KEYINPUT89), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n609), .A2(KEYINPUT90), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n609), .A2(KEYINPUT90), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n646), .A2(KEYINPUT33), .A3(new_n608), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n188), .A2(G478), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n642), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n567), .A3(new_n621), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n482), .A2(new_n502), .A3(new_n448), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n513), .B1(new_n653), .B2(new_n514), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n641), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT91), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT34), .B(G104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  NOR2_X1   g473(.A1(new_n627), .A2(new_n622), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n559), .A2(new_n560), .A3(new_n519), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n662), .A2(new_n663), .B1(new_n564), .B2(new_n565), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n661), .A2(new_n621), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n654), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n641), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n246), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(new_n245), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n257), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n256), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT92), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n256), .A2(KEYINPUT92), .A3(new_n673), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n638), .A2(new_n639), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n634), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT93), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G12));
  AOI22_X1  g498(.A1(new_n348), .A2(new_n360), .B1(new_n676), .B2(new_n677), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n442), .A2(new_n632), .A3(new_n444), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n632), .B1(new_n442), .B2(new_n444), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n513), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n503), .B2(new_n511), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n617), .B(KEYINPUT94), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(G900), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n692), .B1(new_n693), .B2(new_n618), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n661), .A2(new_n664), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n685), .A2(new_n688), .A3(new_n690), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  XOR2_X1   g512(.A(new_n694), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n688), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT97), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(KEYINPUT97), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n701), .B2(new_n703), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n629), .A2(new_n660), .A3(new_n689), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n676), .A2(new_n677), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT96), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n512), .A2(new_n516), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n350), .A2(new_n352), .ZN(new_n712));
  INV_X1    g526(.A(new_n265), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n712), .A2(new_n713), .B1(new_n334), .B2(new_n264), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n714), .B2(G902), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n348), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n708), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n704), .A2(new_n705), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n279), .ZN(G45));
  NAND2_X1  g535(.A1(new_n685), .A2(new_n688), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n651), .A2(new_n567), .A3(new_n695), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n723), .A2(new_n654), .A3(KEYINPUT98), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT98), .B1(new_n723), .B2(new_n654), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  NAND2_X1  g542(.A1(new_n429), .A2(new_n402), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n425), .A2(new_n422), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n406), .A2(new_n729), .B1(new_n730), .B2(new_n437), .ZN(new_n731));
  OAI21_X1  g545(.A(G469), .B1(new_n731), .B2(G902), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n444), .A3(new_n431), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n361), .A2(new_n655), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND2_X1  g551(.A1(new_n348), .A2(new_n360), .ZN(new_n738));
  INV_X1    g552(.A(new_n259), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n739), .A3(new_n666), .A4(new_n734), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  NOR2_X1   g555(.A1(new_n733), .A2(new_n654), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n738), .A2(new_n631), .A3(new_n678), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  NAND2_X1  g558(.A1(new_n503), .A2(new_n511), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n706), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n732), .A2(new_n444), .A3(new_n431), .A4(new_n621), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n331), .A2(new_n335), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n353), .A2(new_n318), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n713), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n338), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n638), .A2(new_n259), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  INV_X1    g569(.A(new_n723), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n638), .A2(new_n752), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n678), .A2(new_n742), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT99), .B(G125), .Z(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G27));
  AOI21_X1  g574(.A(new_n689), .B1(new_n512), .B2(new_n516), .ZN(new_n761));
  INV_X1    g575(.A(new_n444), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n415), .A2(new_n419), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n418), .A2(new_n396), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n763), .A2(new_n764), .B1(new_n395), .B2(new_n396), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n383), .B1(new_n765), .B2(new_n382), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n406), .B1(new_n435), .B2(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n407), .B(new_n402), .C1(new_n432), .C2(new_n433), .ZN(new_n768));
  AOI21_X1  g582(.A(G902), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n440), .B1(new_n769), .B2(new_n363), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n762), .B1(new_n770), .B2(new_n439), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n761), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT100), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(KEYINPUT42), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n361), .A3(new_n756), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n761), .A2(new_n771), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n339), .A2(new_n347), .B1(G472), .B2(new_n359), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n777), .A2(new_n778), .A3(new_n259), .A4(new_n723), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NAND3_X1  g596(.A1(new_n772), .A2(new_n361), .A3(new_n696), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  AND2_X1   g598(.A1(new_n436), .A2(new_n438), .ZN(new_n785));
  OAI21_X1  g599(.A(G469), .B1(new_n785), .B2(KEYINPUT45), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT101), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n786), .A2(KEYINPUT101), .B1(KEYINPUT45), .B2(new_n785), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n440), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(KEYINPUT46), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n431), .B1(new_n789), .B2(KEYINPUT46), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n444), .B(new_n699), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n761), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n651), .A2(new_n629), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n679), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n797), .A3(new_n678), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n793), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n792), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g616(.A(KEYINPUT102), .B(G137), .Z(new_n803));
  XNOR2_X1  g617(.A(new_n802), .B(new_n803), .ZN(G39));
  NOR4_X1   g618(.A1(new_n738), .A2(new_n793), .A3(new_n739), .A4(new_n723), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT103), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n444), .B1(new_n790), .B2(new_n791), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n205), .ZN(G42));
  NOR2_X1   g627(.A1(new_n769), .A2(new_n363), .ZN(new_n814));
  AOI211_X1 g628(.A(G469), .B(G902), .C1(new_n767), .C2(new_n768), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT49), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n794), .A2(new_n259), .A3(new_n762), .A4(new_n689), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n711), .A2(new_n717), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n735), .A2(new_n740), .A3(new_n743), .A4(new_n754), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT104), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT88), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT88), .B1(new_n628), .B2(new_n629), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(new_n444), .A3(new_n690), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n826), .A2(new_n685), .B1(new_n748), .B2(new_n753), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT104), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n735), .A4(new_n740), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n821), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n678), .A2(new_n757), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT107), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n756), .A4(new_n772), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n678), .A2(new_n756), .A3(new_n757), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT107), .B1(new_n834), .B2(new_n777), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n664), .A2(new_n660), .A3(new_n695), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n689), .B(new_n837), .C1(new_n516), .C2(new_n512), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n685), .A2(new_n688), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(new_n783), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n781), .A2(new_n836), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n830), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n661), .A2(new_n629), .A3(new_n621), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n446), .A3(new_n640), .A4(new_n633), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n634), .B2(new_n680), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n843), .A2(new_n652), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n446), .A3(new_n640), .A4(new_n633), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n362), .B2(new_n634), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n847), .B1(KEYINPUT105), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT105), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n849), .B(new_n852), .C1(new_n362), .C2(new_n634), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT106), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n850), .A2(KEYINPUT105), .ZN(new_n855));
  INV_X1    g669(.A(new_n847), .ZN(new_n856));
  AND4_X1   g670(.A1(KEYINPUT106), .A2(new_n855), .A3(new_n853), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n842), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT108), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n842), .B(KEYINPUT108), .C1(new_n854), .C2(new_n857), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n445), .A2(new_n674), .A3(new_n694), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n716), .A3(new_n745), .A4(new_n706), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n727), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n697), .A2(new_n758), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(KEYINPUT52), .B(new_n864), .C1(new_n722), .C2(new_n726), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n860), .A2(new_n861), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT53), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  INV_X1    g686(.A(new_n868), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n697), .A2(KEYINPUT109), .A3(new_n758), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT109), .B1(new_n697), .B2(new_n758), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT110), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT110), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n873), .B(new_n879), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n867), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n860), .A2(new_n872), .A3(new_n861), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n871), .A2(KEYINPUT54), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n870), .A2(new_n872), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n854), .A2(new_n857), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n820), .B(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n888), .A2(new_n872), .A3(new_n841), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n881), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n885), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n883), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n883), .B2(new_n892), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n816), .A2(new_n762), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n810), .A2(new_n811), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n796), .A2(new_n692), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n898), .A2(new_n753), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n761), .A3(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n689), .A3(new_n711), .A4(new_n734), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT50), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n793), .A2(new_n733), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n739), .A2(new_n617), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n904), .A2(new_n717), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n651), .A2(new_n567), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n904), .ZN(new_n909));
  INV_X1    g723(.A(new_n831), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n907), .A2(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n900), .A2(new_n903), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n909), .A2(new_n362), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT48), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n899), .A2(new_n742), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n616), .B(KEYINPUT115), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n651), .A2(new_n567), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n918), .B(new_n919), .C1(new_n920), .C2(new_n907), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n912), .A2(KEYINPUT113), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n912), .A2(KEYINPUT113), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n903), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT114), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n900), .A2(KEYINPUT51), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n915), .B(new_n922), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n894), .A2(new_n895), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(G952), .A2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n819), .B1(new_n930), .B2(new_n931), .ZN(G75));
  AOI21_X1  g746(.A(new_n890), .B1(new_n870), .B2(new_n872), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n188), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT116), .B1(new_n934), .B2(G210), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT116), .ZN(new_n936));
  INV_X1    g750(.A(G210), .ZN(new_n937));
  NOR4_X1   g751(.A1(new_n933), .A2(new_n936), .A3(new_n937), .A4(new_n188), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n505), .A2(new_n506), .A3(new_n454), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n482), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT55), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n935), .A2(new_n938), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n217), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT56), .B1(new_n934), .B2(G210), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n944), .A2(new_n948), .ZN(G51));
  XNOR2_X1  g763(.A(new_n440), .B(KEYINPUT57), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n933), .A2(new_n885), .ZN(new_n951));
  AOI211_X1 g765(.A(KEYINPUT54), .B(new_n890), .C1(new_n872), .C2(new_n870), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n731), .B(KEYINPUT117), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n934), .A2(new_n787), .A3(new_n788), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n945), .B1(new_n955), .B2(new_n956), .ZN(G54));
  NAND3_X1  g771(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n958));
  INV_X1    g772(.A(new_n559), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n961), .A3(new_n945), .ZN(G60));
  NAND2_X1  g776(.A1(G478), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT59), .Z(new_n964));
  NOR2_X1   g778(.A1(new_n649), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n951), .B2(new_n952), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n946), .ZN(new_n967));
  INV_X1    g781(.A(new_n964), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n894), .B2(new_n895), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n967), .B1(new_n969), .B2(new_n649), .ZN(G63));
  INV_X1    g784(.A(new_n933), .ZN(new_n971));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT60), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n971), .A2(new_n672), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n247), .B(new_n250), .C1(new_n933), .C2(new_n973), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n975), .A2(new_n946), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT61), .A4(new_n946), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(G66));
  OAI21_X1  g795(.A(G953), .B1(new_n619), .B2(new_n452), .ZN(new_n982));
  INV_X1    g796(.A(new_n830), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n886), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n480), .B(new_n481), .C1(G898), .C2(new_n217), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  OAI21_X1  g802(.A(G953), .B1(new_n404), .B2(new_n693), .ZN(new_n989));
  XNOR2_X1  g803(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n333), .B(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT120), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n548), .A2(new_n549), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n989), .B1(new_n995), .B2(KEYINPUT124), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n727), .B1(new_n875), .B2(new_n876), .ZN(new_n998));
  OR3_X1    g812(.A1(new_n720), .A2(KEYINPUT62), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n661), .A2(new_n629), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n793), .B1(new_n920), .B2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n701), .A2(new_n361), .A3(new_n703), .A4(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n792), .B2(new_n801), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT121), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n812), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT62), .B1(new_n720), .B2(new_n998), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n999), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n995), .B1(new_n1008), .B2(new_n217), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n792), .A2(new_n362), .A3(new_n746), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n781), .A2(new_n783), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n812), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OR3_X1    g827(.A1(new_n802), .A2(new_n998), .A3(KEYINPUT122), .ZN(new_n1014));
  OAI21_X1  g828(.A(KEYINPUT122), .B1(new_n802), .B2(new_n998), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(G953), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT123), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n217), .A2(G900), .ZN(new_n1019));
  OR3_X1    g833(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1018), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n997), .B(new_n1010), .C1(new_n1022), .C2(new_n994), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n994), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n996), .B1(new_n1024), .B2(new_n1009), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(G72));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT63), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT125), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(new_n984), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n334), .B(KEYINPUT126), .Z(new_n1032));
  NOR2_X1   g846(.A1(new_n1032), .A2(new_n264), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n945), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1029), .B1(new_n1008), .B2(new_n984), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(new_n264), .A3(new_n1032), .ZN(new_n1036));
  INV_X1    g850(.A(new_n358), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1028), .B1(new_n1037), .B2(new_n329), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n871), .A2(new_n882), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1034), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT127), .ZN(G57));
endmodule


