//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(G8gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n203), .B2(new_n206), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT83), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(new_n207), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT17), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n228), .B1(new_n224), .B2(new_n225), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n210), .B(new_n213), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(KEYINPUT84), .Z(new_n232));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n208), .A2(new_n233), .A3(new_n209), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n208), .B2(new_n209), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n226), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n230), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n232), .A4(new_n237), .ZN(new_n241));
  INV_X1    g040(.A(new_n236), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n224), .B(new_n225), .C1(new_n242), .C2(new_n234), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n237), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n232), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(G169gat), .B(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT12), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n238), .A2(new_n239), .B1(new_n244), .B2(new_n245), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n253), .B1(new_n256), .B2(new_n241), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(G169gat), .A3(G176gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT26), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n264), .A2(KEYINPUT68), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT68), .B1(new_n264), .B2(new_n267), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n263), .B(new_n266), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G183gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT27), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n276), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n272), .A2(new_n274), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n275), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n270), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G169gat), .B2(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n264), .A2(KEYINPUT23), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n261), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT24), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n289), .A2(new_n291), .B1(new_n271), .B2(new_n275), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT25), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n291), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G183gat), .B2(G190gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n271), .A2(new_n275), .A3(KEYINPUT65), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n282), .A2(G169gat), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT25), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n282), .A2(new_n265), .B1(new_n260), .B2(new_n262), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n281), .A2(new_n293), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n281), .A2(new_n308), .A3(new_n293), .A4(new_n305), .ZN(new_n309));
  AND2_X1   g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(KEYINPUT29), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n293), .A2(new_n305), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(new_n310), .A3(new_n281), .ZN(new_n314));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(G211gat), .ZN(new_n316));
  INV_X1    g115(.A(G218gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(KEYINPUT22), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(new_n314), .A3(new_n321), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n306), .A2(new_n311), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n309), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n310), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT74), .B(new_n322), .C1(new_n325), .C2(new_n321), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n312), .A2(new_n314), .A3(new_n327), .A4(new_n321), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G1gat), .B(G29gat), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT0), .ZN(new_n335));
  XNOR2_X1  g134(.A(G57gat), .B(G85gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n338));
  XOR2_X1   g137(.A(G141gat), .B(G148gat), .Z(new_n339));
  INV_X1    g138(.A(G155gat), .ZN(new_n340));
  INV_X1    g139(.A(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(KEYINPUT2), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G141gat), .B(G148gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n343), .B(new_n342), .C1(new_n347), .C2(KEYINPUT2), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G113gat), .A2(G120gat), .ZN(new_n350));
  INV_X1    g149(.A(G113gat), .ZN(new_n351));
  INV_X1    g150(.A(G120gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT1), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n350), .B(new_n353), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n352), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n350), .ZN(new_n359));
  INV_X1    g158(.A(G134gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G127gat), .ZN(new_n361));
  INV_X1    g160(.A(G127gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n355), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n356), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n346), .A3(new_n356), .A4(new_n366), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n338), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT76), .B1(new_n369), .B2(KEYINPUT4), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n346), .A2(new_n348), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n367), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n346), .A2(new_n348), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n356), .A2(new_n366), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(new_n386), .A3(new_n371), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n373), .B1(new_n377), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(new_n371), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n382), .A2(new_n383), .A3(new_n376), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n369), .A2(new_n385), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(new_n338), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n337), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT6), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  INV_X1    g196(.A(new_n369), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n348), .A2(new_n346), .B1(new_n356), .B2(new_n366), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n372), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n381), .A2(new_n386), .A3(new_n371), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n369), .A2(new_n376), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n403), .B(KEYINPUT76), .C1(KEYINPUT4), .C2(new_n369), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n337), .B1(new_n389), .B2(new_n392), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n397), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT79), .B1(new_n407), .B2(new_n395), .ZN(new_n408));
  INV_X1    g207(.A(new_n337), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n405), .B2(new_n393), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n381), .A2(new_n371), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n390), .A2(new_n338), .A3(new_n391), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT6), .B1(new_n388), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n333), .A2(new_n396), .A3(new_n408), .A4(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n332), .A2(KEYINPUT38), .ZN(new_n418));
  INV_X1    g217(.A(new_n321), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n325), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n312), .A2(new_n314), .A3(new_n419), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT37), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT37), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(new_n329), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT80), .B1(new_n417), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n408), .A2(new_n396), .A3(new_n416), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n329), .A2(new_n424), .ZN(new_n429));
  INV_X1    g228(.A(new_n423), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n427), .A2(new_n428), .A3(new_n431), .A4(new_n333), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n326), .A2(KEYINPUT37), .A3(new_n328), .ZN(new_n433));
  INV_X1    g232(.A(new_n332), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT38), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n426), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n380), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n321), .B1(new_n438), .B2(KEYINPUT29), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT3), .B1(new_n419), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n441), .B2(new_n382), .ZN(new_n442));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g243(.A(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G22gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT31), .B(G50gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  MUX2_X1   g248(.A(G22gat), .B(new_n446), .S(new_n449), .Z(new_n450));
  XNOR2_X1  g249(.A(new_n444), .B(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n326), .A2(new_n328), .A3(new_n434), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT30), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n434), .B1(new_n326), .B2(new_n328), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI211_X1 g254(.A(KEYINPUT30), .B(new_n434), .C1(new_n326), .C2(new_n328), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n381), .A2(new_n390), .A3(new_n391), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n459), .A2(KEYINPUT78), .A3(new_n372), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT78), .B1(new_n459), .B2(new_n372), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n372), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(KEYINPUT78), .A3(new_n372), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n370), .A2(new_n372), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(new_n458), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n462), .A2(new_n469), .A3(KEYINPUT40), .A4(new_n337), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n470), .A2(new_n410), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n462), .A2(new_n469), .A3(new_n337), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n451), .B1(new_n457), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n437), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n313), .A2(KEYINPUT70), .A3(new_n383), .A4(new_n281), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n281), .A2(new_n383), .A3(new_n293), .A4(new_n305), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n306), .A2(new_n367), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT64), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT72), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT32), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n483), .B2(new_n485), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT33), .B1(new_n483), .B2(new_n485), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G43gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G71gat), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n496));
  INV_X1    g295(.A(G71gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n495), .A2(new_n499), .A3(G99gat), .ZN(new_n500));
  AOI21_X1  g299(.A(G99gat), .B1(new_n495), .B2(new_n499), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n491), .A2(new_n492), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n487), .A2(KEYINPUT72), .ZN(new_n505));
  AOI221_X4 g304(.A(new_n490), .B1(new_n502), .B2(KEYINPUT33), .C1(new_n483), .C2(new_n485), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n505), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n483), .A2(new_n485), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT32), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT33), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n512), .A3(new_n502), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n491), .B1(new_n492), .B2(new_n503), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n489), .B1(new_n507), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n517));
  INV_X1    g316(.A(new_n489), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(new_n508), .A3(new_n514), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n516), .A2(KEYINPUT36), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT36), .B1(new_n516), .B2(new_n520), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n407), .A2(new_n395), .ZN(new_n524));
  AOI211_X1 g323(.A(new_n397), .B(new_n337), .C1(new_n388), .C2(new_n394), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n455), .B2(new_n456), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n451), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n477), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n451), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n518), .B1(new_n517), .B2(new_n519), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT35), .B1(new_n534), .B2(new_n528), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n451), .B1(new_n516), .B2(new_n520), .ZN(new_n536));
  INV_X1    g335(.A(new_n427), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n333), .A2(KEYINPUT30), .A3(new_n452), .ZN(new_n538));
  INV_X1    g337(.A(new_n456), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT81), .B(KEYINPUT35), .Z(new_n541));
  NAND4_X1  g340(.A1(new_n536), .A2(new_n537), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n258), .B1(new_n530), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n545));
  NOR2_X1   g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(G71gat), .B2(G78gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT86), .B1(G71gat), .B2(G78gat), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n547), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G64gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(G57gat), .ZN(new_n556));
  INV_X1    g355(.A(G57gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G64gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT9), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n556), .A2(new_n558), .B1(new_n559), .B2(new_n550), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n545), .B1(new_n554), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n547), .A2(new_n549), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n558), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n550), .A2(new_n559), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n550), .B(new_n551), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT88), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT89), .B(G57gat), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT90), .B(new_n556), .C1(new_n569), .C2(new_n555), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n546), .A2(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n550), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n569), .A2(new_n555), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n570), .B(new_n572), .C1(new_n573), .C2(KEYINPUT90), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT21), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G127gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n568), .A2(new_n574), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT91), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n580), .A2(KEYINPUT21), .B1(new_n235), .B2(new_n236), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n578), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G155gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(G85gat), .ZN(new_n593));
  INV_X1    g392(.A(G92gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G99gat), .B(G106gat), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n591), .A3(new_n595), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n227), .B2(new_n229), .ZN(new_n602));
  INV_X1    g401(.A(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT92), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n226), .A2(new_n603), .B1(KEYINPUT41), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n612));
  XOR2_X1   g411(.A(G190gat), .B(G218gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT93), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n611), .B(new_n615), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n589), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n601), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n580), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n598), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n596), .A2(KEYINPUT95), .A3(new_n597), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n568), .A3(new_n574), .A4(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n579), .A2(KEYINPUT94), .A3(new_n601), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT94), .B1(new_n579), .B2(new_n601), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n620), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n619), .B1(new_n622), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  OAI21_X1  g433(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n619), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n631), .A2(KEYINPUT96), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n634), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n639), .B2(new_n630), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n618), .B(KEYINPUT97), .Z(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n622), .B2(new_n629), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n636), .ZN(new_n645));
  INV_X1    g444(.A(new_n634), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n617), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n544), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n527), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT98), .B(G1gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1324gat));
  NOR2_X1   g452(.A1(new_n650), .A2(new_n540), .ZN(new_n654));
  NAND2_X1  g453(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n205), .A2(new_n204), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n204), .B2(new_n654), .ZN(new_n658));
  MUX2_X1   g457(.A(new_n657), .B(new_n658), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n532), .A2(new_n533), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n650), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT99), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n650), .A2(new_n660), .A3(new_n523), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n531), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT100), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR3_X1   g468(.A1(new_n589), .A2(new_n616), .A3(new_n648), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n544), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n218), .A3(new_n526), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n616), .B1(new_n530), .B2(new_n543), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n247), .A2(new_n254), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n256), .A2(new_n241), .A3(new_n253), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n680), .A2(KEYINPUT101), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT101), .B1(new_n680), .B2(new_n681), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(new_n589), .A3(new_n648), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(new_n526), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n674), .B1(new_n688), .B2(new_n218), .ZN(G1328gat));
  NOR3_X1   g488(.A1(new_n671), .A2(G36gat), .A3(new_n540), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT46), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n687), .A2(new_n457), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n692), .B2(new_n214), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1329gat));
  NOR3_X1   g494(.A1(new_n671), .A2(G43gat), .A3(new_n661), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n523), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n698), .A3(new_n686), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT105), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G43gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n699), .A2(KEYINPUT105), .ZN(new_n702));
  OAI211_X1 g501(.A(KEYINPUT47), .B(new_n697), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(G43gat), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT47), .B1(new_n704), .B2(new_n697), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n705), .A2(KEYINPUT104), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(KEYINPUT104), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(G1330gat));
  NOR3_X1   g507(.A1(new_n671), .A2(G50gat), .A3(new_n531), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n687), .A2(new_n451), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(G50gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g511(.A1(new_n471), .A2(new_n474), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n531), .B1(new_n540), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n525), .B1(new_n524), .B2(new_n415), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n431), .A2(new_n715), .A3(new_n333), .A4(new_n408), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n716), .A2(KEYINPUT80), .B1(KEYINPUT38), .B2(new_n435), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n714), .B1(new_n717), .B2(new_n432), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT36), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n532), .B2(new_n533), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n516), .A2(KEYINPUT36), .A3(new_n520), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n529), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT35), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n526), .B1(new_n538), .B2(new_n539), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n536), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n540), .A2(new_n537), .A3(new_n541), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n534), .A2(new_n726), .ZN(new_n727));
  OAI22_X1  g526(.A1(new_n718), .A2(new_n722), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n637), .A2(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n617), .A2(new_n729), .A3(new_n684), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n526), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(new_n569), .ZN(G1332gat));
  AOI21_X1  g532(.A(new_n540), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT108), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n735), .B(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1333gat));
  AOI21_X1  g539(.A(new_n497), .B1(new_n731), .B2(new_n698), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n661), .A2(G71gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n731), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n731), .A2(new_n451), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n589), .A2(new_n684), .ZN(new_n748));
  INV_X1    g547(.A(new_n616), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n728), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n750), .B2(KEYINPUT110), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n675), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n747), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(KEYINPUT110), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n675), .A2(new_n752), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT51), .A4(new_n748), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n729), .A2(G85gat), .A3(new_n527), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT111), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n589), .A2(new_n729), .A3(new_n684), .ZN(new_n762));
  INV_X1    g561(.A(new_n676), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n616), .B(new_n763), .C1(new_n530), .C2(new_n543), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n678), .B1(new_n728), .B2(new_n749), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT109), .B(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n526), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n761), .B1(new_n771), .B2(new_n593), .ZN(G1336gat));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  OAI21_X1  g572(.A(G92gat), .B1(new_n766), .B2(new_n540), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n729), .B1(new_n754), .B2(new_n757), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n457), .A2(new_n594), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n773), .B(new_n774), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n768), .A2(new_n457), .A3(new_n769), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n779), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT112), .B1(new_n779), .B2(G92gat), .ZN(new_n781));
  AOI211_X1 g580(.A(new_n729), .B(new_n777), .C1(new_n754), .C2(new_n757), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(new_n783), .B2(new_n773), .ZN(G1337gat));
  NAND2_X1  g583(.A1(new_n770), .A2(new_n698), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G99gat), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n661), .A2(G99gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n776), .B2(new_n787), .ZN(G1338gat));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT113), .B(G106gat), .Z(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n768), .A2(new_n451), .A3(new_n769), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n531), .A2(G106gat), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n791), .A2(new_n792), .B1(new_n775), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n775), .A2(new_n793), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n791), .B1(new_n766), .B2(new_n531), .ZN(new_n798));
  XOR2_X1   g597(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n797), .A2(KEYINPUT116), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802));
  INV_X1    g601(.A(new_n793), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n729), .B(new_n803), .C1(new_n754), .C2(new_n757), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n800), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n792), .A2(new_n791), .ZN(new_n808));
  OAI211_X1 g607(.A(KEYINPUT114), .B(KEYINPUT53), .C1(new_n808), .C2(new_n804), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n796), .A2(new_n807), .A3(new_n809), .ZN(G1339gat));
  INV_X1    g609(.A(new_n589), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n622), .A2(new_n629), .ZN(new_n813));
  INV_X1    g612(.A(new_n642), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n622), .A2(new_n629), .A3(KEYINPUT117), .A4(new_n642), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n815), .A2(KEYINPUT54), .A3(new_n631), .A4(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  AOI211_X1 g618(.A(new_n818), .B(new_n634), .C1(new_n643), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n641), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n634), .B1(new_n643), .B2(new_n819), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT55), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT118), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n817), .A2(new_n823), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n818), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n817), .A2(new_n820), .B1(new_n637), .B2(new_n640), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n825), .A2(new_n684), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n244), .A2(new_n245), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n232), .B1(new_n230), .B2(new_n237), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n252), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n681), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT119), .B1(new_n648), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n729), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n749), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n616), .A2(new_n835), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n825), .A2(new_n842), .A3(new_n830), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n811), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n649), .A2(new_n685), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n527), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n540), .A3(new_n536), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n684), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n451), .B1(new_n844), .B2(new_n845), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n540), .A2(new_n526), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n661), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n258), .A2(new_n351), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(G1340gat));
  AOI21_X1  g654(.A(G120gat), .B1(new_n848), .B2(new_n648), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n729), .A2(new_n352), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(G1341gat));
  INV_X1    g657(.A(new_n853), .ZN(new_n859));
  OAI21_X1  g658(.A(G127gat), .B1(new_n859), .B2(new_n811), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n848), .A2(new_n362), .A3(new_n589), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1342gat));
  NAND3_X1  g661(.A1(new_n848), .A2(new_n360), .A3(new_n749), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n859), .B2(new_n616), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n698), .A2(new_n852), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n844), .A2(new_n845), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n869), .B2(new_n451), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n531), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n822), .A2(new_n258), .A3(new_n824), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n729), .A2(new_n835), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n616), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n811), .B1(new_n877), .B2(new_n843), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n873), .B1(new_n878), .B2(new_n845), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n868), .B1(new_n870), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n258), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n698), .A2(new_n531), .A3(new_n457), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n846), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(G141gat), .A3(new_n258), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(KEYINPUT58), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n684), .B(new_n868), .C1(new_n870), .C2(new_n879), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n887), .A2(KEYINPUT120), .A3(G141gat), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT120), .B1(new_n887), .B2(G141gat), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(new_n884), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(G1344gat));
  AOI21_X1  g691(.A(new_n873), .B1(new_n844), .B2(new_n845), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n842), .A2(new_n827), .A3(new_n829), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n589), .B1(new_n876), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n258), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n617), .A2(new_n897), .A3(new_n648), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n451), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n871), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n901), .A2(new_n648), .A3(new_n868), .ZN(new_n902));
  INV_X1    g701(.A(G148gat), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT59), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(KEYINPUT59), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n880), .B2(new_n729), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n883), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n903), .A3(new_n648), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1345gat));
  OAI21_X1  g709(.A(G155gat), .B1(new_n880), .B2(new_n811), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n340), .A3(new_n589), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n880), .B2(new_n616), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n908), .A2(new_n341), .A3(new_n749), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1347gat));
  AOI21_X1  g715(.A(new_n526), .B1(new_n844), .B2(new_n845), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n534), .A2(new_n540), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n919), .A2(G169gat), .A3(new_n685), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n457), .A2(new_n527), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n661), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n850), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n258), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n921), .B1(new_n922), .B2(new_n926), .ZN(G1348gat));
  INV_X1    g726(.A(new_n919), .ZN(new_n928));
  AOI21_X1  g727(.A(G176gat), .B1(new_n928), .B2(new_n648), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n925), .A2(new_n301), .A3(new_n729), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(G1349gat));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n589), .A2(new_n278), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n850), .A2(new_n589), .A3(new_n924), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G183gat), .ZN(new_n936));
  XNOR2_X1  g735(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n937));
  AND4_X1   g736(.A1(new_n932), .A2(new_n934), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n934), .A2(new_n936), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n932), .B1(new_n939), .B2(new_n937), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n275), .A3(new_n749), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  OAI21_X1  g744(.A(G190gat), .B1(new_n925), .B2(new_n616), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(G1351gat));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951));
  INV_X1    g750(.A(new_n900), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n893), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n894), .A2(KEYINPUT126), .A3(new_n900), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n698), .A2(new_n923), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n953), .A2(new_n954), .A3(new_n897), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G197gat), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n523), .A2(new_n451), .A3(new_n457), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT125), .Z(new_n959));
  NAND2_X1  g758(.A1(new_n917), .A2(new_n959), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n960), .A2(G197gat), .A3(new_n685), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n957), .A2(new_n964), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1352gat));
  AND3_X1   g765(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(new_n648), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G204gat), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n960), .A2(G204gat), .A3(new_n729), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n901), .A2(new_n589), .A3(new_n955), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n589), .A2(new_n316), .ZN(new_n976));
  OAI22_X1  g775(.A1(new_n974), .A2(new_n975), .B1(new_n960), .B2(new_n976), .ZN(G1354gat));
  NOR2_X1   g776(.A1(new_n616), .A2(new_n317), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n917), .A2(new_n749), .A3(new_n959), .ZN(new_n979));
  AOI22_X1  g778(.A1(new_n967), .A2(new_n978), .B1(new_n317), .B2(new_n979), .ZN(G1355gat));
endmodule


