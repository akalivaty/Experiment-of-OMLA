//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT79), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT65), .B1(new_n190), .B2(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n190), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  OAI21_X1  g012(.A(G128), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n202), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n200), .A2(KEYINPUT75), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G104), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n205), .A3(G104), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(G107), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n209), .B(new_n215), .C1(new_n203), .C2(KEYINPUT75), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n204), .A2(KEYINPUT76), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n218));
  INV_X1    g032(.A(new_n216), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n200), .A2(KEYINPUT75), .A3(new_n203), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n193), .A2(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n195), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n199), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n203), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n209), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n217), .A2(new_n221), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G137), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G131), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT12), .B1(new_n228), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n227), .A2(new_n225), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT76), .B1(new_n204), .B2(new_n216), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n219), .A2(new_n218), .A3(new_n220), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n243), .A2(new_n244), .A3(new_n237), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n189), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT10), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n217), .B2(new_n221), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n249), .B(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n223), .A2(new_n256), .A3(KEYINPUT64), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT64), .B1(new_n223), .B2(new_n256), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT66), .B(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n252), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n227), .A2(new_n225), .A3(KEYINPUT10), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n248), .A2(new_n237), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G140), .ZN(new_n266));
  INV_X1    g080(.A(G227), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G953), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n266), .B(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n228), .A2(KEYINPUT12), .A3(new_n238), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n244), .B1(new_n243), .B2(new_n237), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT79), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n246), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n263), .A2(new_n264), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT10), .B1(new_n241), .B2(new_n242), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT78), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT78), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n248), .A2(new_n279), .A3(new_n263), .A4(new_n264), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n280), .A3(new_n238), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n270), .B1(new_n281), .B2(new_n265), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n275), .B1(new_n282), .B2(KEYINPUT80), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n284));
  AOI211_X1 g098(.A(new_n284), .B(new_n270), .C1(new_n281), .C2(new_n265), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n187), .B(new_n188), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n272), .A2(new_n273), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT77), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n265), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n288), .B1(new_n287), .B2(new_n265), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n269), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n271), .A2(new_n281), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(G469), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(G469), .A2(G902), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n286), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  OAI21_X1  g111(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G237), .A2(G953), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G214), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n190), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(G143), .A3(G214), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(KEYINPUT18), .A3(G131), .ZN(new_n305));
  INV_X1    g119(.A(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G125), .ZN(new_n307));
  INV_X1    g121(.A(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G146), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n309), .A3(new_n193), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(KEYINPUT18), .A2(G131), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n302), .A2(new_n303), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n305), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n300), .A2(G143), .A3(G214), .ZN(new_n317));
  AOI21_X1  g131(.A(G143), .B1(new_n300), .B2(G214), .ZN(new_n318));
  OAI21_X1  g132(.A(G131), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n302), .A2(new_n236), .A3(new_n303), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT17), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n306), .A3(G125), .ZN(new_n326));
  OAI211_X1 g140(.A(G146), .B(new_n326), .C1(new_n310), .C2(new_n325), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n310), .B2(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n193), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n304), .A2(KEYINPUT17), .A3(G131), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n316), .B1(new_n324), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G113), .B(G122), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(new_n207), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n336), .B(new_n316), .C1(new_n324), .C2(new_n333), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n188), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G475), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT19), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT19), .B1(new_n307), .B2(new_n309), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n193), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT86), .A3(new_n327), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n319), .A2(new_n320), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT86), .B1(new_n345), .B2(new_n327), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n316), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n336), .B1(new_n350), .B2(KEYINPUT87), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n352), .B(new_n316), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  INV_X1    g167(.A(new_n316), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n322), .B(KEYINPUT88), .ZN(new_n355));
  INV_X1    g169(.A(new_n333), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n351), .A2(new_n353), .B1(new_n357), .B2(new_n336), .ZN(new_n358));
  NOR2_X1   g172(.A1(G475), .A2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n358), .A2(KEYINPUT20), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n351), .A2(new_n353), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n339), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n362), .B1(new_n364), .B2(new_n359), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n342), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT89), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT20), .B1(new_n358), .B2(new_n360), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n362), .A3(new_n359), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n368), .A2(new_n369), .B1(G475), .B2(new_n341), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G217), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n297), .A2(new_n374), .A3(G953), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT95), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n378));
  INV_X1    g192(.A(G122), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(G116), .ZN(new_n380));
  INV_X1    g194(.A(G116), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT90), .A3(G122), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G116), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n205), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT91), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n201), .B2(G143), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n190), .A2(KEYINPUT91), .A3(G128), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(G128), .B2(new_n190), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(G134), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(G134), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n385), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n380), .A2(new_n394), .A3(new_n382), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n384), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT93), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT93), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n383), .A2(new_n399), .A3(KEYINPUT14), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT94), .B1(new_n401), .B2(new_n205), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n399), .B1(new_n383), .B2(KEYINPUT14), .ZN(new_n403));
  AOI211_X1 g217(.A(KEYINPUT93), .B(new_n394), .C1(new_n380), .C2(new_n382), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n384), .B(new_n395), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT94), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(G107), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n393), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n383), .A2(new_n384), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G107), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n385), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(G134), .B2(new_n390), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n387), .A2(new_n388), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT13), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n190), .A2(G128), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT92), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT92), .ZN(new_n417));
  OAI221_X1 g231(.A(new_n417), .B1(G128), .B2(new_n190), .C1(new_n413), .C2(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(KEYINPUT13), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n412), .B1(new_n420), .B2(G134), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n377), .B1(new_n408), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n393), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n401), .A2(KEYINPUT94), .A3(new_n205), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n406), .B1(new_n405), .B2(G107), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(G134), .ZN(new_n427));
  INV_X1    g241(.A(new_n412), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n429), .A3(new_n376), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n422), .A2(new_n430), .A3(new_n188), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT96), .B1(new_n431), .B2(KEYINPUT97), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT96), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n422), .A2(new_n430), .A3(new_n433), .A4(new_n188), .ZN(new_n434));
  INV_X1    g248(.A(G478), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n432), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n373), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G952), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G953), .ZN(new_n442));
  NAND2_X1  g256(.A1(G234), .A2(G237), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(G902), .A3(G953), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(G898), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n452));
  INV_X1    g266(.A(G119), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(G116), .ZN(new_n454));
  XOR2_X1   g268(.A(G116), .B(G119), .Z(new_n455));
  OAI211_X1 g269(.A(G113), .B(new_n454), .C1(new_n455), .C2(new_n452), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT2), .B(G113), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n226), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n455), .B(new_n457), .Z(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n252), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n462), .B2(KEYINPUT81), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n252), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G122), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n463), .A2(new_n467), .A3(new_n465), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(KEYINPUT6), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n225), .A2(G125), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(G125), .B2(new_n259), .ZN(new_n473));
  INV_X1    g287(.A(G224), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G953), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT82), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n473), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n466), .A2(new_n478), .A3(new_n468), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT85), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n475), .B2(KEYINPUT84), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n473), .B(new_n485), .C1(KEYINPUT84), .C2(new_n475), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n458), .B(new_n227), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n467), .B(KEYINPUT8), .Z(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n472), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n484), .B2(new_n475), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n473), .B2(KEYINPUT83), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n494), .B2(new_n470), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n480), .A2(new_n483), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n483), .B1(new_n480), .B2(new_n495), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n450), .B(new_n451), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n299), .A2(new_n440), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n201), .A2(G119), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n453), .A2(G128), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT72), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT24), .B(G110), .Z(new_n506));
  NAND3_X1  g320(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n507));
  INV_X1    g321(.A(new_n502), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n503), .B(new_n507), .C1(new_n508), .C2(KEYINPUT23), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n505), .A2(new_n506), .B1(G110), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n505), .A2(new_n506), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n509), .A2(G110), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n327), .B(new_n312), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT22), .B(G137), .ZN(new_n516));
  INV_X1    g330(.A(G953), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n517), .A2(G221), .A3(G234), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n516), .B(new_n518), .Z(new_n519));
  XNOR2_X1  g333(.A(new_n515), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n188), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n374), .B1(G234), .B2(new_n188), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n520), .B(KEYINPUT74), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(G902), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G472), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n300), .A2(G210), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT27), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT26), .B(G101), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n261), .A2(new_n238), .A3(new_n262), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n235), .A2(G131), .ZN(new_n538));
  INV_X1    g352(.A(new_n232), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n230), .A2(G137), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n225), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n460), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(KEYINPUT71), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n537), .A2(new_n542), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n461), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n537), .A2(new_n550), .A3(new_n460), .A4(new_n542), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI211_X1 g366(.A(new_n536), .B(new_n546), .C1(new_n552), .C2(KEYINPUT28), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n537), .A2(KEYINPUT30), .A3(new_n542), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n542), .B1(new_n237), .B2(new_n259), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n460), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n543), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT29), .B1(new_n559), .B2(new_n536), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n537), .A2(KEYINPUT28), .A3(new_n460), .A4(new_n542), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n461), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n545), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n535), .B(KEYINPUT68), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n564), .A2(KEYINPUT29), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n553), .A2(new_n560), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n531), .B1(new_n566), .B2(new_n188), .ZN(new_n567));
  NOR2_X1   g381(.A1(G472), .A2(G902), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n543), .A2(new_n535), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n554), .B2(new_n557), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n571), .A2(new_n572), .B1(new_n563), .B2(new_n564), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n554), .A2(new_n557), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT31), .B1(new_n574), .B2(new_n570), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT67), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n558), .A2(new_n543), .A3(new_n535), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT67), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT31), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT69), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT69), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n573), .A2(new_n582), .A3(new_n576), .A4(new_n579), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n569), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n567), .B1(new_n584), .B2(KEYINPUT32), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT31), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n578), .B1(new_n577), .B2(KEYINPUT31), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n582), .B1(new_n588), .B2(new_n573), .ZN(new_n589));
  AND4_X1   g403(.A1(new_n582), .A2(new_n573), .A3(new_n576), .A4(new_n579), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n568), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n530), .B1(new_n585), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n500), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n598));
  AOI21_X1  g412(.A(G902), .B1(new_n581), .B2(new_n583), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n529), .B(new_n591), .C1(new_n531), .C2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n600), .B2(new_n299), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n188), .B1(new_n589), .B2(new_n590), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n584), .B1(new_n602), .B2(G472), .ZN(new_n603));
  INV_X1    g417(.A(new_n298), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n287), .A2(new_n265), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT77), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n289), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n607), .A2(new_n269), .B1(new_n281), .B2(new_n271), .ZN(new_n608));
  OAI21_X1  g422(.A(G469), .B1(new_n608), .B2(G902), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n604), .B1(new_n609), .B2(new_n286), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n603), .A2(new_n610), .A3(KEYINPUT98), .A4(new_n529), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n431), .A2(new_n435), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n422), .A2(new_n430), .A3(KEYINPUT33), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT33), .B1(new_n422), .B2(new_n430), .ZN(new_n617));
  OAI211_X1 g431(.A(G478), .B(new_n188), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n367), .A3(new_n372), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n499), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n612), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  NOR3_X1   g438(.A1(new_n499), .A2(new_n366), .A3(new_n439), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n612), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  OAI21_X1  g442(.A(new_n591), .B1(new_n599), .B2(new_n531), .ZN(new_n629));
  INV_X1    g443(.A(new_n525), .ZN(new_n630));
  INV_X1    g444(.A(new_n519), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n515), .B(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(new_n527), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n500), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  OAI21_X1  g453(.A(new_n451), .B1(new_n497), .B2(new_n498), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n630), .A2(new_n634), .ZN(new_n642));
  OAI211_X1 g456(.A(KEYINPUT32), .B(new_n568), .C1(new_n589), .C2(new_n590), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n566), .A2(new_n188), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G472), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n584), .A2(new_n592), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n641), .B(new_n642), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n447), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n444), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n370), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n439), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n610), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT100), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n635), .B1(new_n585), .B2(new_n594), .ZN(new_n656));
  INV_X1    g470(.A(new_n653), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n299), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n656), .A2(new_n658), .A3(new_n659), .A4(new_n641), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  INV_X1    g476(.A(new_n451), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n438), .A2(new_n367), .A3(new_n372), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n642), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n651), .B(KEYINPUT39), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n610), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n571), .B1(new_n564), .B2(new_n552), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n594), .A2(new_n643), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n497), .A2(new_n498), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n666), .A2(new_n669), .A3(new_n670), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  INV_X1    g493(.A(new_n651), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n620), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n656), .A2(new_n610), .A3(new_n641), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  OAI211_X1 g497(.A(new_n643), .B(new_n645), .C1(new_n584), .C2(new_n592), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n188), .B1(new_n283), .B2(new_n285), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n686), .A2(new_n298), .A3(new_n286), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n684), .A2(new_n687), .A3(new_n529), .A4(new_n621), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n595), .A2(KEYINPUT102), .A3(new_n621), .A4(new_n687), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT103), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n692), .B(new_n694), .ZN(G15));
  NAND4_X1  g509(.A1(new_n684), .A2(new_n625), .A3(new_n687), .A4(new_n529), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  NAND3_X1  g511(.A1(new_n686), .A2(new_n298), .A3(new_n286), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n640), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n373), .A2(new_n439), .A3(new_n450), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n699), .A2(new_n684), .A3(new_n642), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G119), .ZN(G21));
  AND2_X1   g517(.A1(new_n552), .A2(KEYINPUT28), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n564), .B1(new_n704), .B2(new_n546), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n577), .B(new_n572), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n569), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n599), .B2(new_n531), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n602), .A2(KEYINPUT104), .A3(G472), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n707), .B(new_n530), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n438), .A2(new_n367), .A3(new_n713), .A4(new_n372), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n499), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n715), .A2(new_n687), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n711), .A2(new_n717), .A3(KEYINPUT106), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  INV_X1    g533(.A(new_n707), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT104), .B1(new_n602), .B2(G472), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n599), .A2(new_n708), .A3(new_n531), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n529), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n715), .A2(new_n687), .A3(new_n716), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  AOI21_X1  g541(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n642), .A3(new_n681), .A4(new_n699), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT107), .B(G125), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G27));
  NAND2_X1  g545(.A1(new_n480), .A2(new_n495), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n482), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n604), .A2(new_n663), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n496), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n609), .B2(new_n286), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT108), .ZN(new_n737));
  INV_X1    g551(.A(new_n735), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n296), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  OR3_X1    g557(.A1(new_n584), .A2(new_n743), .A3(KEYINPUT32), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n743), .B1(new_n584), .B2(KEYINPUT32), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n585), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n742), .A2(new_n746), .A3(new_n529), .A4(new_n681), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n296), .A2(new_n738), .A3(KEYINPUT108), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT108), .B1(new_n296), .B2(new_n738), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n684), .A2(new_n529), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n620), .A2(KEYINPUT42), .A3(new_n680), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n747), .A2(KEYINPUT42), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  NAND3_X1  g569(.A1(new_n742), .A2(new_n595), .A3(new_n653), .ZN(new_n756));
  XOR2_X1   g570(.A(KEYINPUT110), .B(G134), .Z(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G36));
  NAND2_X1  g572(.A1(new_n675), .A2(new_n451), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n373), .A2(new_n619), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT43), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n761), .A2(new_n603), .A3(new_n635), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n292), .A2(new_n293), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n187), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n608), .A2(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT46), .B1(new_n770), .B2(new_n295), .ZN(new_n771));
  INV_X1    g585(.A(new_n286), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(KEYINPUT46), .A3(new_n295), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n604), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n667), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n765), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n233), .ZN(G39));
  NOR2_X1   g593(.A1(new_n759), .A2(new_n529), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n681), .A3(new_n594), .A4(new_n585), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n776), .A2(KEYINPUT47), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n306), .ZN(G42));
  NOR2_X1   g600(.A1(new_n761), .A2(new_n444), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n711), .ZN(new_n788));
  INV_X1    g602(.A(new_n784), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n782), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n686), .A2(new_n286), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n604), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n759), .B(new_n788), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n698), .A2(new_n759), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n674), .A2(new_n529), .A3(new_n445), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT117), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n373), .A3(new_n615), .A4(new_n618), .ZN(new_n798));
  INV_X1    g612(.A(new_n788), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n451), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n676), .A2(new_n687), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n799), .B(new_n803), .C1(new_n800), .C2(new_n801), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n787), .A2(new_n795), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n642), .A3(new_n728), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n798), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n793), .A2(new_n794), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n794), .B1(new_n793), .B2(new_n809), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(new_n529), .A3(new_n746), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT48), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n799), .A2(new_n699), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n442), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n620), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n797), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n655), .A2(new_n660), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n640), .B1(new_n712), .B2(new_n714), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n642), .A2(new_n680), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n673), .A4(new_n610), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n729), .A2(new_n682), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT52), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n682), .A2(new_n822), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n661), .A4(new_n729), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n702), .A2(new_n696), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n690), .B2(new_n691), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n754), .A2(new_n830), .A3(new_n726), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n438), .A2(new_n652), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n684), .A2(new_n642), .A3(new_n736), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n656), .A2(KEYINPUT113), .A3(new_n736), .A4(new_n833), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n742), .A2(new_n642), .A3(new_n681), .A4(new_n728), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n756), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n440), .B1(new_n373), .B2(new_n619), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n499), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n601), .A2(new_n611), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n500), .B1(new_n595), .B2(new_n636), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n832), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n829), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT106), .B1(new_n711), .B2(new_n717), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n723), .A2(new_n724), .A3(new_n719), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n850), .B(new_n692), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n752), .A2(new_n753), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n846), .A3(new_n824), .A4(new_n827), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n849), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT115), .B1(new_n840), .B2(new_n845), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n839), .A2(new_n756), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n843), .A2(new_n844), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n838), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n832), .A2(new_n868), .A3(KEYINPUT53), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n858), .A2(new_n847), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n818), .A2(new_n873), .B1(G952), .B2(G953), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT49), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n791), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT112), .Z(new_n877));
  NAND2_X1  g691(.A1(new_n529), .A2(new_n734), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT111), .ZN(new_n879));
  INV_X1    g693(.A(new_n760), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n674), .A2(new_n879), .A3(new_n676), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n875), .B2(new_n791), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n874), .B1(new_n877), .B2(new_n882), .ZN(G75));
  NOR2_X1   g697(.A1(new_n517), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n188), .B1(new_n869), .B2(new_n870), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT56), .B1(new_n886), .B2(new_n482), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n471), .A2(new_n479), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(new_n477), .Z(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT55), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n885), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n887), .B2(new_n891), .ZN(G51));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n188), .B(new_n770), .C1(new_n869), .C2(new_n870), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n295), .B(KEYINPUT57), .Z(new_n896));
  AND3_X1   g710(.A1(new_n869), .A2(new_n871), .A3(new_n870), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n871), .B1(new_n869), .B2(new_n870), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n283), .A2(new_n285), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n895), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n894), .B1(new_n902), .B2(new_n884), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n864), .A2(new_n866), .A3(new_n838), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n828), .A2(new_n904), .A3(new_n831), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n857), .A2(KEYINPUT53), .A3(new_n824), .A4(new_n827), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n863), .A2(new_n867), .ZN(new_n907));
  OAI22_X1  g721(.A1(new_n905), .A2(new_n848), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n872), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n900), .B1(new_n910), .B2(new_n896), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT118), .B(new_n885), .C1(new_n911), .C2(new_n895), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n903), .A2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(new_n358), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n358), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n884), .ZN(G60));
  OR2_X1    g731(.A1(new_n616), .A2(new_n617), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT59), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n910), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n885), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n918), .B1(new_n873), .B2(new_n921), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT119), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n884), .B1(new_n910), .B2(new_n922), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n920), .B1(new_n862), .B2(new_n872), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n927), .B(new_n928), .C1(new_n918), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n926), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n908), .A2(new_n633), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n869), .B2(new_n870), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n633), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n885), .A2(KEYINPUT61), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n526), .B1(new_n908), .B2(new_n934), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(KEYINPUT122), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n940), .B(new_n943), .C1(KEYINPUT122), .C2(new_n942), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT121), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(new_n885), .C1(new_n937), .C2(new_n526), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT121), .B1(new_n942), .B2(new_n884), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n940), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n944), .B1(new_n948), .B2(KEYINPUT61), .ZN(G66));
  NAND3_X1  g763(.A1(new_n830), .A2(new_n726), .A3(new_n866), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n517), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT123), .Z(new_n952));
  OAI21_X1  g766(.A(G953), .B1(new_n448), .B2(new_n474), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT124), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n888), .B1(G898), .B2(new_n517), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  OAI21_X1  g771(.A(G953), .B1(new_n267), .B2(new_n649), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT126), .Z(new_n959));
  NOR4_X1   g773(.A1(new_n751), .A2(new_n668), .A3(new_n759), .A4(new_n841), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n785), .A2(new_n778), .A3(new_n960), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n661), .A2(new_n682), .A3(new_n729), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n678), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n517), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n555), .A2(new_n556), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n554), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n343), .A2(new_n344), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(G900), .B2(G953), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n746), .A2(new_n529), .A3(new_n820), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n777), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n756), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n977), .A2(new_n856), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n790), .B2(new_n781), .ZN(new_n980));
  INV_X1    g794(.A(new_n778), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n962), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT125), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n984), .A3(new_n962), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n980), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n975), .B1(new_n986), .B2(new_n517), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n959), .B1(new_n973), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n959), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n986), .A2(new_n517), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n989), .B(new_n972), .C1(new_n990), .C2(new_n975), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n966), .B2(new_n950), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n559), .B(KEYINPUT127), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n535), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n885), .ZN(new_n998));
  INV_X1    g812(.A(new_n994), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n571), .B1(new_n536), .B2(new_n559), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n999), .B(new_n1000), .C1(new_n849), .C2(new_n860), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n996), .A2(new_n535), .ZN(new_n1002));
  INV_X1    g816(.A(new_n950), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n986), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1002), .B1(new_n1004), .B2(new_n994), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n998), .A2(new_n1001), .A3(new_n1005), .ZN(G57));
endmodule


