//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n210), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(G50), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n208), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n213), .A2(new_n224), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  INV_X1    g0046(.A(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n215), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n246), .B(new_n252), .ZN(G351));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT71), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n208), .A2(G33), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT15), .B(G87), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n257), .B1(new_n208), .B2(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n227), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(new_n227), .A3(new_n262), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n258), .B1(new_n207), .B2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n265), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n267), .A2(new_n268), .B1(new_n258), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1698), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G232), .ZN(new_n277));
  INV_X1    g0077(.A(G107), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n274), .A2(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G1698), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n277), .B1(new_n278), .B2(new_n279), .C1(new_n216), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(G1), .A2(G13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(KEYINPUT69), .A3(new_n282), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n286), .B2(new_n282), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT68), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n207), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n291), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n283), .A2(new_n292), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(G244), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n271), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(G190), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(G200), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n264), .A3(new_n270), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g0109(.A(new_n309), .B(KEYINPUT72), .Z(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n262), .A2(new_n311), .A3(new_n227), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n262), .B2(new_n227), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n269), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(G50), .C1(G1), .C2(new_n208), .ZN(new_n316));
  INV_X1    g0116(.A(G150), .ZN(new_n317));
  INV_X1    g0117(.A(new_n256), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n254), .A2(new_n259), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n208), .B1(new_n201), .B2(new_n247), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n314), .B1(new_n247), .B2(new_n269), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n297), .A2(G226), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n276), .A2(G222), .ZN(new_n325));
  INV_X1    g0125(.A(G223), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n325), .B1(new_n258), .B2(new_n279), .C1(new_n326), .C2(new_n280), .ZN(new_n327));
  AOI211_X1 g0127(.A(new_n296), .B(new_n324), .C1(new_n327), .C2(new_n288), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n323), .B1(new_n328), .B2(G169), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n301), .B2(new_n328), .ZN(new_n330));
  XOR2_X1   g0130(.A(new_n323), .B(KEYINPUT9), .Z(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT73), .B1(new_n328), .B2(G190), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n328), .ZN(new_n334));
  OR3_X1    g0134(.A1(new_n331), .A2(new_n334), .A3(KEYINPUT10), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT10), .B1(new_n331), .B2(new_n334), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n330), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n256), .A2(G50), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n338), .B(new_n339), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n259), .A2(new_n258), .B1(new_n208), .B2(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n314), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT11), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT12), .B1(new_n265), .B2(G68), .ZN(new_n346));
  OR3_X1    g0146(.A1(new_n265), .A2(KEYINPUT12), .A3(G68), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n215), .B1(new_n207), .B2(G20), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n346), .A2(new_n347), .B1(new_n267), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n344), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n291), .A2(new_n294), .A3(KEYINPUT74), .A4(new_n295), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n283), .A2(G238), .A3(new_n292), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G226), .A2(G1698), .ZN(new_n354));
  INV_X1    g0154(.A(G232), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(G1698), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n279), .B1(G33), .B2(G97), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n285), .A2(new_n287), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n352), .B(new_n353), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n291), .A2(new_n294), .A3(new_n295), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT74), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT76), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n353), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G97), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n355), .A2(G1698), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(G226), .B2(G1698), .ZN(new_n368));
  AND2_X1   g0168(.A1(KEYINPUT3), .A2(G33), .ZN(new_n369));
  NOR2_X1   g0169(.A1(KEYINPUT3), .A2(G33), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n366), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n365), .B1(new_n288), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(new_n362), .A4(new_n352), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n364), .A2(new_n375), .A3(KEYINPUT13), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n377));
  NAND4_X1  g0177(.A1(new_n373), .A2(new_n377), .A3(new_n362), .A4(new_n352), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G179), .ZN(new_n379));
  INV_X1    g0179(.A(new_n377), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n359), .B2(new_n363), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n303), .B1(new_n381), .B2(new_n378), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT14), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n376), .A2(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT79), .B1(new_n382), .B2(new_n383), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n382), .A2(KEYINPUT79), .A3(new_n383), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n351), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n381), .A2(new_n378), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G200), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n351), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n364), .A2(new_n375), .A3(KEYINPUT13), .ZN(new_n392));
  INV_X1    g0192(.A(G190), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n359), .A2(new_n363), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n377), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT77), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n395), .A3(KEYINPUT77), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n388), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n279), .B2(G20), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n371), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n215), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  OAI21_X1  g0207(.A(G20), .B1(new_n407), .B2(new_n201), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n256), .A2(G159), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n402), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT7), .B1(new_n371), .B2(new_n208), .ZN(new_n412));
  NOR4_X1   g0212(.A1(new_n369), .A2(new_n370), .A3(new_n403), .A4(G20), .ZN(new_n413));
  OAI21_X1  g0213(.A(G68), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n410), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(new_n263), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n254), .B1(new_n207), .B2(G20), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n315), .A2(new_n418), .B1(new_n269), .B2(new_n254), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G1698), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n326), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G226), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n422), .B(new_n424), .C1(new_n369), .C2(new_n370), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT80), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(KEYINPUT80), .A3(new_n426), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n358), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n283), .A2(G232), .A3(new_n292), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT81), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT81), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n283), .A2(new_n292), .A3(new_n434), .A4(G232), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n360), .ZN(new_n437));
  OAI21_X1  g0237(.A(G169), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n425), .A2(KEYINPUT80), .A3(new_n426), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT80), .B1(new_n425), .B2(new_n426), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n288), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n296), .B1(new_n433), .B2(new_n435), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(G179), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n420), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT18), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n431), .A2(new_n437), .A3(G190), .ZN(new_n447));
  AOI21_X1  g0247(.A(G200), .B1(new_n441), .B2(new_n442), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n419), .B(new_n417), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n315), .A2(new_n418), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n254), .A2(new_n269), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n263), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n414), .A2(new_n415), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n402), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n416), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n333), .B1(new_n431), .B2(new_n437), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n441), .A2(new_n442), .A3(new_n393), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n461), .A3(KEYINPUT17), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT18), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n420), .A2(new_n444), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n446), .A2(new_n451), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n310), .A2(new_n337), .A3(new_n401), .A4(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n207), .A2(G33), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G116), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n267), .A2(KEYINPUT85), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT85), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n266), .B2(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n265), .A2(G116), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT86), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(G20), .B1(new_n273), .B2(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT82), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT82), .B1(G33), .B2(G283), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G116), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n262), .A2(new_n227), .B1(G20), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n485), .A2(KEYINPUT87), .A3(KEYINPUT20), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT20), .B1(new_n485), .B2(new_n487), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n485), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n479), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(G264), .B(G1698), .C1(new_n369), .C2(new_n370), .ZN(new_n496));
  OAI211_X1 g0296(.A(G257), .B(new_n421), .C1(new_n369), .C2(new_n370), .ZN(new_n497));
  INV_X1    g0297(.A(G303), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n496), .B(new_n497), .C1(new_n498), .C2(new_n279), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n288), .ZN(new_n500));
  INV_X1    g0300(.A(G41), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n207), .B(G45), .C1(new_n501), .C2(KEYINPUT5), .ZN(new_n504));
  OAI211_X1 g0304(.A(G270), .B(new_n283), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G45), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G1), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT83), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n507), .B(new_n508), .C1(KEYINPUT5), .C2(new_n501), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n504), .A2(KEYINPUT83), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n509), .A2(new_n510), .A3(new_n291), .A4(new_n502), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n500), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G169), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n468), .B1(new_n495), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n276), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n279), .A2(G257), .A3(G1698), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n358), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G264), .B(new_n283), .C1(new_n503), .C2(new_n504), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n303), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n517), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n301), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n259), .A2(new_n486), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT90), .B1(new_n208), .B2(G107), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT23), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI211_X1 g0327(.A(KEYINPUT90), .B(new_n527), .C1(new_n208), .C2(G107), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n208), .B(G87), .C1(new_n369), .C2(new_n370), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n530), .A2(KEYINPUT22), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(KEYINPUT22), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT24), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n529), .C1(new_n531), .C2(new_n532), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n455), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  XOR2_X1   g0337(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n538));
  NOR2_X1   g0338(.A1(new_n265), .A2(G107), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n312), .A2(new_n313), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n265), .A3(new_n469), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n544), .B2(new_n278), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n521), .B(new_n523), .C1(new_n537), .C2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n499), .A2(new_n288), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n511), .A2(new_n505), .ZN(new_n548));
  OAI211_X1 g0348(.A(KEYINPUT21), .B(G169), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n500), .A2(G179), .A3(new_n505), .A4(new_n511), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n485), .A2(new_n487), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n494), .B(new_n488), .C1(KEYINPUT20), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n475), .A3(new_n478), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n551), .A2(KEYINPUT88), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT88), .B1(new_n551), .B2(new_n554), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n514), .B(new_n546), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G238), .B(new_n421), .C1(new_n369), .C2(new_n370), .ZN(new_n558));
  OAI211_X1 g0358(.A(G244), .B(G1698), .C1(new_n369), .C2(new_n370), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n273), .C2(new_n486), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n288), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n507), .A2(new_n290), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n218), .B1(new_n506), .B2(G1), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n283), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n208), .B1(new_n366), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G87), .B2(new_n205), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n208), .B(G68), .C1(new_n369), .C2(new_n370), .ZN(new_n570));
  INV_X1    g0370(.A(G97), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n259), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n263), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n260), .A2(new_n269), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n543), .A2(G87), .A3(new_n265), .A4(new_n469), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n564), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n560), .B2(new_n288), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G190), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n566), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n565), .A2(new_n303), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n574), .B(new_n575), .C1(new_n260), .C2(new_n544), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n301), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n520), .A2(G200), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n522), .A2(G190), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n537), .A2(new_n545), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT6), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n592), .A2(new_n571), .A3(G107), .ZN(new_n593));
  XNOR2_X1  g0393(.A(G97), .B(G107), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n595), .A2(new_n208), .B1(new_n258), .B2(new_n318), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n278), .B1(new_n404), .B2(new_n405), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n263), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OR2_X1    g0398(.A1(new_n544), .A2(new_n571), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n265), .A2(G97), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT84), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n598), .A2(new_n599), .A3(new_n604), .A4(new_n601), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G257), .B(new_n283), .C1(new_n503), .C2(new_n504), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(G244), .B(new_n421), .C1(new_n369), .C2(new_n370), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT4), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n421), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n483), .A2(new_n484), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n611), .A2(new_n612), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n608), .B1(new_n615), .B2(new_n288), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n511), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G169), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(G179), .A3(new_n511), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n606), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n512), .A2(G200), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n495), .B(new_n622), .C1(new_n393), .C2(new_n512), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n617), .A2(G200), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n616), .A2(G190), .A3(new_n511), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n591), .A2(new_n621), .A3(new_n623), .A4(new_n627), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n467), .A2(new_n557), .A3(new_n628), .ZN(G372));
  NAND2_X1  g0429(.A1(new_n335), .A2(new_n336), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT92), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n398), .A2(new_n399), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n350), .B1(G200), .B2(new_n389), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n305), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n388), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n451), .A2(new_n462), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n399), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT77), .B1(new_n392), .B2(new_n395), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n634), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n305), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n389), .A2(new_n383), .A3(G169), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT79), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n389), .A2(G169), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT14), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n392), .A2(G179), .A3(new_n378), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n646), .A2(new_n648), .A3(new_n649), .A4(new_n387), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n350), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n643), .A2(new_n651), .A3(KEYINPUT92), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n636), .A2(new_n638), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n446), .A2(new_n464), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n631), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT93), .B1(new_n655), .B2(new_n330), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT93), .ZN(new_n657));
  INV_X1    g0457(.A(new_n330), .ZN(new_n658));
  INV_X1    g0458(.A(new_n654), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n643), .A2(new_n651), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n637), .B1(new_n660), .B2(new_n632), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n661), .B2(new_n652), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n657), .B(new_n658), .C1(new_n662), .C2(new_n631), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n467), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n551), .A2(new_n554), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n546), .A2(new_n514), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n591), .A2(new_n667), .A3(new_n621), .A4(new_n627), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n621), .B2(new_n586), .ZN(new_n669));
  INV_X1    g0469(.A(new_n585), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n616), .A2(G179), .A3(new_n511), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n303), .B1(new_n616), .B2(new_n511), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n602), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n586), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n668), .A2(new_n669), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n665), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n664), .A2(new_n678), .ZN(G369));
  NAND2_X1  g0479(.A1(new_n534), .A2(new_n536), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n263), .ZN(new_n681));
  INV_X1    g0481(.A(new_n545), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n681), .A2(new_n587), .A3(new_n682), .A4(new_n588), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n683), .B1(new_n590), .B2(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n546), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n546), .A2(new_n689), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n514), .B1(new_n555), .B2(new_n556), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(new_n690), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n693), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n694), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n495), .A2(new_n690), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n514), .A2(new_n666), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n623), .ZN(new_n703));
  INV_X1    g0503(.A(new_n701), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(new_n695), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n699), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n211), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G1), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n204), .A2(new_n217), .A3(new_n486), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT94), .Z(new_n714));
  OAI22_X1  g0514(.A1(new_n712), .A2(new_n714), .B1(new_n225), .B2(new_n711), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n581), .A2(new_n585), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(new_n606), .A3(new_n675), .A4(new_n620), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT26), .B1(new_n673), .B2(new_n586), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n718), .A2(new_n585), .A3(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n603), .A2(new_n605), .B1(new_n618), .B2(new_n619), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n557), .A2(new_n723), .A3(new_n591), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n689), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT29), .B1(new_n677), .B2(new_n690), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n628), .A2(new_n557), .A3(new_n689), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n522), .A2(new_n579), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n301), .A3(new_n512), .A4(new_n617), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n515), .A2(new_n516), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n288), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(new_n579), .A3(new_n511), .A4(new_n518), .ZN(new_n734));
  INV_X1    g0534(.A(new_n616), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n734), .A2(new_n735), .A3(new_n550), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n731), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NOR4_X1   g0538(.A1(new_n734), .A2(new_n735), .A3(new_n550), .A4(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n689), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n741), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n689), .B(new_n743), .C1(new_n737), .C2(new_n739), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(G330), .B1(new_n729), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n728), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n716), .B1(new_n748), .B2(G1), .ZN(G364));
  NAND2_X1  g0549(.A1(new_n208), .A2(G13), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT97), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G45), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G1), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n710), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n709), .A2(new_n371), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n756), .A2(G355), .B1(new_n486), .B2(new_n709), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n709), .A2(new_n279), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n226), .B2(G45), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n252), .A2(new_n506), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT98), .ZN(new_n762));
  OR3_X1    g0562(.A1(new_n762), .A2(G13), .A3(G33), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(G13), .B2(G33), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n227), .B1(G20), .B2(new_n303), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n755), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n768), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n393), .A2(new_n333), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n208), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n333), .A2(G190), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n774), .A2(new_n498), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n208), .A2(new_n301), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n780), .A2(new_n393), .A3(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n279), .B1(new_n781), .B2(G322), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n779), .A2(new_n775), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT33), .B(G317), .Z(new_n787));
  OAI221_X1 g0587(.A(new_n782), .B1(new_n783), .B2(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n773), .A2(new_n784), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n778), .B(new_n788), .C1(G329), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n779), .A2(new_n772), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  INV_X1    g0593(.A(G326), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n393), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n208), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT101), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n797), .A2(new_n571), .ZN(new_n800));
  INV_X1    g0600(.A(new_n786), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(G68), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT99), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n371), .B1(new_n781), .B2(G58), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  OR3_X1    g0605(.A1(new_n789), .A2(KEYINPUT32), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT32), .B1(new_n789), .B2(new_n805), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n774), .A2(new_n217), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n776), .A2(new_n278), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n792), .A2(new_n247), .B1(new_n785), .B2(new_n258), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n791), .A2(new_n799), .B1(new_n803), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n767), .B(KEYINPUT102), .Z(new_n814));
  OAI221_X1 g0614(.A(new_n770), .B1(new_n771), .B2(new_n813), .C1(new_n705), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n705), .A2(G330), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT96), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n706), .A2(new_n755), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n765), .A2(new_n768), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n258), .ZN(new_n821));
  INV_X1    g0621(.A(new_n785), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n781), .A2(G143), .B1(G159), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n792), .C1(new_n317), .C2(new_n786), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n279), .B1(new_n774), .B2(new_n247), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n776), .A2(new_n215), .B1(new_n789), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n797), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n829), .B(new_n831), .C1(G58), .C2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n827), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n776), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n279), .B(new_n800), .C1(G87), .C2(new_n835), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n486), .A2(new_n785), .B1(new_n786), .B2(new_n777), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT103), .ZN(new_n838));
  INV_X1    g0638(.A(new_n792), .ZN(new_n839));
  INV_X1    g0639(.A(new_n774), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G303), .A2(new_n839), .B1(new_n840), .B2(G107), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n781), .A2(G294), .B1(G311), .B2(new_n790), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n836), .A2(new_n838), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n834), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n754), .B(new_n821), .C1(new_n844), .C2(new_n771), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n271), .A2(new_n689), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n308), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n305), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n642), .A2(new_n690), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n845), .B1(new_n850), .B2(new_n765), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n677), .A2(new_n690), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n850), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n305), .A2(new_n689), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n305), .B2(new_n847), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n677), .A2(new_n690), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n857), .A2(new_n746), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n754), .B1(new_n857), .B2(new_n746), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n851), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  INV_X1    g0661(.A(new_n595), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n486), .B(new_n229), .C1(new_n862), .C2(KEYINPUT35), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(KEYINPUT35), .B2(new_n862), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT36), .Z(new_n865));
  OR3_X1    g0665(.A1(new_n225), .A2(new_n258), .A3(new_n407), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n207), .B(G13), .C1(new_n866), .C2(new_n248), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OR3_X1    g0668(.A1(new_n467), .A2(new_n726), .A3(new_n727), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n664), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n856), .A2(new_n849), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n350), .A2(new_n689), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n651), .A2(new_n641), .A3(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n350), .B(new_n689), .C1(new_n400), .C2(new_n650), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT105), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n411), .A2(new_n314), .A3(new_n416), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n419), .ZN(new_n881));
  INV_X1    g0681(.A(new_n687), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n458), .A2(new_n461), .B1(new_n881), .B2(new_n444), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(KEYINPUT104), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n444), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n886), .A2(KEYINPUT104), .A3(new_n449), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n879), .B(KEYINPUT37), .C1(new_n885), .C2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n883), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n465), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n420), .A2(new_n882), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n445), .A2(new_n892), .A3(new_n449), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT105), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n884), .A2(KEYINPUT104), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n886), .A2(new_n449), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT104), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n899), .A3(new_n883), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n895), .B1(new_n900), .B2(KEYINPUT37), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n878), .B1(new_n891), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n895), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT104), .B1(new_n886), .B2(new_n449), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n887), .A2(new_n904), .A3(new_n889), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n905), .B2(new_n893), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n906), .A2(KEYINPUT38), .A3(new_n888), .A4(new_n890), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n877), .A2(new_n908), .B1(new_n659), .B2(new_n687), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n445), .A2(new_n892), .A3(new_n449), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n894), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n466), .B2(new_n892), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n878), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n651), .A2(new_n689), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n907), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n870), .B(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n850), .B1(new_n873), .B2(new_n874), .ZN(new_n924));
  AND4_X1   g0724(.A1(new_n621), .A2(new_n627), .A3(new_n683), .A4(new_n717), .ZN(new_n925));
  INV_X1    g0725(.A(new_n557), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n925), .A2(new_n926), .A3(new_n623), .A4(new_n690), .ZN(new_n927));
  NOR2_X1   g0727(.A1(KEYINPUT106), .A2(KEYINPUT31), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n740), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n689), .B(new_n928), .C1(new_n737), .C2(new_n739), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n907), .B2(new_n902), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT40), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n915), .A2(KEYINPUT40), .A3(new_n924), .A4(new_n933), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n665), .A2(new_n933), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(G330), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n923), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n207), .B2(new_n751), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n923), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n868), .B1(new_n944), .B2(new_n945), .ZN(G367));
  OR2_X1    g0746(.A1(new_n577), .A2(new_n690), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n717), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n585), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT43), .Z(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n723), .B1(new_n625), .B2(new_n690), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n620), .A2(new_n602), .A3(new_n689), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n694), .A3(new_n696), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT107), .ZN(new_n958));
  INV_X1    g0758(.A(new_n955), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n621), .B1(new_n959), .B2(new_n546), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n960), .A2(new_n690), .B1(KEYINPUT42), .B2(new_n956), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n952), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT109), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n958), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(KEYINPUT109), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT108), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n963), .A2(new_n969), .A3(new_n965), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n707), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n959), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n970), .A3(new_n973), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n710), .B(KEYINPUT41), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n699), .A2(new_n959), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n699), .A2(new_n959), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n972), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n694), .B(new_n696), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n705), .A2(KEYINPUT110), .A3(G330), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT110), .B1(new_n705), .B2(G330), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n985), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n747), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n979), .A2(new_n972), .A3(new_n982), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n984), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n977), .B1(new_n992), .B2(new_n748), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT111), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n753), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n993), .B2(new_n994), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n975), .B(new_n976), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n769), .B1(new_n211), .B2(new_n260), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n758), .A2(new_n241), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n754), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n835), .A2(G77), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n824), .B2(new_n789), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n371), .B(new_n1003), .C1(G58), .C2(new_n840), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n832), .A2(G68), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n793), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(G143), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n781), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1008), .A2(new_n317), .B1(new_n786), .B2(new_n805), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G50), .B2(new_n822), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n371), .B1(new_n785), .B2(new_n777), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n840), .A2(G116), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .C1(new_n278), .C2(new_n797), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n781), .A2(G303), .B1(G317), .B2(new_n790), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G294), .A2(new_n801), .B1(new_n835), .B2(G97), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n783), .C2(new_n793), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1011), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT47), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1001), .B1(new_n1021), .B2(new_n768), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n814), .B2(new_n950), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n998), .A2(new_n1023), .ZN(G387));
  INV_X1    g0824(.A(new_n990), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n989), .A2(new_n747), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1025), .A2(new_n710), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n756), .A2(new_n714), .B1(new_n278), .B2(new_n709), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n255), .A2(new_n247), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT50), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n506), .B1(new_n215), .B2(new_n258), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1030), .A2(new_n714), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n758), .B1(new_n237), .B2(new_n506), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1028), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n755), .B1(new_n1034), .B2(new_n769), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n371), .B1(new_n835), .B2(G97), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n215), .B2(new_n785), .C1(new_n258), .C2(new_n774), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1008), .A2(new_n247), .B1(new_n254), .B2(new_n786), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n792), .A2(new_n805), .B1(new_n789), .B2(new_n317), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n797), .A2(new_n260), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n781), .A2(G317), .B1(G311), .B2(new_n801), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n498), .B2(new_n785), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G322), .B2(new_n1006), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT48), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(KEYINPUT48), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n832), .A2(G283), .B1(new_n840), .B2(G294), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n371), .B1(new_n789), .B2(new_n794), .C1(new_n486), .C2(new_n776), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1049), .B2(KEYINPUT49), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1041), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1035), .B1(new_n694), .B2(new_n814), .C1(new_n1053), .C2(new_n771), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1027), .B(new_n1054), .C1(new_n996), .C2(new_n989), .ZN(G393));
  INV_X1    g0855(.A(new_n991), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1025), .B1(new_n1056), .B2(new_n983), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n992), .A3(new_n710), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n245), .A2(new_n709), .A3(new_n279), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n769), .B1(new_n571), .B2(new_n211), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n797), .A2(new_n258), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n371), .B(new_n1061), .C1(G87), .C2(new_n835), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n247), .A2(new_n786), .B1(new_n774), .B2(new_n215), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G143), .B2(new_n790), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n255), .B2(new_n822), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n781), .A2(G159), .B1(new_n839), .B2(G150), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  AOI22_X1  g0868(.A1(G303), .A2(new_n801), .B1(new_n790), .B2(G322), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n777), .B2(new_n774), .C1(new_n795), .C2(new_n785), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n797), .A2(new_n486), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1070), .A2(new_n279), .A3(new_n810), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n781), .A2(G311), .B1(new_n839), .B2(G317), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT52), .Z(new_n1074));
  AOI22_X1  g0874(.A1(new_n1066), .A2(new_n1068), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n754), .B1(new_n1059), .B2(new_n1060), .C1(new_n1075), .C2(new_n771), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n959), .B2(new_n767), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1056), .A2(new_n983), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n753), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1058), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT112), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1058), .A2(new_n1079), .A3(KEYINPUT112), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(KEYINPUT113), .ZN(new_n1085));
  INV_X1    g0885(.A(G330), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n927), .B2(new_n932), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1087), .A2(new_n924), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n856), .A2(new_n849), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n918), .B1(new_n1089), .B2(new_n875), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n917), .B2(new_n919), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n918), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n915), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n854), .B1(new_n725), .B2(new_n848), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n876), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1092), .B1(new_n871), .B2(new_n876), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n907), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n907), .B2(new_n914), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n915), .B(new_n1092), .C1(new_n876), .C2(new_n1094), .ZN(new_n1102));
  OAI211_X1 g0902(.A(G330), .B(new_n855), .C1(new_n729), .C2(new_n745), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(new_n876), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1103), .A2(new_n876), .B1(new_n1087), .B2(new_n924), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1094), .B1(new_n1103), .B2(new_n876), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n875), .B1(new_n1087), .B2(new_n855), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1107), .A2(new_n871), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n665), .A2(new_n1087), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n664), .A2(new_n1110), .A3(new_n869), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1085), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  AND4_X1   g0913(.A1(new_n664), .A2(new_n1110), .A3(new_n869), .A4(new_n1111), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1114), .A2(KEYINPUT113), .A3(new_n1105), .A4(new_n1097), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1106), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n710), .C1(new_n1117), .C2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n765), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n820), .A2(new_n254), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n774), .A2(new_n317), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT53), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n781), .A2(G132), .B1(G125), .B2(new_n790), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n1123), .C1(new_n785), .C2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G128), .A2(new_n839), .B1(new_n801), .B2(G137), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n371), .B1(new_n835), .B2(G50), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n805), .C2(new_n797), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n792), .A2(new_n777), .B1(new_n776), .B2(new_n215), .ZN(new_n1129));
  OR4_X1    g0929(.A1(new_n279), .A2(new_n1129), .A3(new_n1061), .A4(new_n809), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G97), .A2(new_n822), .B1(new_n801), .B2(G107), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n795), .B2(new_n789), .C1(new_n486), .C2(new_n1008), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1125), .A2(new_n1128), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n755), .B(new_n1120), .C1(new_n1133), .C2(new_n768), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1117), .A2(new_n753), .B1(new_n1119), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1118), .A2(new_n1135), .ZN(G378));
  OAI211_X1 g0936(.A(new_n323), .B(new_n882), .C1(new_n631), .C2(new_n330), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n323), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n337), .B1(new_n1138), .B2(new_n687), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1137), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n936), .A2(G330), .A3(new_n1145), .A4(new_n937), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n937), .B(G330), .C1(new_n935), .C2(KEYINPUT40), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT116), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(new_n921), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(new_n996), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1147), .A2(new_n765), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n371), .A2(new_n501), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n247), .C1(G33), .C2(G41), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n571), .A2(new_n786), .B1(new_n785), .B2(new_n260), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G116), .C2(new_n839), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n781), .A2(G107), .B1(G77), .B2(new_n840), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G58), .A2(new_n835), .B1(new_n790), .B2(G283), .ZN(new_n1160));
  AND4_X1   g0960(.A1(new_n1005), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT114), .Z(new_n1162));
  OAI21_X1  g0962(.A(new_n1156), .B1(new_n1162), .B2(KEYINPUT58), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT115), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n781), .A2(G128), .B1(G132), .B2(new_n801), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n317), .B2(new_n797), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n774), .A2(new_n1124), .ZN(new_n1167));
  INV_X1    g0967(.A(G125), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n792), .A2(new_n1168), .B1(new_n785), .B2(new_n824), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT59), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n835), .A2(G159), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1162), .B2(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n771), .B1(new_n1164), .B2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n755), .B(new_n1178), .C1(new_n247), .C2(new_n820), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1153), .B1(new_n1154), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n664), .A2(new_n869), .A3(new_n1111), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT117), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1116), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT118), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1150), .B2(new_n921), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1150), .A2(new_n921), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1146), .A2(new_n922), .A3(new_n1149), .A4(KEYINPUT118), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1183), .A2(KEYINPUT57), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(KEYINPUT119), .A3(new_n710), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT57), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1183), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n1152), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT119), .B1(new_n1189), .B2(new_n710), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1180), .B1(new_n1194), .B2(new_n1195), .ZN(G375));
  INV_X1    g0996(.A(new_n1110), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1181), .A2(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT120), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT120), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1114), .A2(new_n977), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1110), .A2(new_n753), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT121), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n876), .A2(new_n765), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n755), .B1(new_n215), .B2(new_n820), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT122), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n781), .A2(G137), .B1(G150), .B2(new_n822), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n830), .B2(new_n792), .C1(new_n786), .C2(new_n1124), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G159), .A2(new_n840), .B1(new_n790), .B2(G128), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n371), .B1(new_n835), .B2(G58), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n247), .C2(new_n797), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G116), .A2(new_n801), .B1(new_n790), .B2(G303), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n278), .B2(new_n785), .C1(new_n777), .C2(new_n1008), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G294), .A2(new_n839), .B1(new_n840), .B2(G97), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1040), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(new_n371), .A3(new_n1216), .A4(new_n1002), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1209), .A2(new_n1212), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1207), .B1(new_n768), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1204), .B1(new_n1205), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1202), .A2(new_n1220), .ZN(G381));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1222), .A2(new_n998), .A3(new_n1023), .A4(new_n1223), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1224), .ZN(G407));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n688), .A2(G213), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G375), .C2(new_n1229), .ZN(G409));
  OAI211_X1 g1030(.A(G378), .B(new_n1180), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1192), .A2(new_n1152), .A3(new_n977), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1188), .A2(new_n753), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1154), .A2(new_n1179), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1226), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1231), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1112), .A2(KEYINPUT60), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1199), .A2(new_n1200), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1198), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n711), .B1(new_n1240), .B2(KEYINPUT60), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1220), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n860), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(G384), .A3(new_n1220), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1237), .A2(new_n1227), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT62), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1237), .A2(new_n1227), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1228), .A2(G2897), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1246), .A2(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1244), .A2(G2897), .A3(new_n1228), .A4(new_n1245), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1250), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT62), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1237), .A2(new_n1256), .A3(new_n1227), .A4(new_n1247), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1249), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(G393), .B(G396), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n998), .A2(G390), .A3(new_n1023), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G390), .B1(new_n998), .B2(new_n1023), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G387), .A2(new_n1222), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1260), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n998), .A2(G390), .A3(new_n1023), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1259), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT63), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1246), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1237), .A2(new_n1227), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1237), .A2(new_n1271), .A3(KEYINPUT125), .A4(new_n1227), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1263), .A2(new_n1267), .A3(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1252), .A2(KEYINPUT124), .A3(new_n1253), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT124), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1278), .B1(new_n1250), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT123), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1228), .B(new_n1246), .C1(new_n1231), .C2(new_n1236), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(KEYINPUT63), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1248), .A2(KEYINPUT123), .A3(new_n1270), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1276), .A2(new_n1282), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1269), .A2(new_n1287), .ZN(G405));
  AND2_X1   g1088(.A1(G375), .A2(new_n1226), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1231), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT127), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1247), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1247), .A2(new_n1292), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1246), .A2(KEYINPUT127), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1294), .B(new_n1295), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1268), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1293), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(G402));
endmodule


