//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n452), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(KEYINPUT67), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G137), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n463), .A2(KEYINPUT68), .A3(G101), .A4(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  INV_X1    g051(.A(new_n472), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n463), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(new_n484));
  INV_X1    g059(.A(G2104), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n484), .A2(new_n487), .B1(new_n488), .B2(G136), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n493), .B(new_n494), .C1(new_n472), .C2(new_n471), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n494), .B1(new_n462), .B2(new_n493), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n462), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n463), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G50), .A3(G543), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n507), .B1(G651), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT71), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n505), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n518), .A2(G88), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G166));
  NAND2_X1  g099(.A1(new_n505), .A2(KEYINPUT72), .ZN(new_n525));
  INV_X1    g100(.A(new_n516), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n525), .A2(G543), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n533), .A2(new_n534), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n518), .A2(new_n521), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n531), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AND2_X1   g115(.A1(new_n518), .A2(new_n521), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n530), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(new_n541), .A2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n530), .A2(G43), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n545), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT73), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  AND2_X1   g135(.A1(KEYINPUT74), .A2(G53), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n525), .A2(G543), .A3(new_n529), .A4(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n505), .B2(KEYINPUT72), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n566), .A2(KEYINPUT9), .A3(new_n529), .A4(new_n561), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n518), .A2(G91), .A3(new_n521), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n511), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n564), .A2(new_n567), .A3(new_n568), .A4(new_n572), .ZN(G299));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  INV_X1    g149(.A(new_n522), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n513), .A2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(new_n506), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n574), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n514), .A2(KEYINPUT75), .A3(new_n522), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(G303));
  OAI21_X1  g155(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n541), .A2(G87), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n530), .B2(G49), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n566), .A2(new_n529), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  NOR3_X1   g161(.A1(new_n585), .A2(KEYINPUT76), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n581), .B(new_n582), .C1(new_n584), .C2(new_n587), .ZN(G288));
  NAND3_X1  g163(.A1(new_n505), .A2(G48), .A3(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n541), .B2(G86), .ZN(new_n591));
  OAI21_X1  g166(.A(G61), .B1(new_n509), .B2(new_n510), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(KEYINPUT77), .B1(G73), .B2(G543), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n519), .A2(new_n594), .A3(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n545), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(KEYINPUT78), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n598));
  AOI211_X1 g173(.A(new_n598), .B(new_n545), .C1(new_n593), .C2(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n597), .B2(new_n599), .ZN(G305));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n538), .A2(new_n601), .B1(new_n585), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n511), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n545), .B1(new_n608), .B2(KEYINPUT79), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(KEYINPUT79), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(G290));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NOR2_X1   g187(.A1(G301), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n518), .A2(G92), .A3(new_n521), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G54), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n585), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n530), .A2(KEYINPUT81), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n511), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n618), .A2(new_n619), .B1(G651), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n613), .B1(new_n626), .B2(new_n612), .ZN(G284));
  AOI21_X1  g202(.A(new_n613), .B1(new_n626), .B2(new_n612), .ZN(G321));
  OR3_X1    g203(.A1(G168), .A2(KEYINPUT83), .A3(new_n612), .ZN(new_n629));
  OAI21_X1  g204(.A(KEYINPUT83), .B1(G168), .B2(new_n612), .ZN(new_n630));
  NAND2_X1  g205(.A1(G299), .A2(new_n612), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(G297));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n626), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n553), .A2(new_n612), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n625), .A2(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n481), .A2(G123), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(KEYINPUT84), .ZN(new_n642));
  INV_X1    g217(.A(G111), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n641), .A2(KEYINPUT84), .B1(new_n643), .B2(G2105), .ZN(new_n644));
  AOI22_X1  g219(.A1(G135), .A2(new_n488), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(G2100), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(G2100), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(G2096), .ZN(new_n654));
  NAND4_X1  g229(.A1(new_n647), .A2(new_n652), .A3(new_n653), .A4(new_n654), .ZN(G156));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2430), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT15), .B(G2435), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n660), .B(new_n666), .Z(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n675), .B2(new_n672), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2096), .B(G2100), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n685), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT20), .Z(new_n693));
  AOI211_X1 g268(.A(new_n691), .B(new_n693), .C1(new_n685), .C2(new_n690), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT88), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT87), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NOR2_X1   g278(.A1(G171), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G5), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G1961), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G19), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n554), .B2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n707), .B1(G1341), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G1341), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G32), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n481), .A2(G129), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT26), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n715), .B(new_n717), .C1(G141), .C2(new_n488), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n713), .B1(new_n720), .B2(new_n712), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT94), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT25), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n488), .A2(G139), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n726), .B(new_n727), .C1(new_n463), .C2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G33), .B(new_n729), .S(G29), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2072), .ZN(new_n731));
  INV_X1    g306(.A(G2067), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n712), .A2(G26), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT28), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n481), .A2(G128), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G116), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n488), .B2(G140), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(G29), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n723), .B(new_n731), .C1(new_n732), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n712), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n712), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT29), .Z(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n721), .A2(new_n722), .B1(new_n732), .B2(new_n741), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n712), .A2(G27), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G164), .B2(new_n712), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2078), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(KEYINPUT24), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n712), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G160), .B2(new_n712), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2084), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n748), .A2(new_n751), .A3(new_n757), .ZN(new_n758));
  AND4_X1   g333(.A1(new_n711), .A2(new_n742), .A3(new_n747), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G11), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT97), .B(G28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(new_n712), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n640), .A2(G29), .A3(new_n645), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(KEYINPUT96), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n767), .B1(KEYINPUT96), .B2(new_n766), .C1(new_n705), .C2(new_n706), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n703), .A2(G21), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G168), .B2(new_n703), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT95), .B(G1966), .Z(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n770), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT98), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n703), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT23), .Z(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G299), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1956), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n745), .B2(new_n746), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT99), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n703), .A2(G4), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n626), .B2(new_n703), .ZN(new_n783));
  INV_X1    g358(.A(G1348), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n759), .A2(new_n775), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G23), .B(G288), .S(G16), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT33), .B(G1976), .Z(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n703), .A2(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n703), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1971), .ZN(new_n793));
  OR3_X1    g368(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT32), .B(G1981), .Z(new_n796));
  XOR2_X1   g371(.A(new_n795), .B(new_n796), .Z(new_n797));
  NOR2_X1   g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT34), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT92), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n801), .B(KEYINPUT34), .C1(new_n794), .C2(new_n797), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G290), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT91), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT91), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n703), .B1(G290), .B2(new_n806), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n805), .A2(new_n807), .B1(new_n703), .B2(G24), .ZN(new_n808));
  INV_X1    g383(.A(G1986), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n488), .A2(G131), .ZN(new_n811));
  NOR2_X1   g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT90), .Z(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n481), .A2(G119), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT89), .B1(new_n481), .B2(G119), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n811), .B1(new_n813), .B2(new_n814), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G25), .B(new_n819), .S(G29), .Z(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT35), .B(G1991), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n808), .A2(new_n809), .ZN(new_n823));
  NOR4_X1   g398(.A1(new_n810), .A2(new_n822), .A3(new_n823), .A4(KEYINPUT93), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n798), .A2(new_n799), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n803), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n786), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n828), .A2(KEYINPUT100), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT100), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(G311));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n829), .ZN(G150));
  XOR2_X1   g408(.A(KEYINPUT102), .B(G93), .Z(new_n834));
  AOI22_X1  g409(.A1(new_n541), .A2(new_n834), .B1(new_n530), .B2(G55), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(KEYINPUT101), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(KEYINPUT101), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n837), .A2(G651), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NOR2_X1   g417(.A1(new_n625), .A2(new_n634), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n554), .B(new_n840), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n846), .A2(new_n847), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n842), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(G145));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n719), .B(new_n740), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n729), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n496), .B2(new_n497), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n493), .B1(new_n471), .B2(new_n472), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT4), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n861), .A2(KEYINPUT104), .A3(new_n495), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n503), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n857), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n819), .B(new_n649), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n481), .A2(G130), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G118), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n867), .A2(new_n868), .B1(new_n870), .B2(G2105), .ZN(new_n871));
  AOI22_X1  g446(.A1(G142), .A2(new_n488), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n865), .B(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT106), .B1(new_n864), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n865), .B(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n857), .A2(new_n863), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n857), .A2(new_n863), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n877), .A2(KEYINPUT106), .A3(new_n878), .A4(new_n879), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n490), .B(new_n646), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G160), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n864), .B2(new_n875), .ZN(new_n887));
  AOI21_X1  g462(.A(G37), .B1(new_n887), .B2(new_n880), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n886), .B1(new_n885), .B2(new_n888), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n855), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(KEYINPUT40), .A3(new_n889), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n892), .A2(new_n894), .ZN(G395));
  XNOR2_X1  g470(.A(G290), .B(new_n523), .ZN(new_n896));
  XOR2_X1   g471(.A(G305), .B(G288), .Z(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(KEYINPUT109), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(KEYINPUT109), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n624), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(G299), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT108), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(G299), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n904), .A2(KEYINPUT108), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT41), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n904), .A2(KEYINPUT108), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n906), .A4(new_n905), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n840), .B(new_n553), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n637), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n637), .A2(new_n913), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n909), .B(new_n912), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n910), .A2(new_n906), .A3(new_n905), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n914), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n902), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n902), .A3(new_n920), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n900), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n923), .ZN(new_n925));
  INV_X1    g500(.A(new_n900), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n925), .A2(new_n926), .A3(new_n921), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n840), .A2(new_n612), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n926), .B1(new_n925), .B2(new_n921), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n922), .A2(new_n900), .A3(new_n923), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n612), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n930), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT110), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n928), .A2(new_n930), .ZN(G331));
  XNOR2_X1  g513(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n939));
  OR2_X1    g514(.A1(G171), .A2(KEYINPUT112), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n845), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G286), .B1(G171), .B2(KEYINPUT112), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n913), .B(new_n940), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n942), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n946), .A3(new_n919), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n945), .B(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n909), .A2(new_n912), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n898), .ZN(new_n951));
  INV_X1    g526(.A(new_n898), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(new_n947), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n951), .A2(new_n953), .A3(new_n957), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n939), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n939), .ZN(new_n962));
  AOI211_X1 g537(.A(KEYINPUT111), .B(new_n962), .C1(new_n956), .C2(new_n958), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(G1956), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n501), .A2(new_n502), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n479), .B2(G126), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n861), .A2(KEYINPUT104), .A3(new_n495), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT104), .B1(new_n861), .B2(new_n495), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G40), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n470), .A2(new_n475), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n498), .B2(new_n503), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n965), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n568), .A2(new_n567), .A3(new_n572), .ZN(new_n979));
  NOR2_X1   g554(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n979), .A2(new_n564), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(G299), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n971), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n985));
  INV_X1    g560(.A(new_n475), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n986), .A2(G40), .A3(new_n464), .A4(new_n469), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(new_n976), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT56), .B(G2072), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n985), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n978), .A2(new_n983), .A3(new_n984), .A4(new_n991), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n978), .A2(new_n991), .B1(new_n983), .B2(new_n984), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n863), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n861), .A2(new_n495), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n995), .B2(new_n968), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n975), .B1(new_n996), .B2(new_n966), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n784), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n863), .A2(G1384), .A3(new_n987), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n732), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n624), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n992), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT61), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n985), .A2(new_n989), .A3(new_n990), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT50), .B1(new_n863), .B2(G1384), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n987), .B1(new_n996), .B2(new_n966), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1956), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n983), .A2(new_n984), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1003), .B1(new_n1009), .B2(new_n993), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT121), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT121), .B(new_n1003), .C1(new_n1009), .C2(new_n993), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n985), .A2(new_n989), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT58), .B(G1341), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n1015), .A2(G1996), .B1(new_n999), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n554), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT59), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1020), .A3(new_n554), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n998), .A2(KEYINPUT60), .A3(new_n1000), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n624), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n998), .A2(new_n1000), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT60), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n903), .A2(new_n998), .A3(KEYINPUT60), .A4(new_n1000), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n993), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n992), .A3(KEYINPUT61), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1022), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1002), .B1(new_n1014), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT122), .B(new_n1002), .C1(new_n1014), .C2(new_n1032), .ZN(new_n1036));
  INV_X1    g611(.A(G2078), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n985), .A2(new_n989), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n706), .B1(new_n994), .B2(new_n997), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n988), .B1(new_n863), .B2(G1384), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n987), .B1(new_n996), .B2(KEYINPUT45), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1039), .A2(G2078), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1041), .A2(KEYINPUT125), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT125), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G171), .ZN(new_n1049));
  AOI21_X1  g624(.A(G171), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n863), .B2(G1384), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n971), .A2(new_n1052), .A3(new_n972), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1053), .A3(new_n988), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n975), .A2(new_n1044), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n863), .A2(G1384), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(KEYINPUT45), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(new_n1041), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT54), .B1(new_n1049), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1050), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G171), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(KEYINPUT54), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  INV_X1    g641(.A(G8), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT45), .B1(new_n971), .B2(new_n972), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n975), .B1(new_n976), .B2(new_n988), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n771), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n971), .A2(new_n966), .A3(new_n972), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n987), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n1072));
  INV_X1    g647(.A(G2084), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1067), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G286), .A2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(G286), .A2(KEYINPUT123), .A3(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1065), .B(new_n1066), .C1(new_n1075), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1074), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n772), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1083));
  OAI21_X1  g658(.A(G8), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1078), .A2(new_n1079), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1081), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1064), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1971), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1015), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1005), .A2(new_n746), .A3(new_n1006), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1067), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n994), .A2(G2090), .A3(new_n997), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1971), .B1(new_n985), .B2(new_n989), .ZN(new_n1097));
  OAI21_X1  g672(.A(G8), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n578), .A2(G8), .A3(new_n579), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n578), .A2(KEYINPUT55), .A3(new_n579), .A4(G8), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  MUX2_X1   g678(.A(new_n1095), .B(new_n1098), .S(new_n1103), .Z(new_n1104));
  INV_X1    g679(.A(G1976), .ZN(new_n1105));
  OR2_X1    g680(.A1(G288), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT52), .B1(G288), .B2(new_n1105), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n971), .A2(new_n972), .A3(new_n975), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT116), .B1(new_n1108), .B2(G8), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1106), .B(new_n1107), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n999), .B2(new_n1067), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1109), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1117), .A2(KEYINPUT117), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G1981), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n591), .B(new_n1120), .C1(new_n597), .C2(new_n599), .ZN(new_n1121));
  INV_X1    g696(.A(G86), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n589), .B1(new_n538), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(G1981), .B1(new_n1123), .B2(new_n596), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT118), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1126), .A2(KEYINPUT49), .B1(new_n1116), .B2(new_n1109), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT49), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(KEYINPUT118), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1127), .A2(new_n1129), .B1(new_n1130), .B2(KEYINPUT52), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1104), .A2(new_n1119), .A3(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1060), .A2(new_n1091), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1035), .A2(new_n1036), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1084), .A2(G286), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1104), .A2(new_n1119), .A3(new_n1131), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT119), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1140), .A3(new_n1137), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1119), .A2(new_n1131), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1103), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1098), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(new_n1137), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1098), .A2(new_n1143), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1142), .A2(new_n1135), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1139), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1149));
  OR2_X1    g724(.A1(G288), .A2(G1976), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1121), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1142), .A2(new_n1144), .B1(new_n1151), .B2(new_n1117), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1134), .A2(new_n1148), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1134), .A2(new_n1148), .A3(KEYINPUT126), .A4(new_n1152), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1090), .A2(KEYINPUT62), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT127), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1132), .A2(new_n1049), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1158), .B(new_n1159), .C1(KEYINPUT62), .C2(new_n1090), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1155), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1054), .A2(new_n987), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT115), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n740), .A2(G2067), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n735), .A2(new_n732), .A3(new_n739), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(G1996), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(new_n720), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1162), .A2(G1996), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1163), .A2(new_n1168), .B1(new_n720), .B2(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n819), .A2(new_n821), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n819), .A2(new_n821), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1163), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n804), .A2(new_n809), .ZN(new_n1175));
  NAND2_X1  g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1162), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1161), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1163), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(new_n1165), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1169), .B(KEYINPUT46), .Z(new_n1183));
  INV_X1    g758(.A(new_n1166), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1163), .B1(new_n719), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT47), .Z(new_n1187));
  INV_X1    g762(.A(new_n1174), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1175), .A2(new_n1162), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT48), .Z(new_n1190));
  AOI211_X1 g765(.A(new_n1182), .B(new_n1187), .C1(new_n1188), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1179), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g767(.A1(new_n893), .A2(new_n889), .ZN(new_n1194));
  NOR4_X1   g768(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n1194), .A2(new_n959), .A3(new_n1195), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


