//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT65), .B1(new_n187), .B2(G146), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n190), .B2(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n187), .A2(KEYINPUT66), .A3(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  AND4_X1   g011(.A1(new_n192), .A2(new_n194), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n187), .A2(G146), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT64), .B1(new_n190), .B2(G143), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(new_n187), .A3(G146), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT0), .B(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  AOI22_X1  g022(.A1(KEYINPUT68), .A2(new_n207), .B1(new_n208), .B2(G137), .ZN(new_n209));
  OAI22_X1  g023(.A1(KEYINPUT68), .A2(new_n207), .B1(new_n208), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT11), .A4(G134), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n209), .A2(new_n210), .A3(new_n216), .A4(new_n213), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n215), .A2(KEYINPUT70), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT70), .B1(new_n215), .B2(new_n217), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n206), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n212), .A2(KEYINPUT69), .A3(G134), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n212), .B2(G134), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n208), .A2(G137), .ZN(new_n224));
  OAI211_X1 g038(.A(G131), .B(new_n221), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  OAI21_X1  g041(.A(G128), .B1(new_n199), .B2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n200), .A2(new_n202), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n199), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n192), .A2(new_n194), .A3(new_n195), .A4(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n226), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n220), .A2(KEYINPUT30), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT2), .A2(G113), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT2), .A2(G113), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n241), .B(new_n244), .Z(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n247));
  OAI22_X1  g061(.A1(new_n247), .A2(new_n196), .B1(new_n203), .B2(new_n204), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n248), .A2(new_n249), .B1(new_n217), .B2(new_n215), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n206), .A2(KEYINPUT67), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n234), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n236), .B(new_n246), .C1(KEYINPUT30), .C2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT31), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(G101), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n220), .A2(new_n245), .A3(new_n235), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n253), .A2(new_n254), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n253), .A2(new_n259), .A3(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT31), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n262), .A3(KEYINPUT31), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n260), .A2(KEYINPUT28), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n260), .A2(KEYINPUT28), .ZN(new_n269));
  OAI22_X1  g083(.A1(new_n268), .A2(new_n269), .B1(new_n245), .B2(new_n252), .ZN(new_n270));
  INV_X1    g084(.A(new_n259), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(G472), .A2(G902), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT72), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n273), .A2(KEYINPUT32), .A3(new_n276), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n220), .A2(new_n235), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(new_n246), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n268), .B2(new_n269), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n260), .A2(KEYINPUT73), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n271), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n253), .A2(new_n260), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n271), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n291), .B(new_n287), .C1(new_n271), .C2(new_n270), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G472), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n279), .A2(new_n280), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n280), .A4(new_n294), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  INV_X1    g114(.A(G953), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(G221), .A3(G234), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT79), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT22), .B(G137), .Z(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G125), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(KEYINPUT16), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT16), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n308), .B1(new_n311), .B2(KEYINPUT77), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n307), .A2(new_n313), .A3(KEYINPUT16), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n190), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n314), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n317), .B2(KEYINPUT16), .ZN(new_n318));
  OAI211_X1 g132(.A(G146), .B(new_n316), .C1(new_n318), .C2(new_n308), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n319), .A3(KEYINPUT78), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n321), .B(new_n190), .C1(new_n312), .C2(new_n314), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(G119), .B2(new_n231), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n237), .A2(KEYINPUT23), .A3(G128), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n324), .A2(new_n325), .B1(G119), .B2(new_n231), .ZN(new_n326));
  XNOR2_X1  g140(.A(G119), .B(G128), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT24), .B(G110), .Z(new_n328));
  AOI22_X1  g142(.A1(new_n326), .A2(G110), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n320), .A2(new_n322), .A3(new_n329), .ZN(new_n330));
  OAI22_X1  g144(.A1(new_n326), .A2(G110), .B1(new_n327), .B2(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n317), .A2(new_n190), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n319), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n305), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(KEYINPUT80), .A3(new_n333), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n300), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(KEYINPUT81), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(KEYINPUT81), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT75), .B(G217), .ZN(new_n347));
  INV_X1    g161(.A(G234), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(G902), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT76), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n340), .B2(new_n343), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n338), .A2(new_n339), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n300), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n346), .A2(new_n352), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G113), .B(G122), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT92), .B(G104), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n301), .A3(G214), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT91), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G143), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(G143), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n187), .A2(KEYINPUT91), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G214), .A4(new_n255), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT18), .A3(G131), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(new_n368), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT18), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n317), .B(new_n190), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n216), .ZN(new_n375));
  AND4_X1   g189(.A1(new_n370), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n365), .A2(new_n368), .A3(G131), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n317), .B(KEYINPUT19), .Z(new_n380));
  OAI211_X1 g194(.A(new_n379), .B(new_n319), .C1(G146), .C2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n361), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT17), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n375), .A2(new_n383), .A3(new_n378), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n369), .A2(KEYINPUT93), .A3(KEYINPUT17), .A4(G131), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT93), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n378), .B2(new_n383), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n320), .A2(new_n322), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n361), .A3(new_n377), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT94), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n376), .B1(new_n388), .B2(new_n389), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT94), .A3(new_n361), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n382), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(G475), .A2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(KEYINPUT20), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n382), .ZN(new_n400));
  AND4_X1   g214(.A1(KEYINPUT94), .A2(new_n390), .A3(new_n361), .A4(new_n377), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT94), .B1(new_n394), .B2(new_n361), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n397), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n394), .A2(new_n361), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n393), .B2(new_n395), .ZN(new_n409));
  OAI21_X1  g223(.A(G475), .B1(new_n409), .B2(G902), .ZN(new_n410));
  OAI211_X1 g224(.A(G952), .B(new_n301), .C1(new_n348), .C2(new_n362), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT95), .ZN(new_n412));
  OAI211_X1 g226(.A(G902), .B(G953), .C1(new_n348), .C2(new_n362), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT96), .Z(new_n414));
  XOR2_X1   g228(.A(KEYINPUT21), .B(G898), .Z(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G116), .B(G122), .ZN(new_n417));
  INV_X1    g231(.A(G107), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(KEYINPUT14), .A2(G107), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n239), .B2(G122), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n420), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n187), .A2(G128), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n231), .A2(G143), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(G134), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n422), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT13), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n208), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n430), .A2(new_n426), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n426), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n419), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT9), .B(G234), .Z(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n301), .A3(new_n347), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n428), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n300), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n441), .A2(new_n443), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n410), .A2(new_n416), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT97), .B1(new_n407), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n410), .A2(new_n446), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT97), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n406), .A4(new_n416), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G221), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n435), .B2(new_n300), .ZN(new_n454));
  INV_X1    g268(.A(G104), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n455), .A2(KEYINPUT3), .A3(G107), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(KEYINPUT82), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G104), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n456), .B1(new_n460), .B2(G107), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n459), .A3(new_n418), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT83), .B(G101), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n463), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n465), .A2(KEYINPUT4), .B1(new_n466), .B2(G101), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(KEYINPUT4), .A3(G101), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n206), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OR3_X1    g284(.A1(new_n418), .A2(KEYINPUT84), .A3(G104), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT84), .B1(new_n418), .B2(G104), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n462), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n247), .A2(new_n228), .ZN(new_n475));
  INV_X1    g289(.A(new_n233), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n465), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT10), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n218), .A2(new_n219), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n465), .A2(new_n474), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n230), .A2(new_n233), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(KEYINPUT10), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n470), .A2(new_n479), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G110), .B(G140), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n301), .A2(G227), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n485), .B(new_n486), .Z(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n477), .B1(new_n482), .B2(new_n481), .ZN(new_n492));
  INV_X1    g306(.A(new_n480), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT12), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n215), .A2(new_n217), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n495), .A2(KEYINPUT12), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n489), .B(new_n491), .C1(new_n494), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n470), .A2(new_n479), .A3(new_n483), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n493), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n484), .ZN(new_n501));
  INV_X1    g315(.A(new_n487), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G469), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n300), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n484), .B1(new_n497), .B2(new_n494), .ZN(new_n507));
  INV_X1    g321(.A(new_n488), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n507), .A2(new_n502), .B1(new_n508), .B2(new_n500), .ZN(new_n509));
  OAI21_X1  g323(.A(G469), .B1(new_n509), .B2(G902), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n454), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G214), .B1(G237), .B2(G902), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT86), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n465), .A2(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n466), .A2(G101), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n245), .B1(new_n517), .B2(new_n468), .ZN(new_n518));
  INV_X1    g332(.A(G113), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n239), .A2(G119), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT5), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT5), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n522), .A2(new_n523), .B1(new_n241), .B2(new_n244), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n465), .A2(new_n474), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n514), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n246), .B1(new_n467), .B2(new_n469), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT86), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n513), .B(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n525), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(KEYINPUT87), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n526), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G125), .B1(new_n198), .B2(new_n205), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n230), .A2(new_n309), .A3(new_n233), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT88), .B(G224), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G953), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n537), .B(new_n539), .ZN(new_n540));
  OAI221_X1 g354(.A(new_n514), .B1(KEYINPUT87), .B2(new_n532), .C1(new_n518), .C2(new_n525), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n529), .A2(KEYINPUT8), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n514), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n524), .B1(new_n465), .B2(new_n474), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(new_n525), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n539), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT7), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(KEYINPUT7), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI211_X1 g367(.A(KEYINPUT89), .B(new_n553), .C1(new_n535), .C2(new_n536), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT89), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n537), .B2(new_n552), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(G902), .B1(new_n557), .B2(new_n531), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n542), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G210), .B1(G237), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT90), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n542), .A2(new_n558), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n562), .A3(new_n561), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n511), .A2(new_n512), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n452), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n299), .A2(new_n357), .A3(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n570), .B(new_n464), .Z(G3));
  NAND2_X1  g385(.A1(new_n511), .A2(new_n357), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n273), .A2(new_n300), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G472), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n277), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n542), .A2(new_n558), .A3(new_n560), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT98), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n565), .A2(new_n561), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT98), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n542), .A2(new_n558), .A3(new_n579), .A4(new_n560), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n512), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n572), .A2(new_n575), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n437), .A2(KEYINPUT100), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n439), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n428), .A2(KEYINPUT100), .A3(new_n433), .A4(new_n438), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(KEYINPUT33), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n588));
  NAND2_X1  g402(.A1(new_n440), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n442), .A2(G902), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n591), .A2(KEYINPUT101), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(KEYINPUT101), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n441), .A2(new_n442), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n396), .A2(KEYINPUT20), .A3(new_n398), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n404), .B1(new_n403), .B2(new_n397), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n410), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n416), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n583), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  OR2_X1    g418(.A1(new_n406), .A2(KEYINPUT102), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n597), .A2(KEYINPUT102), .ZN(new_n606));
  INV_X1    g420(.A(new_n446), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(new_n410), .ZN(new_n608));
  AND4_X1   g422(.A1(new_n416), .A2(new_n605), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n583), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  XNOR2_X1  g426(.A(new_n334), .B(KEYINPUT103), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n305), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n346), .A2(new_n352), .B1(new_n356), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n575), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n569), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT37), .B(G110), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G12));
  INV_X1    g434(.A(new_n582), .ZN(new_n621));
  INV_X1    g435(.A(new_n616), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n412), .B1(new_n414), .B2(G900), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n605), .A2(new_n606), .A3(new_n608), .A4(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n506), .A2(new_n510), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n624), .A2(new_n454), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n299), .A2(new_n621), .A3(new_n622), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G128), .ZN(G30));
  INV_X1    g442(.A(new_n567), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT38), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n446), .B1(new_n406), .B2(new_n410), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n567), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n630), .A2(new_n512), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n623), .B(KEYINPUT39), .Z(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n511), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n634), .B1(KEYINPUT40), .B2(new_n637), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n263), .A2(new_n265), .B1(new_n271), .B2(new_n270), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n278), .B(new_n275), .C1(new_n639), .C2(new_n267), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT32), .B1(new_n273), .B2(new_n276), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n290), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n271), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n283), .A2(new_n271), .A3(new_n260), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n300), .A3(new_n285), .ZN(new_n646));
  OAI21_X1  g460(.A(G472), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n622), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n638), .B(new_n648), .C1(KEYINPUT40), .C2(new_n637), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G143), .ZN(G45));
  INV_X1    g464(.A(new_n599), .ZN(new_n651));
  INV_X1    g465(.A(new_n623), .ZN(new_n652));
  AOI211_X1 g466(.A(new_n454), .B(new_n652), .C1(new_n506), .C2(new_n510), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n299), .A2(new_n621), .A3(new_n622), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G146), .ZN(G48));
  AOI21_X1  g470(.A(G902), .B1(new_n498), .B2(new_n503), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G469), .ZN(new_n658));
  INV_X1    g472(.A(new_n454), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n621), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT74), .B1(new_n642), .B2(new_n294), .ZN(new_n662));
  INV_X1    g476(.A(new_n298), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n357), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n601), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT104), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n357), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n297), .B2(new_n298), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n601), .A4(new_n661), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NAND4_X1  g487(.A1(new_n299), .A2(new_n357), .A3(new_n609), .A4(new_n661), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  NOR2_X1   g489(.A1(new_n660), .A2(new_n452), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n299), .A2(new_n676), .A3(new_n622), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  OAI211_X1 g492(.A(new_n265), .B(new_n261), .C1(new_n286), .C2(new_n259), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n276), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n574), .A2(new_n357), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n658), .A2(new_n659), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n681), .A2(new_n682), .A3(new_n600), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n581), .A2(new_n598), .A3(new_n607), .A4(new_n512), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n631), .A2(new_n686), .A3(new_n512), .A4(new_n581), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G122), .ZN(G24));
  NAND3_X1  g504(.A1(new_n622), .A2(new_n574), .A3(new_n680), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n599), .A2(new_n652), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n661), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  NAND2_X1  g509(.A1(new_n693), .A2(KEYINPUT42), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n295), .A2(new_n357), .ZN(new_n697));
  INV_X1    g511(.A(new_n512), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n567), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n511), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n696), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n700), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n668), .A2(new_n693), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n216), .ZN(G33));
  INV_X1    g520(.A(new_n668), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n707), .A2(new_n624), .A3(new_n700), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n208), .ZN(G36));
  NAND2_X1  g523(.A1(new_n507), .A2(new_n502), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n508), .A2(new_n500), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT107), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n505), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n509), .A2(new_n716), .A3(KEYINPUT45), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(G469), .A2(G902), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n718), .A2(KEYINPUT46), .A3(new_n719), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n506), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n659), .A3(new_n636), .A4(new_n699), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n598), .A3(KEYINPUT43), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n598), .A2(KEYINPUT108), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n598), .A2(KEYINPUT108), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n595), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n727), .B1(new_n730), .B2(KEYINPUT43), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n575), .A2(new_n732), .A3(new_n622), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n732), .B1(new_n575), .B2(new_n622), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n725), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n731), .B(KEYINPUT44), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G137), .ZN(G39));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n723), .A2(new_n506), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT46), .B1(new_n718), .B2(new_n719), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n742), .B(new_n659), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n742), .B1(new_n724), .B2(new_n659), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n693), .A2(new_n667), .A3(new_n699), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n299), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G140), .ZN(G42));
  INV_X1    g566(.A(KEYINPUT121), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n658), .A2(new_n699), .A3(new_n659), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n412), .B1(new_n754), .B2(KEYINPUT117), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n658), .A2(new_n699), .A3(new_n756), .A4(new_n659), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n731), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n697), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT48), .Z(new_n760));
  INV_X1    g574(.A(new_n682), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n681), .A2(new_n412), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n731), .A2(new_n621), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n301), .A2(G952), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT120), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n755), .A2(new_n757), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n642), .A2(new_n357), .A3(new_n647), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n651), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n760), .A2(new_n763), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n731), .A2(new_n699), .A3(new_n762), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n724), .A2(new_n659), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT47), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n745), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n658), .A2(new_n454), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n630), .A2(new_n633), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n512), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n731), .A3(new_n761), .A4(new_n762), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT50), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT50), .B1(new_n779), .B2(new_n780), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n776), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n755), .A2(new_n757), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(KEYINPUT118), .A3(new_n692), .A4(new_n731), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n758), .B2(new_n691), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n598), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n768), .A2(new_n790), .A3(new_n726), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(KEYINPUT119), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT119), .B1(new_n789), .B2(new_n791), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n784), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT51), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n748), .A2(KEYINPUT115), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n748), .A2(KEYINPUT115), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n798), .A3(new_n775), .ZN(new_n799));
  INV_X1    g613(.A(new_n771), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n782), .A2(new_n783), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n789), .A2(new_n803), .A3(new_n791), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n753), .B(new_n770), .C1(new_n796), .C2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n783), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n774), .A2(new_n775), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n781), .B(new_n808), .C1(new_n809), .C2(new_n771), .ZN(new_n810));
  INV_X1    g624(.A(new_n794), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n810), .B1(new_n811), .B2(new_n792), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n806), .B1(new_n812), .B2(new_n803), .ZN(new_n813));
  INV_X1    g627(.A(new_n770), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT121), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n807), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n572), .A2(new_n575), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n567), .A2(new_n416), .A3(new_n512), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n790), .A2(new_n607), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n819), .B2(new_n599), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n569), .A2(new_n617), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n570), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n449), .A2(new_n605), .A3(new_n606), .A4(new_n623), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n622), .B(new_n824), .C1(new_n662), .C2(new_n663), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n692), .A2(new_n693), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n700), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n705), .A2(new_n708), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n674), .A2(new_n677), .A3(new_n689), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n671), .A2(new_n829), .A3(KEYINPUT110), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT110), .B1(new_n671), .B2(new_n829), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n823), .B(new_n828), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n627), .A2(new_n655), .A3(new_n694), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n685), .A2(new_n687), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n279), .A2(new_n280), .A3(new_n647), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n616), .A3(new_n653), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n836), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n648), .A2(new_n688), .A3(KEYINPUT111), .A4(new_n653), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n834), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n693), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n844), .A2(new_n691), .A3(new_n660), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n582), .B(new_n616), .C1(new_n297), .C2(new_n298), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n846), .B2(new_n626), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n840), .A2(new_n841), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(KEYINPUT112), .A3(new_n655), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n843), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n850), .B1(new_n843), .B2(new_n849), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n833), .A2(new_n854), .A3(KEYINPUT53), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT52), .B1(new_n835), .B2(new_n842), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n856), .B(new_n857), .C1(new_n832), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n671), .A2(new_n829), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT110), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n671), .A2(new_n829), .A3(KEYINPUT110), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n822), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n828), .A3(new_n851), .A4(new_n858), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n856), .B1(new_n867), .B2(new_n857), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n627), .A2(new_n655), .A3(new_n694), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT112), .B1(new_n871), .B2(new_n848), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n835), .A2(new_n842), .A3(new_n834), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT52), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n851), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n875), .A2(new_n832), .A3(KEYINPUT53), .ZN(new_n876));
  INV_X1    g690(.A(new_n827), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n671), .A2(new_n829), .A3(new_n877), .A4(new_n823), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n705), .A2(new_n708), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n851), .A2(new_n878), .A3(new_n879), .A4(new_n858), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(KEYINPUT53), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n870), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(KEYINPUT114), .B(new_n870), .C1(new_n876), .C2(new_n881), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n816), .A2(new_n869), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(G952), .A2(G953), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n777), .A2(new_n454), .A3(new_n698), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n658), .B(KEYINPUT49), .Z(new_n890));
  OR4_X1    g704(.A1(new_n730), .A2(new_n889), .A3(new_n767), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n301), .A2(G952), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n833), .A2(new_n854), .A3(new_n857), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n880), .A2(KEYINPUT53), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(G210), .A3(G902), .A4(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(KEYINPUT122), .A2(KEYINPUT123), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n534), .A2(new_n541), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(new_n540), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT55), .Z(new_n901));
  AND2_X1   g715(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n898), .B1(new_n902), .B2(KEYINPUT122), .ZN(new_n903));
  NOR2_X1   g717(.A1(KEYINPUT123), .A2(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n901), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n893), .B1(new_n903), .B2(new_n907), .ZN(G51));
  XOR2_X1   g722(.A(new_n719), .B(KEYINPUT57), .Z(new_n909));
  NOR3_X1   g723(.A1(new_n876), .A2(new_n881), .A3(new_n870), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT54), .B1(new_n894), .B2(new_n895), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n504), .ZN(new_n913));
  OR4_X1    g727(.A1(new_n300), .A2(new_n876), .A3(new_n881), .A4(new_n718), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n893), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NOR2_X1   g729(.A1(new_n876), .A2(new_n881), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n917), .A2(new_n396), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n396), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n893), .ZN(G60));
  NAND2_X1  g734(.A1(new_n587), .A2(new_n589), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT59), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n922), .B(new_n924), .C1(new_n910), .C2(new_n911), .ZN(new_n925));
  INV_X1    g739(.A(new_n893), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n869), .A2(new_n884), .A3(new_n885), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n924), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n929), .B2(new_n921), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT60), .Z(new_n932));
  NAND3_X1  g746(.A1(new_n894), .A2(new_n895), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n615), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n926), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n354), .B1(new_n916), .B2(new_n932), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(G66));
  INV_X1    g754(.A(new_n538), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n301), .B1(new_n941), .B2(new_n415), .ZN(new_n942));
  INV_X1    g756(.A(new_n866), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n301), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n899), .B1(G898), .B2(new_n301), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n944), .B(new_n945), .Z(G69));
  MUX2_X1   g760(.A(new_n252), .B(new_n282), .S(KEYINPUT30), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n380), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n649), .A2(new_n627), .A3(new_n655), .A4(new_n694), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AOI22_X1  g765(.A1(new_n738), .A2(new_n739), .B1(new_n748), .B2(new_n750), .ZN(new_n952));
  INV_X1    g766(.A(new_n699), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n953), .B(new_n637), .C1(new_n599), .C2(new_n819), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n668), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n951), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n951), .B2(new_n956), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n948), .B1(new_n960), .B2(G953), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n301), .B1(G227), .B2(G900), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n964));
  OR4_X1    g778(.A1(new_n635), .A2(new_n772), .A3(new_n837), .A4(new_n697), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n879), .A2(new_n952), .A3(new_n871), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n301), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n301), .A2(G900), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n964), .A3(new_n969), .ZN(new_n971));
  INV_X1    g785(.A(new_n948), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n961), .B(new_n963), .C1(new_n970), .C2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n973), .B2(new_n970), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n967), .A2(new_n969), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT125), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n978), .A2(KEYINPUT126), .A3(new_n972), .A4(new_n971), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n976), .A2(new_n961), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n980), .A2(new_n981), .A3(new_n962), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n980), .B2(new_n962), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n974), .B1(new_n982), .B2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n943), .B2(new_n966), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n290), .A2(new_n259), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n893), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n986), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n960), .B2(new_n866), .ZN(new_n991));
  INV_X1    g805(.A(new_n644), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n861), .A2(new_n868), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n291), .B2(new_n264), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(G57));
endmodule


