//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G134), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n190), .B1(new_n195), .B2(new_n188), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT66), .B1(new_n198), .B2(new_n194), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n192), .A2(G134), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(G137), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n196), .A2(new_n197), .A3(new_n199), .A4(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n195), .B1(G134), .B2(new_n194), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT1), .A3(G146), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n212), .B(new_n214), .C1(G128), .C2(new_n209), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n204), .A2(new_n216), .A3(new_n206), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n208), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT30), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n195), .A2(new_n188), .ZN(new_n220));
  INV_X1    g034(.A(new_n190), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n199), .A2(new_n220), .A3(new_n221), .A4(new_n203), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n204), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n213), .A2(G146), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G143), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n209), .A2(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n224), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n218), .A2(new_n219), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n234), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n223), .B2(new_n204), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n204), .A2(new_n215), .A3(new_n206), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT30), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT2), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G116), .ZN(new_n249));
  INV_X1    g063(.A(G119), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n249), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n250), .A2(G116), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n248), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n255), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT68), .B(G119), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n247), .B(new_n257), .C1(new_n258), .C2(new_n249), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n242), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n191), .A2(new_n193), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n200), .B1(new_n262), .B2(G137), .ZN(new_n263));
  AOI211_X1 g077(.A(KEYINPUT66), .B(new_n194), .C1(new_n191), .C2(new_n193), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n197), .B1(new_n265), .B2(new_n196), .ZN(new_n266));
  INV_X1    g080(.A(new_n204), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n234), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n260), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n204), .A2(new_n215), .A3(new_n206), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT26), .B(G101), .Z(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(G237), .A2(G953), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G210), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT70), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n277), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n239), .A2(new_n240), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(new_n269), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n261), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n242), .A2(new_n260), .B1(KEYINPUT70), .B2(new_n282), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT31), .A3(new_n279), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n269), .B1(new_n218), .B2(new_n236), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n271), .B1(new_n289), .B2(KEYINPUT71), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n291), .B(new_n269), .C1(new_n218), .C2(new_n236), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT28), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n239), .A2(new_n240), .A3(new_n260), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(KEYINPUT28), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n286), .A2(new_n288), .B1(new_n297), .B2(new_n280), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n187), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n260), .B1(new_n239), .B2(new_n240), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n271), .A2(new_n302), .A3(KEYINPUT72), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n281), .A2(new_n304), .A3(new_n269), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(KEYINPUT28), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n280), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n296), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT73), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n313), .A3(new_n310), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n294), .B1(new_n242), .B2(new_n260), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n307), .B1(new_n316), .B2(new_n277), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n204), .A2(new_n216), .A3(new_n206), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n216), .B1(new_n204), .B2(new_n206), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n211), .A2(new_n225), .A3(new_n227), .ZN(new_n320));
  AOI21_X1  g134(.A(G128), .B1(new_n225), .B2(new_n227), .ZN(new_n321));
  INV_X1    g135(.A(new_n214), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n318), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n224), .A2(new_n235), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n260), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n291), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n271), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n295), .B1(new_n329), .B2(KEYINPUT28), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n317), .B1(new_n330), .B2(new_n277), .ZN(new_n331));
  OAI21_X1  g145(.A(G472), .B1(new_n315), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT31), .B1(new_n287), .B2(new_n279), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n269), .B1(new_n237), .B2(new_n241), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n271), .A2(KEYINPUT70), .A3(new_n277), .ZN(new_n335));
  NOR4_X1   g149(.A1(new_n334), .A2(new_n335), .A3(new_n278), .A4(new_n285), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n330), .A2(new_n277), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(KEYINPUT32), .A3(new_n299), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n301), .A2(new_n332), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(G214), .B1(G237), .B2(G902), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n340), .B(KEYINPUT82), .Z(new_n341));
  INV_X1    g155(.A(G104), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT3), .B1(new_n342), .B2(G107), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n344));
  INV_X1    g158(.A(G107), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(G107), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G101), .ZN(new_n349));
  INV_X1    g163(.A(G101), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n343), .A2(new_n346), .A3(new_n350), .A4(new_n347), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(KEYINPUT4), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n353), .A3(G101), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n260), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT5), .B(new_n257), .C1(new_n258), .C2(new_n249), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n254), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n358), .A3(G113), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n345), .A2(G104), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n342), .A2(G107), .ZN(new_n361));
  OAI21_X1  g175(.A(G101), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n259), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT83), .B1(new_n355), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(G110), .B(G122), .Z(new_n367));
  NAND3_X1  g181(.A1(new_n355), .A2(new_n364), .A3(KEYINPUT83), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n366), .A2(KEYINPUT6), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n355), .A2(new_n364), .A3(KEYINPUT83), .ZN(new_n370));
  INV_X1    g184(.A(new_n367), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n370), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n355), .A2(new_n364), .A3(new_n371), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n373), .A2(KEYINPUT6), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n369), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G125), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT84), .B1(new_n234), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n232), .A2(new_n233), .A3(new_n378), .A4(G125), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n323), .A2(new_n376), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G953), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G224), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT85), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n382), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT86), .ZN(new_n388));
  AOI211_X1 g202(.A(KEYINPUT5), .B(new_n249), .C1(new_n251), .C2(new_n253), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(new_n243), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n358), .A2(KEYINPUT86), .A3(G113), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n356), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n392), .A2(new_n393), .A3(new_n259), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n392), .B2(new_n259), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n363), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n367), .A2(KEYINPUT8), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n367), .A2(KEYINPUT8), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n359), .A2(new_n259), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n351), .A2(new_n362), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n381), .B1(new_n376), .B2(new_n234), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT7), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n385), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n385), .A2(new_n404), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n380), .A2(new_n381), .A3(new_n406), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n405), .A2(new_n373), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(G902), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n387), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G210), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n387), .A2(new_n409), .A3(new_n411), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n341), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G140), .B1(new_n376), .B2(KEYINPUT75), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n418));
  INV_X1    g232(.A(G140), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(G125), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G146), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(G125), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n376), .A2(G140), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n226), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n275), .A2(G214), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n213), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n275), .A2(G143), .A3(G214), .ZN(new_n429));
  NAND2_X1  g243(.A1(KEYINPUT18), .A2(G131), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n197), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n432), .A2(KEYINPUT88), .A3(KEYINPUT18), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT88), .B1(new_n432), .B2(KEYINPUT18), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n426), .B(new_n431), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n429), .ZN(new_n436));
  AOI21_X1  g250(.A(G143), .B1(new_n275), .B2(G214), .ZN(new_n437));
  OAI21_X1  g251(.A(G131), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n428), .A2(new_n197), .A3(new_n429), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT17), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n432), .A2(KEYINPUT17), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT16), .B1(new_n419), .B2(G125), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n226), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT16), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n417), .B2(new_n420), .ZN(new_n447));
  OAI21_X1  g261(.A(G146), .B1(new_n447), .B2(new_n443), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n441), .A2(new_n442), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n435), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G113), .B(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(new_n342), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n435), .A2(new_n449), .A3(new_n454), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n310), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n456), .A2(KEYINPUT90), .A3(new_n310), .A4(new_n457), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(G475), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n450), .A2(new_n452), .ZN(new_n463));
  INV_X1    g277(.A(G475), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n438), .A2(new_n439), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n465), .A2(new_n448), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n423), .A2(new_n424), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(KEYINPUT19), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(KEYINPUT19), .B2(new_n421), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n226), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n452), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n435), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n463), .A2(new_n464), .A3(new_n310), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT20), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n450), .A2(new_n452), .B1(new_n471), .B2(new_n435), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT20), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n464), .A4(new_n310), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n462), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(G234), .A2(G237), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n480), .A2(G952), .A3(new_n383), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(G902), .A3(G953), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n482), .B(KEYINPUT93), .Z(new_n483));
  XOR2_X1   g297(.A(KEYINPUT21), .B(G898), .Z(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g301(.A1(KEYINPUT91), .A2(KEYINPUT13), .ZN(new_n488));
  NAND2_X1  g302(.A1(KEYINPUT91), .A2(KEYINPUT13), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(G128), .A3(new_n213), .ZN(new_n491));
  XNOR2_X1  g305(.A(G128), .B(G143), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n488), .A3(new_n489), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n493), .A3(G134), .ZN(new_n494));
  XOR2_X1   g308(.A(G116), .B(G122), .Z(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G107), .ZN(new_n496));
  XNOR2_X1  g310(.A(G116), .B(G122), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n345), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n262), .A2(new_n492), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n494), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n249), .A2(KEYINPUT14), .A3(G122), .ZN(new_n504));
  OAI211_X1 g318(.A(G107), .B(new_n504), .C1(new_n495), .C2(KEYINPUT14), .ZN(new_n505));
  INV_X1    g319(.A(new_n500), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n262), .A2(new_n492), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n505), .B(new_n498), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n494), .A2(new_n499), .A3(KEYINPUT92), .A4(new_n500), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n503), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT9), .B(G234), .Z(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G217), .A3(new_n383), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n512), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n503), .A2(new_n508), .A3(new_n509), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n310), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n516), .B(new_n310), .C1(KEYINPUT15), .C2(new_n518), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n487), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n416), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT22), .B(G137), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n383), .A2(G221), .A3(G234), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n251), .A2(new_n253), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(G128), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n250), .A2(G128), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n531), .B2(G128), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n532), .B1(new_n534), .B2(new_n530), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G110), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n445), .A2(new_n448), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT24), .B(G110), .Z(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n448), .A2(new_n425), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n534), .A2(new_n538), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT76), .B(G110), .Z(new_n543));
  OAI211_X1 g357(.A(new_n532), .B(new_n543), .C1(new_n534), .C2(new_n530), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n529), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n545), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n528), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n551));
  OR2_X1    g365(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n550), .A2(new_n310), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G217), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(G234), .B2(new_n310), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT74), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n546), .A2(new_n549), .A3(new_n310), .A4(new_n552), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n555), .A2(G902), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n550), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n511), .ZN(new_n564));
  OAI21_X1  g378(.A(G221), .B1(new_n564), .B2(G902), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n565), .B(KEYINPUT78), .Z(new_n566));
  XOR2_X1   g380(.A(new_n566), .B(KEYINPUT79), .Z(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n352), .A2(new_n234), .A3(new_n354), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n323), .B2(new_n400), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n215), .A2(new_n363), .A3(KEYINPUT10), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n224), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n215), .A2(new_n363), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n323), .A2(new_n400), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n224), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n224), .A2(KEYINPUT12), .A3(new_n577), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n574), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G110), .B(G140), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n383), .A2(G227), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n583), .B(new_n584), .Z(new_n585));
  NOR2_X1   g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n573), .A2(new_n224), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n585), .B1(new_n573), .B2(new_n224), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT80), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT80), .ZN(new_n592));
  OAI221_X1 g406(.A(new_n592), .B1(new_n589), .B2(new_n588), .C1(new_n582), .C2(new_n585), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n593), .A3(new_n310), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G469), .ZN(new_n595));
  INV_X1    g409(.A(new_n585), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n588), .B2(new_n574), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n580), .A2(new_n581), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(new_n589), .ZN(new_n599));
  INV_X1    g413(.A(G469), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(KEYINPUT81), .A3(new_n600), .A4(new_n310), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n589), .B1(new_n581), .B2(new_n580), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n266), .A2(new_n267), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n603), .A2(new_n571), .A3(new_n569), .A4(new_n572), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n585), .B1(new_n604), .B2(new_n587), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n600), .B(new_n310), .C1(new_n602), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT81), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n568), .B1(new_n595), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n339), .A2(new_n525), .A3(new_n563), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  OAI21_X1  g426(.A(G472), .B1(new_n298), .B2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n286), .A2(new_n288), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT28), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n294), .B1(new_n326), .B2(new_n291), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n328), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n280), .B1(new_n617), .B2(new_n295), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n300), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n613), .A2(new_n620), .A3(new_n563), .A4(new_n610), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n486), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n411), .B1(new_n387), .B2(new_n409), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n414), .B1(new_n623), .B2(KEYINPUT94), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n387), .A2(new_n409), .A3(new_n625), .A4(new_n411), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n341), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n516), .A2(KEYINPUT33), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n513), .A2(new_n629), .A3(new_n515), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(G478), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(G478), .A2(G902), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n516), .A2(new_n518), .A3(new_n310), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n479), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n627), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n622), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n474), .A2(new_n641), .A3(new_n477), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n473), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(new_n462), .A3(new_n522), .A4(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n622), .A2(new_n627), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n613), .A2(new_n620), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n547), .A2(new_n548), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n529), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n560), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n559), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n610), .A2(new_n654), .ZN(new_n655));
  NOR4_X1   g469(.A1(new_n649), .A2(new_n655), .A3(new_n416), .A4(new_n524), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT37), .B(G110), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  AND2_X1   g472(.A1(new_n610), .A2(new_n654), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n481), .B1(new_n483), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT96), .B1(new_n645), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT96), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n644), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n339), .A2(new_n659), .A3(new_n627), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XNOR2_X1  g482(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n661), .B(new_n669), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n610), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT40), .Z(new_n672));
  INV_X1    g486(.A(new_n341), .ZN(new_n673));
  INV_X1    g487(.A(new_n654), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n413), .A2(new_n414), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n672), .A2(new_n673), .A3(new_n674), .A4(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n479), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n523), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n303), .A2(new_n280), .A3(new_n305), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n284), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n301), .A2(new_n338), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n679), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  NAND2_X1  g501(.A1(new_n624), .A2(new_n626), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n479), .A2(new_n634), .A3(new_n662), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n673), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT99), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n627), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n339), .A2(new_n691), .A3(new_n659), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  OAI21_X1  g509(.A(new_n310), .B1(new_n602), .B2(new_n605), .ZN(new_n696));
  AOI221_X4 g510(.A(new_n566), .B1(G469), .B2(new_n696), .C1(new_n601), .C2(new_n608), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n486), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n339), .A2(new_n637), .A3(new_n563), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NOR3_X1   g516(.A1(new_n698), .A2(new_n486), .A3(new_n562), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n339), .A3(new_n627), .A4(new_n645), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NAND3_X1  g519(.A1(new_n688), .A2(new_n697), .A3(new_n673), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n627), .A2(KEYINPUT100), .A3(new_n697), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n524), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n339), .A4(new_n654), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  INV_X1    g527(.A(G472), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n337), .B2(new_n310), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n306), .A2(new_n296), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n280), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n300), .B1(new_n614), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n688), .A2(new_n673), .A3(new_n681), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n699), .A3(new_n720), .A4(new_n563), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR3_X1   g536(.A1(new_n715), .A2(new_n674), .A3(new_n718), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n708), .A3(new_n689), .A4(new_n709), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  NOR2_X1   g539(.A1(new_n675), .A2(new_n341), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n310), .B1(new_n586), .B2(new_n590), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n566), .B1(new_n609), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n339), .A2(new_n563), .A3(new_n689), .A4(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT101), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n338), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n619), .A2(KEYINPUT101), .A3(KEYINPUT32), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n332), .A4(new_n301), .ZN(new_n737));
  AND4_X1   g551(.A1(KEYINPUT42), .A2(new_n726), .A3(new_n729), .A4(new_n689), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n563), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT102), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT102), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n733), .A2(new_n742), .A3(new_n739), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NAND4_X1  g559(.A1(new_n339), .A2(new_n563), .A3(new_n666), .A4(new_n730), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  NAND2_X1  g561(.A1(new_n680), .A2(new_n634), .ZN(new_n748));
  XOR2_X1   g562(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT106), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n748), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n649), .A3(new_n654), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT107), .Z(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n591), .A2(new_n758), .A3(new_n593), .ZN(new_n759));
  OR3_X1    g573(.A1(new_n586), .A2(new_n758), .A3(new_n590), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT103), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n609), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n765), .A2(KEYINPUT103), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n566), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n670), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT104), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n754), .A2(new_n755), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n757), .A2(new_n726), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G137), .ZN(G39));
  XNOR2_X1  g592(.A(new_n771), .B(KEYINPUT47), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n339), .A2(new_n563), .A3(new_n635), .A4(new_n661), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n726), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NAND2_X1  g596(.A1(new_n567), .A2(new_n673), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n696), .A2(G469), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n609), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n680), .B(new_n634), .C1(new_n786), .C2(KEYINPUT49), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n783), .B(new_n787), .C1(KEYINPUT49), .C2(new_n786), .ZN(new_n788));
  INV_X1    g602(.A(new_n685), .ZN(new_n789));
  INV_X1    g603(.A(new_n677), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n788), .A2(new_n563), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n723), .A2(new_n689), .A3(new_n730), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n339), .A2(new_n659), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n523), .A2(new_n462), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n413), .A3(new_n673), .A4(new_n414), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n642), .A2(new_n643), .A3(new_n662), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n797), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n726), .A2(KEYINPUT110), .A3(new_n799), .A4(new_n795), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n793), .A2(KEYINPUT111), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT111), .B1(new_n793), .B2(new_n801), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n746), .B(new_n792), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n621), .A2(new_n416), .A3(new_n486), .A4(new_n635), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n656), .ZN(new_n806));
  INV_X1    g620(.A(new_n621), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n415), .A2(new_n522), .ZN(new_n808));
  INV_X1    g622(.A(new_n487), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT109), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n808), .A2(KEYINPUT109), .A3(new_n809), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n806), .A2(new_n611), .A3(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n712), .A2(new_n700), .A3(new_n704), .A4(new_n721), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n804), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n724), .A2(new_n694), .A3(new_n667), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n684), .B1(new_n619), .B2(KEYINPUT32), .ZN(new_n817));
  INV_X1    g631(.A(new_n338), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n720), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n654), .A2(new_n661), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n729), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n729), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT113), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n824), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n823), .B1(new_n729), .B2(new_n820), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n685), .A4(new_n720), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(new_n816), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n816), .A2(new_n832), .A3(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n733), .B2(new_n739), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n815), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n816), .A2(KEYINPUT52), .A3(new_n832), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n744), .B1(new_n840), .B2(new_n833), .ZN(new_n841));
  INV_X1    g655(.A(new_n814), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n812), .A2(new_n611), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n843), .A2(new_n656), .A3(new_n805), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n746), .A2(new_n792), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n793), .A2(new_n801), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT111), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n793), .A2(KEYINPUT111), .A3(new_n801), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n837), .B1(new_n841), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(KEYINPUT116), .B(new_n837), .C1(new_n841), .C2(new_n851), .ZN(new_n855));
  AOI211_X1 g669(.A(KEYINPUT54), .B(new_n839), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n841), .A2(new_n851), .A3(new_n837), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT115), .Z(new_n859));
  XOR2_X1   g673(.A(new_n852), .B(KEYINPUT114), .Z(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n857), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g677(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n864));
  NAND4_X1  g678(.A1(new_n753), .A2(new_n481), .A3(new_n563), .A4(new_n719), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n341), .A3(new_n790), .A4(new_n697), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT50), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT118), .Z(new_n869));
  NOR2_X1   g683(.A1(new_n786), .A2(new_n567), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n726), .B(new_n866), .C1(new_n779), .C2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n726), .A2(new_n481), .A3(new_n697), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n753), .A2(new_n723), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n789), .A2(new_n872), .A3(new_n563), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n479), .A2(new_n634), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n871), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n864), .B1(new_n869), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n877), .A2(new_n879), .A3(new_n868), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n737), .A2(new_n563), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n753), .A3(new_n872), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT48), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n874), .A2(new_n636), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(G952), .A3(new_n383), .A4(new_n886), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n884), .B(new_n887), .C1(new_n710), .C2(new_n866), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n878), .A2(new_n880), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n863), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n791), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NAND2_X1  g706(.A1(new_n854), .A2(new_n855), .ZN(new_n893));
  INV_X1    g707(.A(new_n839), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n310), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G210), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n375), .B(new_n386), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n896), .B2(new_n897), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n383), .A2(G952), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G51));
  XOR2_X1   g717(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(G469), .A3(G902), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n862), .B1(new_n893), .B2(new_n894), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(new_n856), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n904), .B1(G469), .B2(G902), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n599), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n895), .A2(G469), .A3(new_n760), .A4(new_n759), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(new_n475), .Z(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n902), .ZN(G60));
  NAND2_X1  g728(.A1(new_n628), .A2(new_n630), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT120), .Z(new_n916));
  XNOR2_X1  g730(.A(new_n632), .B(KEYINPUT59), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n863), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n906), .B2(new_n856), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n921));
  INV_X1    g735(.A(new_n902), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n923), .B(new_n919), .C1(new_n906), .C2(new_n856), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n921), .A2(KEYINPUT122), .A3(new_n922), .A4(new_n924), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n918), .B1(new_n927), .B2(new_n928), .ZN(G63));
  XNOR2_X1  g743(.A(new_n550), .B(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n893), .A2(new_n894), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  AOI21_X1  g747(.A(new_n930), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n902), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n931), .A2(new_n933), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n652), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n937), .A3(KEYINPUT61), .ZN(new_n938));
  OAI211_X1 g752(.A(KEYINPUT125), .B(new_n922), .C1(new_n936), .C2(new_n930), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n934), .B2(new_n902), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n939), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g756(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(G66));
  AOI21_X1  g758(.A(new_n383), .B1(new_n484), .B2(G224), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n813), .A2(new_n814), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n947), .B2(new_n383), .ZN(new_n948));
  INV_X1    g762(.A(new_n375), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(G898), .B2(new_n383), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n948), .B(new_n950), .Z(G69));
  NAND3_X1  g765(.A1(new_n777), .A2(new_n744), .A3(new_n781), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n773), .A2(new_n720), .A3(new_n881), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n746), .A3(new_n816), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n383), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n242), .B(new_n469), .Z(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n955), .B(new_n957), .C1(G900), .C2(new_n383), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n686), .A2(new_n816), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  NOR3_X1   g774(.A1(new_n671), .A2(new_n341), .A3(new_n675), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n635), .B1(new_n523), .B2(new_n479), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n339), .A3(new_n563), .A4(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n960), .A2(new_n777), .A3(new_n781), .A4(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n383), .A3(new_n956), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n383), .B1(G227), .B2(G900), .ZN(new_n966));
  AOI22_X1  g780(.A1(new_n958), .A2(new_n965), .B1(KEYINPUT127), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n964), .B2(new_n947), .ZN(new_n972));
  INV_X1    g786(.A(new_n316), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n277), .A3(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n952), .A2(new_n954), .A3(new_n947), .ZN(new_n975));
  INV_X1    g789(.A(new_n971), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n280), .B(new_n316), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n922), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n973), .A2(new_n280), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n861), .B1(new_n284), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n971), .B2(new_n980), .ZN(G57));
endmodule


