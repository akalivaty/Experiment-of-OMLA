//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT86), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G952), .ZN(new_n190));
  AOI211_X1 g004(.A(G953), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT21), .B(G898), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G902), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  AOI211_X1 g009(.A(new_n194), .B(new_n195), .C1(G234), .C2(G237), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n191), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT81), .B1(new_n199), .B2(G104), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT81), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G107), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n199), .A3(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n200), .A2(new_n203), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n210), .A2(new_n211), .A3(new_n205), .A4(new_n207), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n214), .B(G101), .C1(new_n204), .C2(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G116), .B(G119), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT72), .B1(new_n217), .B2(KEYINPUT71), .ZN(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G116), .ZN(new_n220));
  INV_X1    g034(.A(G116), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G119), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT72), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT2), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT70), .B1(KEYINPUT2), .B2(G113), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n230), .A2(new_n231), .B1(KEYINPUT2), .B2(G113), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n218), .A2(new_n226), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n218), .B2(new_n226), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT87), .B1(new_n216), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n220), .A2(KEYINPUT5), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(new_n229), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n238), .A2(new_n239), .B1(new_n232), .B2(new_n217), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n202), .A2(G107), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n199), .A2(G104), .ZN(new_n242));
  OAI21_X1  g056(.A(G101), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n212), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT83), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n212), .B2(new_n243), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n240), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n218), .A2(new_n226), .ZN(new_n249));
  INV_X1    g063(.A(new_n232), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n218), .A2(new_n226), .A3(new_n232), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT87), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n215), .A4(new_n213), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n236), .A2(new_n248), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G110), .B(G122), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n236), .A2(new_n257), .A3(new_n255), .A4(new_n248), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(KEYINPUT6), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT88), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT88), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n259), .A2(new_n263), .A3(KEYINPUT6), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT0), .ZN(new_n275));
  INV_X1    g089(.A(G128), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G125), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n276), .A2(KEYINPUT1), .ZN(new_n280));
  INV_X1    g094(.A(G146), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G143), .ZN(new_n282));
  INV_X1    g096(.A(G143), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G146), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n272), .A2(KEYINPUT68), .A3(new_n280), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT1), .B1(new_n283), .B2(G146), .ZN(new_n290));
  OR2_X1    g104(.A1(KEYINPUT69), .A2(G128), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT69), .A2(G128), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n273), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G125), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n279), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT90), .B(G224), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n195), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n298), .B(new_n300), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT89), .B1(new_n259), .B2(KEYINPUT6), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT89), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT6), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n256), .A2(new_n304), .A3(new_n305), .A4(new_n258), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n265), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n298), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n300), .A2(KEYINPUT7), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n257), .B(KEYINPUT8), .Z(new_n312));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n238), .B1(new_n239), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT91), .B1(new_n217), .B2(KEYINPUT5), .ZN(new_n315));
  OAI22_X1  g129(.A1(new_n314), .A2(new_n315), .B1(new_n250), .B2(new_n223), .ZN(new_n316));
  INV_X1    g130(.A(new_n244), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n240), .A2(new_n244), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n310), .A2(new_n311), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n298), .A2(KEYINPUT7), .A3(new_n300), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n260), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n194), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT92), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n308), .A2(new_n309), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n309), .B1(new_n308), .B2(new_n324), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n189), .B(new_n198), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(G475), .A2(G902), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT16), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n296), .A2(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n331), .B1(new_n334), .B2(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n281), .ZN(new_n336));
  OAI211_X1 g150(.A(G146), .B(new_n331), .C1(new_n334), .C2(new_n329), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G237), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n195), .A3(G214), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT93), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n283), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n283), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT93), .A2(G143), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n342), .B1(new_n345), .B2(new_n340), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT66), .B(G131), .Z(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT95), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT17), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT95), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n352), .A3(new_n347), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n349), .A2(new_n350), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n349), .A2(new_n353), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n338), .B(new_n354), .C1(new_n355), .C2(new_n351), .ZN(new_n356));
  XNOR2_X1  g170(.A(G113), .B(G122), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(new_n202), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT94), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT18), .ZN(new_n360));
  INV_X1    g174(.A(G131), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n346), .A2(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n334), .A2(G146), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n332), .A2(new_n333), .A3(new_n281), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n356), .A2(new_n358), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n349), .A2(new_n353), .A3(new_n350), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n334), .B(KEYINPUT19), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n371), .B(new_n337), .C1(G146), .C2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n358), .B1(new_n373), .B2(new_n369), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n370), .A2(KEYINPUT96), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n369), .ZN(new_n377));
  INV_X1    g191(.A(new_n358), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n356), .A2(new_n358), .A3(new_n369), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT20), .B(new_n328), .C1(new_n375), .C2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n358), .B1(new_n356), .B2(new_n369), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n194), .B1(new_n370), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G475), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n328), .B1(new_n370), .B2(new_n374), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT20), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G116), .B(G122), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n199), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n221), .A2(KEYINPUT14), .A3(G122), .ZN(new_n392));
  INV_X1    g206(.A(new_n390), .ZN(new_n393));
  OAI211_X1 g207(.A(G107), .B(new_n392), .C1(new_n393), .C2(KEYINPUT14), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT69), .B(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G143), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n283), .A2(G128), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G134), .ZN(new_n399));
  INV_X1    g213(.A(G134), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n396), .B2(new_n397), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n391), .B(new_n394), .C1(new_n399), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT13), .B1(new_n395), .B2(G143), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n398), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n396), .A2(KEYINPUT13), .A3(G134), .A4(new_n397), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n390), .B(new_n199), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT97), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(KEYINPUT97), .A3(new_n408), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n403), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT9), .B(G234), .Z(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n415), .A2(new_n416), .A3(G953), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n417), .ZN(new_n419));
  AOI211_X1 g233(.A(new_n419), .B(new_n403), .C1(new_n411), .C2(new_n412), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n194), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n421), .B(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n389), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n327), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n290), .A2(G128), .B1(new_n282), .B2(new_n284), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n287), .B2(new_n288), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n244), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT82), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n433), .B(new_n428), .C1(new_n244), .C2(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT11), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n400), .B2(G137), .ZN(new_n437));
  INV_X1    g251(.A(G137), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT11), .A3(G134), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n400), .A2(G137), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G131), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n441), .A2(new_n347), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(KEYINPUT67), .A3(G131), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n213), .A2(new_n278), .A3(new_n215), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT10), .B(new_n295), .C1(new_n245), .C2(new_n247), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n435), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G140), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n195), .A2(G227), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n452), .B(new_n453), .Z(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n317), .A2(new_n295), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n244), .A2(new_n430), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n447), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n460), .B(KEYINPUT12), .Z(new_n461));
  NAND3_X1  g275(.A1(new_n451), .A2(KEYINPUT84), .A3(new_n454), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n435), .A2(new_n449), .A3(new_n450), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n447), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n451), .ZN(new_n468));
  INV_X1    g282(.A(new_n454), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n457), .A2(KEYINPUT85), .A3(new_n461), .A4(new_n462), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n194), .ZN(new_n474));
  NAND2_X1  g288(.A1(G469), .A2(G902), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n461), .A2(new_n451), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n469), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(new_n451), .A3(new_n454), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(G469), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G221), .B1(new_n415), .B2(G902), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n416), .B1(G234), .B2(new_n194), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT23), .B1(new_n276), .B2(G119), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT76), .B1(new_n219), .B2(G128), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT76), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n276), .A3(G119), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n292), .ZN(new_n489));
  NOR2_X1   g303(.A1(KEYINPUT69), .A2(G128), .ZN(new_n490));
  OAI211_X1 g304(.A(KEYINPUT23), .B(G119), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT77), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n488), .A2(new_n491), .A3(KEYINPUT77), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(G110), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT78), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n395), .A2(G119), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n276), .A2(G119), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n219), .B1(new_n291), .B2(new_n292), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT75), .B1(new_n504), .B2(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT24), .B(G110), .Z(new_n507));
  AOI22_X1  g321(.A1(new_n506), .A2(new_n507), .B1(new_n337), .B2(new_n336), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT78), .A4(G110), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n498), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n506), .A2(new_n507), .B1(G110), .B2(new_n492), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n337), .A3(new_n367), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT80), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT80), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n510), .A2(new_n515), .A3(new_n512), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT79), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n514), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(KEYINPUT80), .A3(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT25), .B1(new_n524), .B2(new_n194), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n526));
  AOI211_X1 g340(.A(new_n526), .B(G902), .C1(new_n522), .C2(new_n523), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n483), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n483), .A2(G902), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(G472), .A2(G902), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n274), .A2(KEYINPUT65), .A3(new_n277), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT65), .ZN(new_n534));
  INV_X1    g348(.A(new_n277), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n272), .B1(new_n269), .B2(new_n270), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n447), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n441), .A2(new_n347), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n289), .B2(new_n294), .ZN(new_n540));
  INV_X1    g354(.A(new_n440), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n400), .A2(G137), .ZN(new_n542));
  OAI21_X1  g356(.A(G131), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n278), .A2(new_n447), .B1(new_n540), .B2(new_n543), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT30), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n253), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n235), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n339), .A2(new_n195), .A3(G210), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT74), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT26), .B(G101), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n550), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n558), .A2(KEYINPUT31), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT31), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n550), .A2(new_n560), .A3(new_n551), .A4(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n545), .A2(new_n253), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT28), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n548), .B2(new_n235), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n447), .A2(new_n278), .ZN(new_n565));
  AND4_X1   g379(.A1(new_n563), .A2(new_n565), .A3(new_n544), .A4(new_n235), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n562), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n557), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n532), .B1(new_n559), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT32), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n558), .A2(KEYINPUT31), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n561), .A3(new_n569), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n532), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(new_n557), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n550), .A2(new_n551), .A3(new_n568), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT29), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n548), .A2(new_n235), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n564), .B2(new_n566), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n557), .A2(KEYINPUT29), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n194), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G472), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n573), .A2(new_n576), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n531), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n427), .A2(new_n482), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  OR2_X1    g403(.A1(new_n413), .A2(new_n417), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n413), .A2(new_n417), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(KEYINPUT33), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n418), .B2(new_n420), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n422), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n421), .A2(G478), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n422), .A2(new_n194), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n389), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT98), .B1(new_n327), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n309), .ZN(new_n601));
  AOI221_X4 g415(.A(new_n301), .B1(new_n303), .B2(new_n306), .C1(new_n262), .C2(new_n264), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n323), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n601), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n308), .A2(new_n309), .A3(new_n324), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n188), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n598), .A2(new_n389), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n607), .A2(new_n608), .A3(new_n198), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n528), .A2(new_n530), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n561), .A2(new_n569), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n613), .B2(new_n574), .ZN(new_n614));
  INV_X1    g428(.A(G472), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n571), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n480), .A2(new_n617), .A3(new_n481), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NAND3_X1  g435(.A1(new_n480), .A2(new_n617), .A3(new_n481), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n375), .A2(new_n381), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n328), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n387), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n382), .A2(new_n385), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n424), .A3(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n622), .A2(new_n327), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G107), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NAND2_X1  g444(.A1(new_n605), .A2(new_n606), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(new_n189), .A3(new_n198), .A4(new_n425), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n616), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n480), .A2(new_n481), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n635));
  INV_X1    g449(.A(new_n483), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n516), .A2(new_n521), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n515), .B1(new_n510), .B2(new_n512), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n523), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n194), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n526), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n524), .A2(KEYINPUT25), .A3(new_n194), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n636), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n513), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n529), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n635), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n528), .A2(KEYINPUT99), .A3(new_n647), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n634), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n633), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(G12));
  OAI211_X1 g470(.A(new_n585), .B(new_n189), .C1(new_n325), .C2(new_n326), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n651), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n196), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n191), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n627), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n482), .A2(new_n658), .A3(new_n659), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT101), .B(G128), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G30));
  XNOR2_X1  g482(.A(new_n663), .B(KEYINPUT39), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n482), .A2(new_n669), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n188), .B(new_n659), .C1(new_n670), .C2(KEYINPUT40), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n573), .A2(new_n576), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n550), .A2(new_n551), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n568), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n568), .A2(new_n551), .A3(new_n580), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n194), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n389), .A2(new_n424), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n670), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n631), .B(new_n685), .Z(new_n686));
  AND3_X1   g500(.A1(new_n671), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT103), .B(G143), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G45));
  NOR2_X1   g503(.A1(new_n599), .A2(new_n664), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n482), .A2(new_n658), .A3(new_n659), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n472), .A2(new_n194), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G469), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n481), .A3(new_n474), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n586), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n611), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n693), .B1(new_n611), .B2(new_n697), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT41), .B(G113), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n695), .A2(new_n198), .A3(new_n481), .A4(new_n474), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n531), .A2(new_n424), .A3(new_n626), .A4(new_n625), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n703), .A2(new_n704), .A3(new_n657), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT105), .B(G116), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G18));
  NOR4_X1   g521(.A1(new_n703), .A2(new_n657), .A3(new_n651), .A4(new_n426), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT106), .B(G119), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G21));
  OAI21_X1  g524(.A(new_n189), .B1(new_n325), .B2(new_n326), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n575), .A2(new_n194), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n532), .B(KEYINPUT107), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n581), .A2(new_n568), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n574), .A2(new_n561), .A3(new_n714), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n712), .A2(G472), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n528), .A3(new_n530), .A4(new_n198), .ZN(new_n717));
  NOR4_X1   g531(.A1(new_n696), .A2(new_n711), .A3(new_n717), .A4(new_n679), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(G122), .Z(G24));
  INV_X1    g533(.A(new_n716), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n651), .A2(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n695), .A2(new_n481), .A3(new_n474), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n722), .A3(new_n607), .A4(new_n690), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n478), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(G469), .A3(new_n477), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n474), .A2(new_n475), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n474), .A2(KEYINPUT109), .A3(new_n475), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n605), .A2(new_n189), .A3(new_n606), .A4(new_n481), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT110), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n587), .A4(new_n690), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n737), .B1(new_n732), .B2(new_n734), .ZN(new_n741));
  AOI211_X1 g555(.A(KEYINPUT110), .B(new_n733), .C1(new_n730), .C2(new_n731), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n587), .B(new_n690), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  OAI211_X1 g561(.A(new_n587), .B(new_n665), .C1(new_n741), .C2(new_n742), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n479), .B1(new_n750), .B2(new_n473), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n726), .A2(KEYINPUT45), .A3(new_n477), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n479), .B(KEYINPUT111), .C1(new_n750), .C2(new_n473), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n475), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n474), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT46), .B1(new_n756), .B2(new_n475), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n481), .B(new_n669), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n595), .ZN(new_n762));
  INV_X1    g576(.A(new_n596), .ZN(new_n763));
  INV_X1    g577(.A(new_n597), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n389), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n765), .B2(new_n389), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n616), .A3(new_n659), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n631), .A2(new_n188), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n761), .A2(new_n773), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  OAI21_X1  g591(.A(new_n481), .B1(new_n758), .B2(new_n759), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n531), .A2(new_n585), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n774), .A2(new_n690), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n782), .B(new_n481), .C1(new_n758), .C2(new_n759), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n666), .A2(new_n691), .A3(new_n723), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n711), .B1(new_n730), .B2(new_n731), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n678), .A2(new_n481), .A3(new_n680), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n644), .A2(new_n648), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n663), .B(KEYINPUT115), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n786), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n652), .B(new_n658), .C1(new_n665), .C2(new_n690), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n786), .A2(new_n792), .A3(new_n794), .A4(new_n723), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n708), .A2(new_n718), .A3(new_n705), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n698), .B2(new_n699), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n626), .A2(new_n424), .A3(new_n388), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n622), .A2(new_n327), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n652), .B2(new_n633), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n632), .A2(new_n634), .A3(new_n586), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n631), .A2(new_n189), .A3(new_n198), .A4(new_n609), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n622), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT113), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n327), .A2(new_n599), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n618), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n588), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n801), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n690), .B(new_n721), .C1(new_n741), .C2(new_n742), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n625), .A2(new_n626), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n424), .A2(new_n664), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n774), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n774), .A2(KEYINPUT114), .A3(new_n813), .A4(new_n814), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n585), .A3(new_n652), .A4(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n748), .A2(new_n812), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n796), .A2(new_n811), .A3(new_n746), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n748), .A2(new_n812), .A3(new_n819), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n798), .A3(new_n810), .ZN(new_n825));
  INV_X1    g639(.A(new_n792), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n666), .A2(new_n691), .A3(new_n723), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT116), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .ZN(new_n829));
  OAI211_X1 g643(.A(KEYINPUT116), .B(new_n786), .C1(new_n826), .C2(new_n827), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n825), .A2(new_n831), .A3(KEYINPUT53), .A4(new_n746), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n825), .A2(new_n746), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n822), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT117), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n821), .A2(new_n822), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n835), .A2(new_n839), .A3(new_n822), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n834), .B1(new_n841), .B2(KEYINPUT54), .ZN(new_n842));
  INV_X1    g656(.A(new_n770), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n531), .A2(new_n191), .A3(new_n716), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n188), .ZN(new_n846));
  INV_X1    g660(.A(new_n686), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n722), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT50), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n846), .B2(new_n848), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n722), .A2(new_n191), .A3(new_n774), .ZN(new_n853));
  INV_X1    g667(.A(new_n678), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n531), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n598), .A2(new_n389), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n850), .A2(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n843), .A2(new_n853), .ZN(new_n859));
  INV_X1    g673(.A(new_n721), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n845), .A2(new_n774), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT118), .Z(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n779), .A2(new_n783), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n695), .A2(new_n474), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n866), .A2(KEYINPUT119), .B1(new_n481), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n866), .A2(KEYINPUT119), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n858), .A2(new_n861), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n867), .A2(new_n481), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n779), .B2(new_n783), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n864), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(G952), .B(new_n195), .C1(new_n872), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n859), .A2(new_n586), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT48), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n853), .A2(new_n599), .A3(new_n855), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n871), .A2(new_n876), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n845), .A2(new_n607), .A3(new_n722), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n842), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(G952), .B2(G953), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n531), .A2(new_n189), .A3(new_n481), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT112), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(new_n766), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n867), .B(KEYINPUT49), .Z(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n847), .A3(new_n854), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n883), .A2(new_n888), .ZN(G75));
  AOI21_X1  g703(.A(new_n194), .B1(new_n823), .B2(new_n832), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT56), .B1(new_n890), .B2(G210), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n265), .A2(new_n307), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n302), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n891), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n195), .A2(G952), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(G51));
  XNOR2_X1  g711(.A(new_n833), .B(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n475), .A2(KEYINPUT57), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n475), .A2(KEYINPUT57), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n472), .ZN(new_n902));
  INV_X1    g716(.A(new_n756), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n890), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n896), .B1(new_n902), .B2(new_n904), .ZN(G54));
  NAND2_X1  g719(.A1(KEYINPUT58), .A2(G475), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT120), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n890), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(new_n623), .Z(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n896), .ZN(G60));
  NAND2_X1  g724(.A1(new_n592), .A2(new_n594), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n597), .B(KEYINPUT59), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n842), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n896), .ZN(new_n914));
  INV_X1    g728(.A(new_n912), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n898), .A2(new_n594), .A3(new_n592), .A4(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT121), .Z(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT60), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n833), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT122), .ZN(new_n922));
  INV_X1    g736(.A(new_n524), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n833), .A2(new_n924), .A3(new_n920), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n833), .B2(new_n920), .ZN(new_n927));
  INV_X1    g741(.A(new_n920), .ZN(new_n928));
  AOI211_X1 g742(.A(KEYINPUT122), .B(new_n928), .C1(new_n823), .C2(new_n832), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n646), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n896), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n926), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n931), .A2(new_n932), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n935), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n926), .A2(new_n930), .A3(new_n937), .A4(new_n933), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(G66));
  NOR2_X1   g753(.A1(new_n811), .A2(G953), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n195), .B1(new_n192), .B2(new_n299), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT124), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(KEYINPUT124), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n892), .B1(G898), .B2(new_n195), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  AOI21_X1  g759(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n547), .A2(new_n549), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n372), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(G900), .A2(G953), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n746), .A2(new_n776), .A3(new_n784), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n760), .A2(new_n586), .A3(new_n711), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n827), .B1(new_n952), .B2(new_n680), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n951), .A2(KEYINPUT126), .A3(new_n748), .A4(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n776), .A2(new_n784), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(new_n746), .A3(new_n748), .A4(new_n953), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n949), .B(new_n950), .C1(new_n959), .C2(G953), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n946), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n687), .A2(new_n827), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n586), .B1(new_n599), .B2(new_n799), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n682), .A2(new_n774), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n955), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(new_n195), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n960), .B1(new_n968), .B2(new_n949), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n962), .B(new_n969), .Z(G72));
  XOR2_X1   g784(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n971));
  NOR2_X1   g785(.A1(new_n615), .A2(new_n194), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n811), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n959), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n673), .A3(new_n568), .ZN(new_n976));
  INV_X1    g790(.A(new_n674), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n841), .A2(new_n578), .A3(new_n977), .A4(new_n973), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n973), .B1(new_n967), .B2(new_n974), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n674), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n914), .A2(new_n976), .A3(new_n978), .A4(new_n980), .ZN(G57));
endmodule


