//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n439), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(G567), .A2(new_n455), .B1(new_n453), .B2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT3), .B1(new_n461), .B2(KEYINPUT68), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n460), .A3(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n470), .B1(new_n478), .B2(new_n468), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(new_n468), .B2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n476), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OR3_X1    g059(.A1(new_n483), .A2(KEYINPUT69), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n476), .A2(new_n468), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n485), .A2(new_n486), .B1(G124), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND3_X1  g067(.A1(new_n473), .A2(new_n475), .A3(G126), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n468), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n461), .A2(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n496), .A2(G102), .ZN(new_n497));
  OR3_X1    g072(.A1(new_n495), .A2(KEYINPUT70), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n468), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n502), .B1(new_n462), .B2(new_n463), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT4), .A2(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n507));
  OAI211_X1 g082(.A(G138), .B(new_n504), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n500), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT70), .B1(new_n495), .B2(new_n497), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n498), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(G543), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n518), .A2(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT72), .Z(new_n528));
  OAI21_X1  g103(.A(G651), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n520), .B2(new_n534), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT73), .Z(new_n536));
  NAND3_X1  g111(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n537));
  INV_X1    g112(.A(new_n523), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  AOI22_X1  g116(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n520), .A2(new_n545), .B1(new_n546), .B2(new_n523), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n543), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n520), .A2(new_n551), .B1(new_n552), .B2(new_n523), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  AOI22_X1  g136(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT75), .Z(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  XNOR2_X1  g139(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n523), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n538), .A2(new_n568), .A3(KEYINPUT9), .A4(G53), .ZN(new_n569));
  INV_X1    g144(.A(new_n520), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G91), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n564), .A2(new_n567), .A3(new_n569), .A4(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  NAND2_X1  g148(.A1(new_n570), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n538), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n515), .A2(new_n517), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT76), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n538), .A2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n570), .A2(G86), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n538), .A2(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n588), .B2(new_n520), .C1(new_n543), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n518), .A2(G92), .A3(new_n519), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT77), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(KEYINPUT10), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n593), .A2(KEYINPUT10), .B1(G54), .B2(new_n538), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n518), .A2(G66), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n543), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n554), .A2(new_n604), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n600), .A2(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n464), .A2(new_n496), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT13), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n487), .A2(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n482), .A2(G135), .ZN(new_n619));
  NOR2_X1   g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT78), .Z(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT15), .B(G2435), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2443), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n642), .A2(new_n643), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(KEYINPUT17), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(new_n644), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n645), .B(KEYINPUT80), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n647), .B(new_n651), .C1(new_n649), .C2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT81), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n659), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT82), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n667), .B2(KEYINPUT20), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n668), .B(new_n669), .C1(KEYINPUT20), .C2(new_n667), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1986), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1981), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1991), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT33), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1976), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n677), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(G1971), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(G1971), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n677), .A2(G6), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G305), .B2(G16), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT32), .B(G1981), .Z(new_n689));
  AOI211_X1 g264(.A(new_n685), .B(new_n686), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n682), .B(new_n690), .C1(new_n688), .C2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT84), .B(KEYINPUT34), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n487), .A2(G119), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n482), .A2(G131), .ZN(new_n697));
  NOR2_X1   g272(.A1(G95), .A2(G2105), .ZN(new_n698));
  OAI21_X1  g273(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT83), .Z(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n692), .A2(new_n694), .ZN(new_n705));
  MUX2_X1   g280(.A(G24), .B(G290), .S(G16), .Z(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(G1986), .Z(new_n707));
  NAND4_X1  g282(.A1(new_n695), .A2(new_n704), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT36), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT28), .ZN(new_n710));
  INV_X1    g285(.A(G26), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n482), .A2(G140), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT86), .ZN(new_n715));
  OR2_X1    g290(.A1(G104), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT87), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n487), .A2(G128), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n715), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n713), .B1(new_n720), .B2(G29), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n712), .B1(new_n721), .B2(new_n710), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(G2067), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G21), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G168), .B2(G16), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(G1966), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT93), .Z(new_n727));
  NOR2_X1   g302(.A1(G5), .A2(G16), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G171), .B2(G16), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n725), .A2(G1966), .B1(G1961), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G34), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT24), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT24), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n471), .A2(new_n480), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2084), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n727), .A2(new_n730), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G29), .A2(G32), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n487), .A2(G129), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n482), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n496), .A2(G105), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n743), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n740), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n729), .A2(G1961), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n622), .A2(KEYINPUT92), .A3(new_n734), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT30), .B(G28), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n734), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  OAI21_X1  g331(.A(KEYINPUT92), .B1(new_n622), .B2(new_n734), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n752), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n601), .A2(new_n677), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G4), .B2(new_n677), .ZN(new_n760));
  INV_X1    g335(.A(G1348), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n739), .A2(new_n751), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n677), .A2(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n555), .B2(new_n677), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G1341), .Z(new_n767));
  NOR2_X1   g342(.A1(G164), .A2(new_n734), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G27), .B2(new_n734), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT23), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n677), .A2(G20), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n772), .B(new_n773), .C1(G299), .C2(G16), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT94), .B(G1956), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n734), .A2(G35), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G162), .B2(new_n734), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT29), .B(G2090), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n779), .B(new_n780), .Z(new_n781));
  AOI22_X1  g356(.A1(G2067), .A2(new_n722), .B1(new_n769), .B2(new_n770), .ZN(new_n782));
  AND4_X1   g357(.A1(new_n771), .A2(new_n777), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n734), .A2(G33), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n496), .A2(G103), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT88), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT25), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n482), .A2(G139), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n787), .B(new_n788), .C1(new_n468), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT89), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n784), .B1(new_n791), .B2(new_n734), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT90), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2072), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n764), .A2(new_n767), .A3(new_n783), .A4(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n709), .A2(new_n723), .A3(new_n796), .ZN(G311));
  NAND3_X1  g372(.A1(new_n709), .A2(new_n723), .A3(new_n796), .ZN(G150));
  NAND2_X1  g373(.A1(G80), .A2(G543), .ZN(new_n799));
  INV_X1    g374(.A(G67), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n579), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(new_n543), .ZN(new_n804));
  INV_X1    g379(.A(G93), .ZN(new_n805));
  INV_X1    g380(.A(G55), .ZN(new_n806));
  OAI22_X1  g381(.A1(new_n520), .A2(new_n805), .B1(new_n806), .B2(new_n523), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G860), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT37), .Z(new_n810));
  OR3_X1    g385(.A1(new_n555), .A2(new_n807), .A3(new_n804), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n555), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n601), .A2(G559), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n819));
  AOI21_X1  g394(.A(G860), .B1(new_n819), .B2(KEYINPUT97), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(KEYINPUT97), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n810), .B1(new_n821), .B2(new_n822), .ZN(G145));
  INV_X1    g398(.A(G37), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n491), .B(new_n622), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G160), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n510), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n495), .A2(new_n497), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n464), .A2(new_n501), .A3(G138), .A4(new_n504), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(KEYINPUT98), .A3(new_n500), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n791), .A2(new_n720), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n791), .A2(new_n720), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n838), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n833), .A2(KEYINPUT98), .A3(new_n500), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT98), .B1(new_n833), .B2(new_n500), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n495), .A2(new_n497), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n840), .A2(new_n836), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n747), .B1(new_n839), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n487), .A2(G130), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n482), .A2(G142), .ZN(new_n848));
  NOR2_X1   g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(new_n468), .B2(G118), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n615), .Z(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(new_n700), .Z(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n844), .B1(new_n840), .B2(new_n836), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n837), .A2(new_n838), .A3(new_n835), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n856), .A3(new_n748), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n846), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n854), .B1(new_n846), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n827), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(new_n858), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n826), .B1(new_n859), .B2(new_n861), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n824), .B(new_n860), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g441(.A1(new_n808), .A2(new_n604), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n611), .B(new_n813), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n600), .A2(G299), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n600), .A2(G299), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT100), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(KEYINPUT41), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n869), .A2(new_n870), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n873), .B1(new_n879), .B2(new_n868), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(G303), .B(G288), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G290), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(G305), .Z(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n881), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n867), .B1(new_n886), .B2(new_n604), .ZN(G295));
  OAI21_X1  g462(.A(new_n867), .B1(new_n886), .B2(new_n604), .ZN(G331));
  AOI21_X1  g463(.A(G301), .B1(new_n811), .B2(new_n812), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n811), .A2(new_n812), .A3(G301), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(G168), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(G286), .B1(new_n893), .B2(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n877), .A3(new_n874), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n894), .A3(new_n871), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n885), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n899));
  OR3_X1    g474(.A1(new_n898), .A2(new_n899), .A3(G37), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n885), .A3(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n898), .B2(G37), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT43), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n897), .B1(new_n896), .B2(KEYINPUT102), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n878), .B2(new_n895), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n884), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(KEYINPUT103), .B(new_n884), .C1(new_n905), .C2(new_n907), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n824), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n904), .B1(KEYINPUT43), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n912), .B2(KEYINPUT43), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n900), .A2(new_n918), .A3(new_n901), .A4(new_n902), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n911), .A2(new_n824), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n878), .A2(new_n906), .A3(new_n895), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n896), .A2(KEYINPUT102), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n897), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n924), .A2(new_n884), .B1(KEYINPUT103), .B2(new_n901), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  AND4_X1   g501(.A1(new_n916), .A2(new_n926), .A3(KEYINPUT44), .A4(new_n919), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n915), .B1(new_n920), .B2(new_n927), .ZN(G397));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n844), .B2(G1384), .ZN(new_n930));
  NAND2_X1  g505(.A1(G160), .A2(G40), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G2067), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n720), .B(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT106), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n747), .B(G1996), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n700), .B(new_n703), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(G290), .A2(G1986), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(KEYINPUT105), .ZN(new_n942));
  NAND2_X1  g517(.A1(G290), .A2(G1986), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n942), .B(new_n943), .Z(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(new_n932), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n679), .A2(G1976), .ZN(new_n946));
  INV_X1    g521(.A(G1976), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT52), .B1(G288), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT108), .B1(new_n844), .B2(G1384), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n835), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n931), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n931), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n835), .A2(new_n950), .A3(new_n951), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n950), .B1(new_n835), .B2(new_n951), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT110), .B1(new_n960), .B2(G8), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n946), .B(new_n948), .C1(new_n956), .C2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT49), .ZN(new_n964));
  NAND2_X1  g539(.A1(G305), .A2(G1981), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT111), .B(G1981), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(KEYINPUT49), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI211_X1 g545(.A(new_n963), .B(KEYINPUT49), .C1(new_n965), .C2(new_n967), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n956), .B2(new_n961), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n954), .B1(new_n953), .B2(new_n955), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n960), .A2(KEYINPUT110), .A3(G8), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n975), .A2(new_n976), .B1(G1976), .B2(new_n679), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n962), .B(new_n973), .C1(new_n974), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n958), .B2(new_n959), .ZN(new_n980));
  INV_X1    g555(.A(G2090), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n512), .A2(new_n951), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n957), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n929), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n835), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n957), .A3(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT107), .B(G1971), .Z(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n955), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(G303), .A2(G8), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n991), .B(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n978), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n958), .A2(new_n959), .A3(new_n979), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n931), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n512), .A2(new_n979), .A3(new_n951), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n949), .A2(KEYINPUT50), .A3(new_n952), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(KEYINPUT113), .A3(new_n957), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n999), .A2(new_n981), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(new_n989), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n993), .B1(new_n1004), .B2(new_n955), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n980), .A2(new_n957), .A3(new_n983), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(G2084), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(new_n931), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n982), .A2(new_n929), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n949), .A2(new_n929), .A3(new_n952), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(KEYINPUT114), .A3(new_n957), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1966), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1017), .A2(new_n955), .A3(G286), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n996), .A2(new_n1005), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT63), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT63), .B1(new_n990), .B2(new_n994), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n978), .A2(new_n995), .A3(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1019), .A2(new_n1020), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n995), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(new_n978), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n973), .A2(new_n947), .A3(new_n679), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1026), .A2(new_n967), .B1(new_n976), .B2(new_n975), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1023), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(G299), .B(KEYINPUT57), .ZN(new_n1029));
  INV_X1    g604(.A(new_n987), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT56), .B(G2072), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1034));
  INV_X1    g609(.A(G1956), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1029), .B(new_n1033), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1032), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1029), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1006), .A2(new_n761), .B1(new_n933), .B2(new_n953), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1040), .A2(new_n600), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT61), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1029), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1037), .B2(new_n1032), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1045), .B2(new_n1036), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n1050));
  INV_X1    g625(.A(G1996), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n985), .A2(new_n957), .A3(new_n1051), .A4(new_n986), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT58), .B(G1341), .Z(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n953), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1050), .B1(new_n1055), .B2(new_n555), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(KEYINPUT116), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n960), .A2(new_n1053), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n554), .B1(new_n1058), .B2(new_n1052), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1050), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1049), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1056), .A2(KEYINPUT116), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1060), .B1(new_n1059), .B2(new_n1050), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(new_n1064), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1046), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1040), .A2(KEYINPUT60), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT119), .B(new_n600), .C1(new_n1040), .C2(KEYINPUT60), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1006), .A2(new_n761), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n953), .A2(new_n933), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(KEYINPUT60), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(new_n601), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1071), .A2(KEYINPUT60), .A3(new_n600), .A4(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT118), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1040), .A2(new_n1078), .A3(KEYINPUT60), .A4(new_n600), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1068), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1067), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1037), .A2(new_n1044), .A3(new_n1032), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1039), .A2(KEYINPUT61), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1039), .A2(new_n1086), .A3(KEYINPUT61), .A4(new_n1083), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1042), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1961), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n985), .A2(new_n957), .A3(new_n770), .A4(new_n986), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1006), .A2(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n770), .A2(KEYINPUT53), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n469), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G40), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n478), .B2(new_n468), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n930), .A2(new_n986), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT54), .B1(new_n1100), .B2(KEYINPUT123), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1093), .B1(new_n1015), .B2(new_n1094), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT122), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1099), .B2(G171), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1107), .A3(G171), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1101), .A2(new_n1104), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1102), .A2(G301), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(KEYINPUT54), .C1(G301), .C2(new_n1099), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n996), .A2(new_n1005), .ZN(new_n1113));
  NAND2_X1  g688(.A1(G286), .A2(G8), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT120), .ZN(new_n1115));
  NAND2_X1  g690(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1115), .B(new_n1117), .C1(new_n1017), .C2(new_n955), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1007), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1013), .A2(KEYINPUT114), .A3(new_n957), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT114), .B1(new_n1013), .B2(new_n957), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1120), .A2(new_n1121), .A3(new_n1011), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1122), .B2(G1966), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(G8), .A3(new_n1116), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT51), .B(new_n1119), .C1(new_n1122), .C2(G1966), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1115), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1118), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1112), .A2(new_n1113), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1028), .B1(new_n1089), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1118), .A2(new_n1124), .A3(new_n1127), .A4(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1113), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1133), .A2(KEYINPUT124), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1135), .A2(new_n1134), .A3(new_n1113), .A4(new_n1132), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n945), .B1(new_n1130), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n932), .B1(new_n935), .B2(new_n747), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n932), .B(new_n1051), .C1(new_n1143), .C2(KEYINPUT46), .ZN(new_n1144));
  XOR2_X1   g719(.A(KEYINPUT126), .B(KEYINPUT46), .Z(new_n1145));
  INV_X1    g720(.A(new_n932), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(G1996), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT47), .Z(new_n1149));
  OR3_X1    g724(.A1(new_n937), .A2(new_n703), .A3(new_n701), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n720), .A2(G2067), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n932), .A2(new_n941), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT48), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1149), .B(new_n1154), .C1(new_n939), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1141), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g733(.A(G229), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n639), .A2(new_n458), .A3(new_n656), .ZN(new_n1161));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n1162));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g737(.A(new_n1163), .B1(new_n1162), .B2(new_n1161), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n913), .A2(new_n865), .A3(new_n1164), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


