//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n211), .A2(new_n212), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(new_n212), .B2(new_n211), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT66), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT67), .B(G77), .Z(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G58), .A2(G232), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n221), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n246), .B(KEYINPUT68), .Z(new_n247));
  INV_X1    g0047(.A(G107), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G97), .ZN(new_n249));
  INV_X1    g0049(.A(G97), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G107), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n247), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G274), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT69), .B(G45), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT75), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(KEYINPUT69), .A2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT69), .A2(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G41), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(KEYINPUT75), .B1(new_n265), .B2(new_n257), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n270), .B(new_n256), .C1(G41), .C2(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n267), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n262), .A2(new_n266), .B1(G238), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G97), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(G226), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n275), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n283), .A2(KEYINPUT74), .A3(new_n267), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT74), .B1(new_n283), .B2(new_n267), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n273), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT13), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT13), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n288), .B(new_n273), .C1(new_n284), .C2(new_n285), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(KEYINPUT76), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT76), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n286), .A2(new_n291), .A3(KEYINPUT13), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(G169), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT14), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT14), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n290), .A2(new_n295), .A3(G169), .A4(new_n292), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n287), .A2(G179), .A3(new_n289), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n242), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n214), .A2(G33), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n304), .A2(G77), .B1(G20), .B2(new_n242), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n202), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n213), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(KEYINPUT11), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n256), .B2(G20), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G68), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n302), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT11), .B1(new_n308), .B2(new_n310), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n298), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n290), .A2(G200), .A3(new_n292), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n286), .B2(KEYINPUT13), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n316), .B1(new_n320), .B2(new_n289), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n274), .A2(G222), .A3(new_n281), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n274), .A2(G1698), .ZN(new_n325));
  INV_X1    g0125(.A(G223), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n324), .B1(new_n222), .B2(new_n274), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n267), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n260), .B1(new_n272), .B2(G226), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(G190), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n204), .A2(G20), .ZN(new_n335));
  INV_X1    g0135(.A(G150), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT71), .B(G58), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT8), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(KEYINPUT8), .B2(G58), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n335), .B1(new_n336), .B2(new_n307), .C1(new_n303), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n310), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n299), .A2(G50), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n312), .B2(G50), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(KEYINPUT9), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT9), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n341), .B2(new_n343), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n334), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT10), .B1(new_n333), .B2(KEYINPUT73), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n349), .B(new_n334), .C1(new_n345), .C2(new_n347), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n344), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n331), .A2(G169), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n330), .A2(G179), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n260), .B1(new_n272), .B2(G232), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n278), .A2(new_n280), .A3(G226), .A4(G1698), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n278), .A2(new_n280), .A3(G223), .A4(new_n281), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G87), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n267), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n360), .A2(G190), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n332), .B1(new_n360), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n274), .B2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n278), .A2(new_n280), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n242), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G159), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n307), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n201), .B1(new_n337), .B2(G68), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n214), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n370), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n373), .B2(new_n214), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n371), .B(G20), .C1(new_n278), .C2(new_n280), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G58), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT71), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G58), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n216), .B1(new_n389), .B2(new_n242), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n377), .B1(new_n390), .B2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n384), .A2(new_n391), .A3(KEYINPUT16), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n381), .A2(new_n392), .A3(new_n310), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n339), .A2(new_n299), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n312), .B2(new_n339), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n368), .A2(new_n369), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n395), .ZN(new_n398));
  INV_X1    g0198(.A(G179), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n360), .A2(new_n399), .A3(new_n365), .ZN(new_n400));
  AOI21_X1  g0200(.A(G169), .B1(new_n360), .B2(new_n365), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT77), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G169), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n364), .A2(new_n267), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n269), .A2(new_n271), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G41), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(G1), .A3(G13), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(G232), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n260), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n403), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n360), .A2(new_n399), .A3(new_n365), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n398), .A2(new_n402), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n398), .A2(KEYINPUT18), .A3(new_n402), .A4(new_n414), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n397), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT15), .B(G87), .Z(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n303), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT8), .B(G58), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n222), .A2(new_n214), .B1(new_n424), .B2(new_n307), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n310), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n312), .A2(G77), .B1(new_n222), .B2(new_n300), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n274), .A2(G232), .A3(new_n281), .ZN(new_n429));
  INV_X1    g0229(.A(G238), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n429), .B1(new_n248), .B2(new_n274), .C1(new_n325), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n267), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n260), .B1(new_n272), .B2(G244), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n428), .B1(new_n435), .B2(new_n332), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT72), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n428), .C1(new_n435), .C2(new_n332), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n437), .B(new_n439), .C1(new_n319), .C2(new_n434), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n428), .B1(new_n434), .B2(new_n403), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(G179), .B2(new_n434), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR4_X1   g0243(.A1(new_n323), .A2(new_n359), .A3(new_n420), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G257), .A3(new_n407), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n446), .A2(new_n447), .A3(new_n449), .A4(G274), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n278), .A2(new_n280), .A3(G244), .A4(new_n281), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT4), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n461), .A2(new_n462), .A3(new_n267), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n461), .B2(new_n267), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n454), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT82), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT82), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n454), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(G200), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n299), .A2(G97), .ZN(new_n470));
  INV_X1    g0270(.A(new_n310), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT80), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n256), .A2(G33), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n471), .A2(new_n472), .A3(new_n299), .A4(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n299), .A2(new_n473), .A3(new_n213), .A4(new_n309), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT80), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n470), .B1(new_n477), .B2(G97), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n453), .B1(new_n461), .B2(new_n267), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n248), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT6), .ZN(new_n483));
  XNOR2_X1  g0283(.A(G97), .B(G107), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G77), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n485), .A2(new_n214), .B1(new_n486), .B2(new_n307), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n248), .B1(new_n372), .B2(new_n374), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n310), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT79), .ZN(new_n490));
  OAI21_X1  g0290(.A(G107), .B1(new_n382), .B2(new_n383), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n481), .B1(new_n252), .B2(KEYINPUT6), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(G20), .B1(G77), .B2(new_n306), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT79), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n495), .A3(new_n310), .ZN(new_n496));
  AOI221_X4 g0296(.A(new_n479), .B1(G190), .B2(new_n480), .C1(new_n490), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n469), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT89), .A2(G87), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n278), .A2(new_n280), .A3(new_n499), .A4(new_n214), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n274), .A2(new_n502), .A3(new_n214), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT90), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n214), .B2(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT23), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n505), .B(new_n508), .C1(new_n214), .C2(G107), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n507), .A2(new_n509), .B1(G116), .B2(new_n304), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n504), .A2(KEYINPUT24), .A3(new_n510), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n310), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n256), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n448), .A2(G41), .ZN(new_n517));
  OAI211_X1 g0317(.A(G264), .B(new_n407), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT92), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n450), .A2(KEYINPUT92), .A3(G264), .A4(new_n407), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n278), .A2(new_n280), .A3(G250), .A4(new_n281), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n278), .A2(new_n280), .A3(G257), .A4(G1698), .ZN(new_n524));
  XOR2_X1   g0324(.A(KEYINPUT91), .B(G294), .Z(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(new_n277), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n267), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n527), .A3(new_n452), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G200), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n477), .A2(G107), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n299), .A2(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT25), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n522), .A2(new_n527), .A3(G190), .A4(new_n452), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n515), .A2(new_n529), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT93), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n471), .B1(new_n511), .B2(new_n512), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n533), .B1(new_n539), .B2(new_n514), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(KEYINPUT93), .A3(new_n535), .A4(new_n529), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n495), .B1(new_n494), .B2(new_n310), .ZN(new_n543));
  AOI211_X1 g0343(.A(KEYINPUT79), .B(new_n471), .C1(new_n491), .C2(new_n493), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n478), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n399), .B(new_n454), .C1(new_n463), .C2(new_n464), .ZN(new_n546));
  INV_X1    g0346(.A(new_n480), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n403), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n477), .A2(new_n421), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n421), .A2(new_n299), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n214), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT84), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT84), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n556), .A3(new_n214), .ZN(new_n557));
  NOR4_X1   g0357(.A1(KEYINPUT85), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  INV_X1    g0360(.A(G87), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n555), .B(new_n557), .C1(new_n558), .C2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n278), .A2(new_n280), .A3(new_n214), .A4(G68), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n303), .B2(new_n250), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n550), .B(new_n552), .C1(new_n568), .C2(new_n471), .ZN(new_n569));
  OAI21_X1  g0369(.A(G250), .B1(new_n445), .B2(G1), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n267), .A2(new_n570), .B1(new_n445), .B2(new_n257), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n278), .A2(new_n280), .A3(G238), .A4(new_n281), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT83), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT83), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n274), .A2(new_n574), .A3(G238), .A4(new_n281), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n274), .A2(G244), .A3(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G116), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n573), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n571), .B1(new_n578), .B2(new_n267), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n399), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n569), .B(new_n580), .C1(G169), .C2(new_n579), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(G190), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n471), .B1(new_n563), .B2(new_n567), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n561), .B1(new_n474), .B2(new_n476), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n583), .A2(new_n584), .A3(new_n551), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n582), .B(new_n585), .C1(new_n332), .C2(new_n579), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n498), .A2(new_n542), .A3(new_n549), .A4(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n274), .A2(G257), .A3(new_n281), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n373), .A2(G303), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n278), .A2(new_n280), .A3(G264), .A4(G1698), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n267), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n450), .A2(G270), .A3(new_n407), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n595), .A2(KEYINPUT86), .A3(new_n452), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT86), .B1(new_n595), .B2(new_n452), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G169), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n300), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n475), .B2(new_n600), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n459), .B(new_n214), .C1(G33), .C2(new_n250), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(G20), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n310), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n604), .B1(new_n310), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT20), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(KEYINPUT20), .B(new_n603), .C1(new_n606), .C2(new_n607), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n602), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n589), .B1(new_n599), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT88), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT88), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n589), .C1(new_n599), .C2(new_n612), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n598), .A2(new_n399), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n589), .B2(new_n599), .ZN(new_n619));
  INV_X1    g0419(.A(new_n612), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n528), .A2(G179), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n403), .B2(new_n528), .ZN(new_n623));
  INV_X1    g0423(.A(new_n540), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n598), .A2(G200), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n626), .B(new_n612), .C1(new_n319), .C2(new_n598), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n617), .A2(new_n621), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n588), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n444), .A2(new_n629), .ZN(G372));
  INV_X1    g0430(.A(KEYINPUT94), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n588), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n490), .A2(new_n496), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(new_n478), .B1(new_n403), .B2(new_n547), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n469), .A2(new_n497), .B1(new_n634), .B2(new_n546), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n581), .A2(new_n586), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n538), .B2(new_n541), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(KEYINPUT94), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n617), .A2(new_n621), .A3(new_n625), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT95), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n617), .A2(KEYINPUT95), .A3(new_n621), .A4(new_n625), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n632), .A2(new_n638), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n581), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n587), .A2(KEYINPUT26), .A3(new_n546), .A4(new_n634), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n549), .B2(new_n636), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n444), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT96), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n317), .A2(new_n442), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n322), .A3(new_n397), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n419), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n353), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n651), .B1(new_n655), .B2(new_n358), .ZN(new_n656));
  AOI211_X1 g0456(.A(KEYINPUT96), .B(new_n357), .C1(new_n654), .C2(new_n353), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n650), .B1(new_n656), .B2(new_n657), .ZN(G369));
  NAND2_X1  g0458(.A1(new_n617), .A2(new_n621), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n214), .A2(G13), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n256), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n612), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n659), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n627), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n625), .A2(new_n667), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT97), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n624), .B1(new_n623), .B2(new_n666), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n542), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n659), .A2(new_n667), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n625), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n667), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT98), .ZN(G399));
  INV_X1    g0486(.A(new_n210), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OR3_X1    g0489(.A1(new_n558), .A2(new_n562), .A3(G116), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n689), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n217), .B2(new_n689), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n666), .B1(new_n643), .B2(new_n648), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n639), .A2(new_n635), .A3(new_n637), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n666), .B1(new_n697), .B2(new_n648), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n629), .A2(new_n667), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n522), .A2(new_n527), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(new_n480), .A3(new_n579), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n703), .B1(new_n618), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n579), .B1(new_n704), .B2(new_n452), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n465), .A3(new_n399), .A4(new_n598), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n618), .A2(new_n705), .A3(new_n703), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n666), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT31), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n701), .B1(new_n702), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n700), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n694), .B1(new_n716), .B2(G1), .ZN(G364));
  NOR3_X1   g0517(.A1(new_n319), .A2(G179), .A3(G200), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n214), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n250), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n399), .A2(new_n332), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n214), .A2(new_n319), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n214), .A2(G190), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G179), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G159), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n274), .B1(new_n202), .B2(new_n723), .C1(new_n728), .C2(KEYINPUT32), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n720), .B(new_n729), .C1(KEYINPUT32), .C2(new_n728), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n332), .A2(G179), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n722), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n561), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n721), .A2(new_n724), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n724), .A2(new_n731), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n242), .B1(new_n735), .B2(new_n248), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n724), .A2(G179), .A3(new_n332), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n733), .B(new_n736), .C1(new_n223), .C2(new_n738), .ZN(new_n739));
  NOR4_X1   g0539(.A1(new_n214), .A2(new_n399), .A3(new_n319), .A4(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT101), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(KEYINPUT101), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n730), .B(new_n739), .C1(new_n389), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n734), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT33), .B(G317), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(new_n727), .B2(G329), .ZN(new_n748));
  INV_X1    g0548(.A(G283), .ZN(new_n749));
  INV_X1    g0549(.A(G322), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n748), .B1(new_n749), .B2(new_n735), .C1(new_n750), .C2(new_n741), .ZN(new_n751));
  INV_X1    g0551(.A(new_n723), .ZN(new_n752));
  INV_X1    g0552(.A(new_n732), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G326), .A2(new_n752), .B1(new_n753), .B2(G303), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n274), .B1(new_n738), .B2(G311), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(new_n525), .C2(new_n719), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n745), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n213), .B1(G20), .B2(new_n403), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OR3_X1    g0559(.A1(KEYINPUT100), .A2(G13), .A3(G33), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT100), .B1(G13), .B2(G33), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n758), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n246), .A2(new_n445), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n687), .A2(new_n274), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n766), .B(new_n768), .C1(new_n218), .C2(new_n258), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n210), .A2(new_n274), .ZN(new_n770));
  INV_X1    g0570(.A(G355), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(G116), .B2(new_n210), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n765), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n256), .B1(new_n660), .B2(G45), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n689), .A2(KEYINPUT99), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT99), .ZN(new_n776));
  INV_X1    g0576(.A(new_n774), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n688), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n759), .A2(new_n773), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT102), .Z(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n670), .B2(new_n764), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n673), .A2(new_n780), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n671), .A2(G330), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n783), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NOR2_X1   g0588(.A1(new_n442), .A2(new_n666), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n440), .B1(new_n428), .B2(new_n667), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n442), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n695), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n649), .A2(new_n667), .A3(new_n791), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n780), .B1(new_n794), .B2(new_n714), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n714), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n762), .A2(new_n758), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n738), .A2(G116), .B1(new_n740), .B2(G294), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n799), .B(new_n373), .C1(new_n561), .C2(new_n735), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n734), .A2(new_n749), .B1(new_n726), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n723), .A2(new_n803), .B1(new_n732), .B2(new_n248), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n800), .A2(new_n720), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n752), .A2(G137), .B1(new_n738), .B2(G159), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n336), .B2(new_n734), .ZN(new_n807));
  INV_X1    g0607(.A(new_n744), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(G143), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT34), .Z(new_n810));
  AOI21_X1  g0610(.A(new_n373), .B1(new_n727), .B2(G132), .ZN(new_n811));
  INV_X1    g0611(.A(new_n735), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G68), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n811), .B(new_n813), .C1(new_n202), .C2(new_n732), .ZN(new_n814));
  INV_X1    g0614(.A(new_n719), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n337), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT103), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n805), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n758), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n780), .B1(G77), .B2(new_n798), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT104), .Z(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n763), .B2(new_n791), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n796), .A2(new_n822), .ZN(G384));
  NOR2_X1   g0623(.A1(new_n660), .A2(new_n256), .ZN(new_n824));
  INV_X1    g0624(.A(new_n664), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n398), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n368), .A2(new_n393), .A3(new_n395), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT37), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT107), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n415), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n398), .A2(KEYINPUT107), .A3(new_n402), .A4(new_n414), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n829), .A2(new_n830), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n402), .A2(new_n414), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT106), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT16), .B1(new_n384), .B2(new_n391), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n837), .B2(new_n471), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n381), .A2(KEYINPUT106), .A3(new_n310), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(new_n392), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n835), .B1(new_n395), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n664), .B1(new_n840), .B2(new_n395), .ZN(new_n842));
  INV_X1    g0642(.A(new_n827), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n834), .B1(new_n844), .B2(new_n830), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n417), .A2(new_n418), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT17), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n396), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n842), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT108), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT108), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n845), .A2(new_n849), .A3(new_n852), .A4(KEYINPUT38), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n420), .A2(new_n398), .A3(new_n825), .ZN(new_n855));
  INV_X1    g0655(.A(new_n415), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n856), .B2(new_n828), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n834), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n316), .A2(new_n666), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n317), .A2(new_n322), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n298), .A2(new_n316), .A3(new_n666), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n790), .A2(new_n442), .ZN(new_n866));
  INV_X1    g0666(.A(new_n789), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n712), .B2(new_n702), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n861), .A2(KEYINPUT40), .A3(new_n865), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n845), .A2(new_n849), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n850), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(new_n869), .A3(new_n865), .ZN(new_n875));
  XOR2_X1   g0675(.A(KEYINPUT110), .B(KEYINPUT40), .Z(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n588), .A2(new_n628), .A3(new_n666), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n711), .B(KEYINPUT31), .Z(new_n880));
  OAI21_X1  g0680(.A(new_n444), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n870), .A2(new_n877), .A3(G330), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n444), .A2(new_n713), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n696), .A2(new_n444), .A3(new_n699), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n656), .B2(new_n657), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n885), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n317), .A2(new_n666), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n840), .A2(new_n395), .ZN(new_n891));
  INV_X1    g0691(.A(new_n835), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n825), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n827), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n896), .A2(new_n834), .B1(new_n420), .B2(new_n842), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n852), .B1(new_n897), .B2(KEYINPUT38), .ZN(new_n898));
  AND4_X1   g0698(.A1(new_n852), .A2(new_n845), .A3(KEYINPUT38), .A4(new_n849), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n890), .B(new_n860), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT109), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n902), .B1(new_n900), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n889), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n789), .B1(new_n695), .B2(new_n791), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n863), .A2(new_n864), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n908), .A2(new_n874), .B1(new_n846), .B2(new_n664), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n824), .B1(new_n888), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n911), .B2(new_n888), .ZN(new_n913));
  OAI211_X1 g0713(.A(G116), .B(new_n215), .C1(new_n492), .C2(KEYINPUT35), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(KEYINPUT35), .B2(new_n492), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  OAI211_X1 g0716(.A(new_n223), .B(new_n218), .C1(new_n242), .C2(new_n389), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n256), .B(G13), .C1(new_n917), .C2(new_n241), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT105), .Z(new_n919));
  NAND3_X1  g0719(.A1(new_n913), .A2(new_n916), .A3(new_n919), .ZN(G367));
  NAND2_X1  g0720(.A1(new_n498), .A2(new_n683), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n666), .B1(new_n921), .B2(new_n549), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n545), .A2(new_n666), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n635), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n634), .A2(new_n546), .A3(new_n666), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n682), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n927), .B2(KEYINPUT42), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(KEYINPUT42), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n585), .A2(new_n667), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n644), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n636), .B2(new_n930), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n926), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n680), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n937), .B(new_n939), .Z(new_n940));
  XNOR2_X1  g0740(.A(new_n688), .B(KEYINPUT41), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n678), .B(new_n681), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n673), .B1(new_n943), .B2(KEYINPUT112), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(KEYINPUT112), .B2(new_n943), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n945), .A2(new_n680), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n946), .A2(new_n716), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT111), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n678), .A2(new_n681), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n625), .B2(new_n666), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n949), .B1(new_n951), .B2(new_n938), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n684), .A2(KEYINPUT45), .A3(new_n926), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT44), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n684), .B2(new_n926), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(KEYINPUT44), .A3(new_n938), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n954), .A2(new_n958), .A3(new_n680), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n680), .B1(new_n954), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n948), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n947), .B(new_n961), .C1(new_n948), .C2(new_n960), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n942), .B1(new_n962), .B2(new_n716), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n940), .B1(new_n963), .B2(new_n777), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n768), .A2(new_n239), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n765), .B1(new_n210), .B2(new_n422), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n780), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n202), .A2(new_n737), .B1(new_n734), .B2(new_n376), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n373), .B(new_n968), .C1(new_n337), .C2(new_n753), .ZN(new_n969));
  AOI22_X1  g0769(.A1(G137), .A2(new_n727), .B1(new_n740), .B2(G150), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G143), .A2(new_n752), .B1(new_n223), .B2(new_n812), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n815), .A2(G68), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT114), .B(G317), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n727), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n525), .B2(new_n734), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n373), .B1(new_n735), .B2(new_n250), .C1(new_n719), .C2(new_n248), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n723), .A2(new_n801), .B1(new_n737), .B2(new_n749), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n803), .B2(new_n744), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT113), .B1(new_n732), .B2(new_n600), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n973), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT47), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n819), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n967), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n764), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n988), .B2(new_n932), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n964), .A2(new_n989), .ZN(G387));
  NAND2_X1  g0790(.A1(new_n946), .A2(new_n777), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n770), .A2(new_n691), .B1(G107), .B2(new_n210), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT115), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n445), .B1(new_n242), .B2(new_n486), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n424), .A2(G50), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT50), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n691), .B(new_n997), .C1(new_n996), .C2(new_n995), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n998), .B(new_n767), .C1(new_n236), .C2(new_n258), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n779), .B1(new_n1000), .B2(new_n765), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G150), .A2(new_n727), .B1(new_n740), .B2(G50), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n376), .B2(new_n723), .C1(new_n339), .C2(new_n734), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n815), .A2(new_n421), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n373), .B1(new_n812), .B2(G97), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n738), .A2(G68), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n223), .A2(new_n753), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n737), .A2(new_n803), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n723), .A2(new_n750), .B1(new_n734), .B2(new_n801), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(new_n808), .C2(new_n974), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT48), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n749), .B2(new_n719), .C1(new_n525), .C2(new_n732), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT49), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n274), .B1(new_n727), .B2(G326), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n600), .B2(new_n735), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1009), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1001), .B1(new_n679), .B2(new_n988), .C1(new_n1020), .C2(new_n819), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n947), .A2(new_n689), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n946), .A2(new_n716), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n991), .B(new_n1021), .C1(new_n1022), .C2(new_n1023), .ZN(G393));
  NOR2_X1   g0824(.A1(new_n959), .A2(new_n960), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n962), .B(new_n688), .C1(new_n947), .C2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n926), .A2(new_n988), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT116), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT116), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n768), .A2(new_n254), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n765), .B1(new_n250), .B2(new_n210), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n780), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n749), .A2(new_n732), .B1(new_n734), .B2(new_n803), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n752), .A2(G317), .B1(new_n740), .B2(G311), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT52), .ZN(new_n1036));
  INV_X1    g0836(.A(G294), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n737), .A2(new_n1037), .B1(new_n726), .B2(new_n750), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n373), .B1(new_n735), .B2(new_n248), .C1(new_n719), .C2(new_n600), .ZN(new_n1039));
  OR4_X1    g0839(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n424), .A2(new_n737), .B1(new_n734), .B2(new_n202), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n719), .A2(new_n486), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT118), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n741), .A2(new_n376), .B1(new_n723), .B2(new_n336), .ZN(new_n1045));
  XOR2_X1   g0845(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n373), .B1(new_n812), .B2(G87), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G68), .A2(new_n753), .B1(new_n727), .B2(G143), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1040), .B1(new_n1044), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1033), .B1(new_n758), .B2(new_n1053), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n1029), .A2(new_n1030), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1025), .B2(new_n777), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1026), .A2(new_n1056), .ZN(G390));
  OAI211_X1 g0857(.A(new_n886), .B(new_n884), .C1(new_n656), .C2(new_n657), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n713), .A2(new_n865), .A3(new_n791), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT120), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT120), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n713), .A2(new_n865), .A3(new_n1062), .A4(new_n791), .ZN(new_n1063));
  OAI211_X1 g0863(.A(G330), .B(new_n791), .C1(new_n880), .C2(new_n879), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n907), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n793), .A2(new_n867), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n697), .A2(new_n648), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(new_n667), .A3(new_n866), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1060), .A2(new_n867), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n1065), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1059), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT119), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n889), .B1(new_n854), .B2(new_n860), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1070), .A2(new_n867), .B1(new_n863), .B2(new_n864), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n859), .B1(new_n851), .B2(new_n853), .ZN(new_n1080));
  NOR4_X1   g0880(.A1(new_n1080), .A2(new_n1077), .A3(KEYINPUT119), .A4(new_n889), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(KEYINPUT39), .B(new_n859), .C1(new_n851), .C2(new_n853), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n890), .B1(new_n873), .B2(new_n850), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT109), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n900), .A2(new_n902), .A3(new_n901), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n889), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n906), .B2(new_n907), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1082), .A2(new_n1089), .A3(new_n1060), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1074), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n889), .B1(new_n1067), .B2(new_n865), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n903), .A2(new_n1095), .A3(new_n904), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n861), .A2(new_n1078), .A3(new_n1087), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT119), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1076), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1091), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1066), .A2(new_n1067), .B1(new_n1071), .B2(new_n1065), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1058), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1082), .A2(new_n1089), .A3(new_n1060), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1094), .A2(new_n1105), .A3(new_n688), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G137), .A2(new_n746), .B1(new_n740), .B2(G132), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n726), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT53), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n732), .B2(new_n336), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n753), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(G128), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n274), .B1(new_n723), .B2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT54), .B(G143), .Z(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1117), .A2(new_n737), .B1(new_n735), .B2(new_n202), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1115), .B(new_n1118), .C1(G159), .C2(new_n815), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT121), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n723), .A2(new_n749), .B1(new_n737), .B2(new_n250), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G107), .B2(new_n746), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT122), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n813), .B1(new_n1037), .B2(new_n726), .C1(new_n600), .C2(new_n741), .ZN(new_n1125));
  OR3_X1    g0925(.A1(new_n1042), .A2(new_n274), .A3(new_n733), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n758), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n779), .B1(new_n339), .B2(new_n797), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT123), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n903), .A2(new_n904), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n762), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n777), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT124), .B1(new_n1106), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1106), .A2(new_n1135), .A3(KEYINPUT124), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(G378));
  NOR2_X1   g0939(.A1(new_n354), .A2(new_n664), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n359), .B(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1141), .B(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n883), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1144), .A2(G330), .A3(new_n877), .A4(new_n870), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n910), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n905), .A3(new_n1147), .A4(new_n909), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1145), .A2(new_n762), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n780), .B1(G50), .B2(new_n798), .ZN(new_n1153));
  INV_X1    g0953(.A(G132), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n741), .A2(new_n1114), .B1(new_n734), .B2(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G137), .A2(new_n738), .B1(new_n753), .B2(new_n1116), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1108), .B2(new_n723), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G150), .C2(new_n815), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT59), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n812), .A2(G159), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G33), .B(G41), .C1(new_n727), .C2(G124), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n735), .A2(new_n389), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G107), .B2(new_n740), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n274), .A2(G41), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1166), .A2(new_n972), .A3(new_n1007), .A4(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n723), .A2(new_n600), .B1(new_n726), .B2(new_n749), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n422), .A2(new_n737), .B1(new_n734), .B2(new_n250), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1167), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1164), .A2(new_n1172), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1153), .B1(new_n1176), .B2(new_n758), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1151), .A2(new_n777), .B1(new_n1152), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1105), .A2(new_n1059), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n1151), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n688), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1105), .A2(new_n1059), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(KEYINPUT57), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1178), .B1(new_n1181), .B2(new_n1183), .ZN(G375));
  NAND2_X1  g0984(.A1(new_n1058), .A2(new_n1102), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1074), .A2(new_n941), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n907), .A2(new_n762), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n798), .A2(G68), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G132), .A2(new_n752), .B1(new_n753), .B2(G159), .ZN(new_n1189));
  INV_X1    g0989(.A(G137), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1189), .B1(new_n1114), .B2(new_n726), .C1(new_n744), .C2(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1117), .A2(new_n734), .B1(new_n737), .B2(new_n336), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1192), .A2(new_n373), .A3(new_n1165), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n202), .B2(new_n719), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n738), .A2(G107), .B1(new_n746), .B2(G116), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n250), .B2(new_n732), .C1(new_n1037), .C2(new_n723), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G303), .A2(new_n727), .B1(new_n740), .B2(G283), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n274), .B1(new_n812), .B2(G77), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n1004), .A3(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n1191), .A2(new_n1194), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1188), .B(new_n779), .C1(new_n1200), .C2(new_n758), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1073), .A2(new_n777), .B1(new_n1187), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1186), .A2(new_n1202), .ZN(G381));
  OR4_X1    g1003(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1204), .A2(G387), .A3(G381), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1106), .A2(new_n1135), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(G375), .A2(KEYINPUT125), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(G375), .A2(KEYINPUT125), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(G407));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n665), .A2(G213), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT126), .Z(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G407), .B(G213), .C1(new_n1211), .C2(new_n1214), .ZN(G409));
  NAND2_X1  g1015(.A1(new_n1182), .A2(new_n941), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1178), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1207), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1106), .A2(new_n1135), .A3(KEYINPUT124), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(new_n1136), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(G375), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT60), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1185), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1058), .A2(new_n1102), .A3(KEYINPUT60), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1223), .A2(new_n688), .A3(new_n1074), .A4(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1225), .A2(G384), .A3(new_n1202), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G384), .B1(new_n1225), .B2(new_n1202), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1221), .A2(new_n1214), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT62), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT61), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT62), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1221), .A2(new_n1232), .A3(new_n1214), .A4(new_n1228), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1213), .A2(G2897), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT127), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1227), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1225), .A2(G384), .A3(new_n1202), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1235), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT127), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1236), .B1(new_n1234), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1178), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1182), .A2(KEYINPUT57), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n689), .B1(new_n1182), .B2(KEYINPUT57), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1246), .A2(G378), .B1(new_n1207), .B2(new_n1217), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1242), .B1(new_n1247), .B2(new_n1213), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1230), .A2(new_n1231), .A3(new_n1233), .A4(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(G393), .B(new_n787), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n964), .A2(new_n989), .A3(G390), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G390), .B1(new_n964), .B2(new_n989), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1251), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1254), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n1250), .A3(new_n1252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1249), .A2(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1221), .A2(new_n1214), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1242), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1221), .A2(KEYINPUT63), .A3(new_n1214), .A4(new_n1228), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1229), .A2(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1260), .A2(new_n1262), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1259), .A2(new_n1266), .ZN(G405));
  NAND2_X1  g1067(.A1(new_n1246), .A2(G378), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G375), .A2(new_n1207), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(new_n1228), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1228), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1260), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1258), .B1(new_n1273), .B2(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(G402));
endmodule


