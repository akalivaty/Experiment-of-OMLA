//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G478), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT15), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT87), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT78), .B(G107), .ZN(new_n190));
  XNOR2_X1  g004(.A(G116), .B(G122), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  INV_X1    g009(.A(G122), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n197), .B2(KEYINPUT14), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n189), .A2(new_n192), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G134), .ZN(new_n200));
  XNOR2_X1  g014(.A(G128), .B(G143), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n199), .B(new_n202), .C1(new_n189), .C2(new_n192), .ZN(new_n203));
  XNOR2_X1  g017(.A(new_n190), .B(new_n191), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n201), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT13), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(G143), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n208), .A2(KEYINPUT86), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n208), .A2(new_n209), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT86), .B1(new_n213), .B2(new_n206), .ZN(new_n214));
  OAI21_X1  g028(.A(G134), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n204), .B(new_n205), .C1(new_n210), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT9), .B(G234), .ZN(new_n218));
  INV_X1    g032(.A(G217), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n218), .A2(new_n219), .A3(G953), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT88), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n203), .A2(new_n216), .A3(new_n223), .A4(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n221), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n226), .A2(KEYINPUT89), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT89), .B1(new_n226), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n188), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n229), .A2(new_n188), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G475), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT71), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G953), .ZN(new_n237));
  INV_X1    g051(.A(G237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n235), .A2(new_n237), .A3(G214), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n212), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT71), .B(G953), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n241), .A2(G143), .A3(G214), .A4(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT18), .A3(G131), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  XNOR2_X1  g059(.A(G125), .B(G140), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G140), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G125), .ZN(new_n250));
  INV_X1    g064(.A(G125), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G140), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(KEYINPUT77), .ZN(new_n254));
  OAI22_X1  g068(.A1(new_n248), .A2(new_n254), .B1(new_n245), .B2(new_n246), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT18), .A2(G131), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n240), .A2(new_n242), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n244), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G113), .B(G122), .ZN(new_n259));
  INV_X1    g073(.A(G104), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n240), .A2(new_n242), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n240), .B2(new_n242), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT17), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n243), .A2(KEYINPUT17), .A3(G131), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT16), .ZN(new_n269));
  OR3_X1    g083(.A1(new_n251), .A2(KEYINPUT16), .A3(G140), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G146), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(G146), .B1(new_n269), .B2(new_n270), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n258), .B(new_n263), .C1(new_n267), .C2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n268), .A2(new_n274), .ZN(new_n277));
  INV_X1    g091(.A(new_n266), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT17), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n240), .A2(new_n242), .A3(new_n264), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n255), .A2(new_n257), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n277), .A2(new_n281), .B1(new_n282), .B2(new_n244), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n276), .B1(new_n283), .B2(new_n261), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n233), .B1(new_n284), .B2(new_n227), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT20), .ZN(new_n287));
  INV_X1    g101(.A(new_n258), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT82), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n247), .B1(new_n289), .B2(KEYINPUT19), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n253), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n246), .B2(new_n247), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT19), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n271), .B1(new_n294), .B2(G146), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n295), .A2(KEYINPUT83), .B1(new_n278), .B2(new_n280), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT83), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n271), .C1(new_n294), .C2(G146), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n288), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n276), .B1(new_n299), .B2(new_n261), .ZN(new_n300));
  NOR2_X1   g114(.A1(G475), .A2(G902), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n287), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n247), .B1(new_n250), .B2(new_n252), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n293), .B1(new_n303), .B2(KEYINPUT82), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n253), .A2(new_n290), .ZN(new_n305));
  AOI21_X1  g119(.A(G146), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT83), .B1(new_n306), .B2(new_n272), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n278), .A2(new_n280), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n298), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n261), .B1(new_n309), .B2(new_n258), .ZN(new_n310));
  INV_X1    g124(.A(new_n276), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n287), .B(new_n301), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n286), .B1(new_n302), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n286), .B(KEYINPUT85), .C1(new_n302), .C2(new_n313), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n232), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G221), .B1(new_n218), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G469), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(new_n227), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n241), .A2(G227), .ZN(new_n323));
  XOR2_X1   g137(.A(G110), .B(G140), .Z(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n195), .A2(KEYINPUT78), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G107), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n328), .A3(G104), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n195), .A2(G104), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT3), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(new_n260), .B2(G107), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G101), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G101), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n330), .B1(new_n190), .B2(G104), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n336), .B(new_n333), .C1(new_n337), .C2(KEYINPUT3), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n338), .A3(KEYINPUT4), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n245), .A2(G143), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n212), .A2(G146), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT0), .A2(G128), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT0), .A2(G128), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G143), .B(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n343), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(G101), .C1(new_n332), .C2(new_n334), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n339), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n190), .A2(G104), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n260), .A2(G107), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G128), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT68), .B1(new_n342), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT68), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n347), .A2(new_n359), .A3(new_n356), .A4(G128), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n340), .A2(KEYINPUT1), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n347), .B1(G128), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n338), .B(new_n355), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n338), .A2(new_n355), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n358), .A2(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT69), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(KEYINPUT1), .C1(new_n212), .C2(G146), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G128), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n369), .B1(new_n340), .B2(KEYINPUT1), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n342), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n365), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n352), .A2(new_n366), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G137), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT11), .ZN(new_n378));
  INV_X1    g192(.A(G134), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT64), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT64), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G134), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(KEYINPUT11), .A3(G134), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT11), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G137), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n383), .A2(new_n264), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT65), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n384), .A2(new_n386), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n390), .A2(KEYINPUT65), .A3(new_n383), .A4(new_n264), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n383), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G131), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n376), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n389), .A2(new_n391), .B1(G131), .B2(new_n393), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n365), .A2(new_n364), .B1(new_n367), .B2(new_n374), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n398), .B2(new_n352), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n325), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n338), .A2(new_n355), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n362), .A2(KEYINPUT69), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(G128), .A3(new_n370), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n403), .A2(new_n342), .B1(new_n360), .B2(new_n358), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n364), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n395), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT12), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n398), .A2(new_n397), .A3(new_n352), .ZN(new_n409));
  INV_X1    g223(.A(new_n325), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT12), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n411), .A3(new_n395), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n408), .A2(new_n409), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n400), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n322), .B1(new_n414), .B2(new_n321), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n406), .B2(new_n395), .ZN(new_n416));
  AOI211_X1 g230(.A(KEYINPUT12), .B(new_n397), .C1(new_n405), .C2(new_n364), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n409), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n325), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n376), .A2(new_n395), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n409), .A3(new_n410), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(G469), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n320), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G116), .B(G119), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(KEYINPUT70), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT2), .B(G113), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n339), .A2(new_n428), .A3(new_n351), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(KEYINPUT5), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n431));
  INV_X1    g245(.A(G119), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(G116), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(G113), .ZN(new_n434));
  INV_X1    g248(.A(new_n427), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n430), .A2(new_n434), .B1(new_n435), .B2(new_n425), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n338), .A2(new_n355), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT79), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n439), .B(KEYINPUT79), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n429), .A2(new_n443), .A3(new_n437), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n438), .A2(new_n446), .A3(new_n441), .ZN(new_n447));
  INV_X1    g261(.A(G224), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(G953), .ZN(new_n449));
  AOI21_X1  g263(.A(G125), .B1(new_n368), .B2(new_n373), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n251), .B1(new_n346), .B2(new_n348), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n449), .ZN(new_n453));
  INV_X1    g267(.A(new_n451), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n453), .B(new_n454), .C1(new_n404), .C2(G125), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(new_n447), .A3(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n428), .A2(new_n351), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n458), .A2(new_n339), .B1(new_n367), .B2(new_n436), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT8), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n443), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n441), .A2(KEYINPUT8), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n435), .A2(new_n425), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT80), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n430), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n434), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n430), .A2(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n463), .B1(new_n367), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n401), .A2(new_n436), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n459), .A2(new_n443), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n453), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n452), .A2(new_n455), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n450), .A2(new_n451), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n473), .A3(new_n453), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(G902), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n457), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n481), .B(KEYINPUT81), .Z(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n457), .A2(new_n479), .A3(new_n482), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n234), .A2(G952), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(G234), .B2(G237), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n227), .B(new_n241), .C1(G234), .C2(G237), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT21), .B(G898), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n318), .A2(new_n424), .A3(new_n488), .A4(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT28), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n381), .A2(G134), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n379), .A2(KEYINPUT64), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n497), .B(new_n377), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G131), .ZN(new_n501));
  AOI21_X1  g315(.A(G137), .B1(new_n380), .B2(new_n382), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n497), .B1(new_n379), .B2(G137), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT67), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n368), .A2(new_n373), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n503), .B1(new_n200), .B2(G137), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n500), .A4(G131), .ZN(new_n510));
  AND4_X1   g324(.A1(new_n392), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n349), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n392), .B2(new_n394), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n428), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n395), .A2(new_n349), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n392), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n516));
  INV_X1    g330(.A(new_n428), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n496), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n518), .A2(new_n496), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n241), .A2(G210), .A3(new_n238), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT26), .B(G101), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT29), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n227), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n519), .B2(new_n521), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n511), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n515), .B2(new_n516), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n428), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n527), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n518), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT29), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G472), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n535), .B1(new_n519), .B2(new_n521), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT30), .B1(new_n511), .B2(new_n513), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n515), .A2(new_n532), .A3(new_n516), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n517), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n518), .A2(new_n527), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT31), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  INV_X1    g359(.A(new_n543), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n534), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n539), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT32), .ZN(new_n549));
  NOR2_X1   g363(.A1(G472), .A2(G902), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n538), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n219), .B1(G234), .B2(new_n227), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n241), .A2(G221), .A3(G234), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT22), .B(G137), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G119), .B(G128), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT73), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT74), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT24), .B(G110), .ZN(new_n563));
  OR3_X1    g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT75), .B1(new_n432), .B2(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT23), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n432), .A2(G128), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT23), .ZN(new_n570));
  OAI211_X1 g384(.A(KEYINPUT75), .B(new_n570), .C1(new_n432), .C2(G128), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n274), .B1(G110), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n248), .A2(new_n254), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n271), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n561), .A2(new_n563), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n572), .A2(G110), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT76), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT76), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n576), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n559), .B1(new_n574), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n582), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n581), .B1(new_n577), .B2(new_n578), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n271), .B(new_n575), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n566), .A2(new_n573), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n558), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(new_n589), .A3(new_n227), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n584), .A2(new_n589), .A3(KEYINPUT25), .A4(new_n227), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n555), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n584), .A2(new_n589), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n554), .A2(G902), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n553), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n495), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n336), .ZN(G3));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n548), .B2(new_n227), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n548), .B2(new_n550), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n487), .A2(new_n493), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n597), .A4(new_n424), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n310), .A2(new_n311), .ZN(new_n606));
  INV_X1    g420(.A(new_n301), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT20), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n285), .B1(new_n608), .B2(new_n312), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n315), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n217), .A2(KEYINPUT90), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n612), .B2(new_n220), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n220), .B2(new_n612), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n226), .A2(new_n611), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n187), .A2(G902), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n226), .A2(new_n227), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n616), .A2(new_n618), .B1(G478), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n605), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  NAND2_X1  g438(.A1(new_n232), .A2(new_n609), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n605), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT35), .B(G107), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NOR2_X1   g442(.A1(new_n574), .A2(new_n583), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n596), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n594), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n603), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n495), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT91), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  NAND2_X1  g453(.A1(new_n414), .A2(new_n321), .ZN(new_n640));
  INV_X1    g454(.A(new_n322), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n423), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n457), .A2(new_n479), .A3(new_n482), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n482), .B1(new_n457), .B2(new_n479), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND4_X1   g459(.A1(new_n485), .A2(new_n642), .A3(new_n645), .A4(new_n319), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n491), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n490), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n625), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n646), .A2(new_n553), .A3(new_n634), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  INV_X1    g466(.A(KEYINPUT92), .ZN(new_n653));
  INV_X1    g467(.A(new_n518), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n527), .B1(new_n542), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n514), .A2(new_n518), .A3(new_n535), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(new_n227), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n653), .B1(new_n658), .B2(G472), .ZN(new_n659));
  AOI211_X1 g473(.A(KEYINPUT92), .B(new_n601), .C1(new_n655), .C2(new_n657), .ZN(new_n660));
  OAI22_X1  g474(.A1(new_n551), .A2(new_n552), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT93), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI221_X1 g477(.A(KEYINPUT93), .B1(new_n659), .B2(new_n660), .C1(new_n551), .C2(new_n552), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n649), .B(KEYINPUT39), .Z(new_n666));
  AND2_X1   g480(.A1(new_n424), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT40), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n645), .B(KEYINPUT38), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n316), .A2(new_n317), .A3(new_n232), .ZN(new_n670));
  INV_X1    g484(.A(new_n485), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n634), .A3(new_n671), .ZN(new_n672));
  AND4_X1   g486(.A1(new_n665), .A2(new_n668), .A3(new_n669), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n212), .ZN(G45));
  INV_X1    g488(.A(new_n649), .ZN(new_n675));
  AND4_X1   g489(.A1(new_n316), .A2(new_n317), .A3(new_n620), .A4(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT94), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n488), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n594), .A2(new_n633), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n548), .A2(new_n550), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT32), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n679), .B1(new_n683), .B2(new_n538), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n316), .A2(new_n317), .A3(new_n620), .A4(new_n675), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT94), .B1(new_n685), .B2(new_n487), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n678), .A2(new_n684), .A3(new_n424), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  INV_X1    g502(.A(new_n598), .ZN(new_n689));
  INV_X1    g503(.A(new_n621), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n400), .A2(new_n413), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n227), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n319), .A3(new_n640), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n689), .A2(new_n690), .A3(new_n604), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  INV_X1    g512(.A(new_n625), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n604), .A3(new_n699), .A4(new_n695), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  NOR2_X1   g515(.A1(new_n694), .A2(new_n487), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n684), .A2(new_n494), .A3(new_n318), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  AOI21_X1  g518(.A(KEYINPUT95), .B1(new_n520), .B2(new_n522), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT95), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n519), .A2(new_n521), .A3(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n705), .A2(new_n707), .A3(new_n527), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n544), .A2(new_n547), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n550), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n548), .A2(new_n227), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT96), .B1(new_n711), .B2(G472), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT96), .ZN(new_n713));
  AOI211_X1 g527(.A(new_n713), .B(new_n601), .C1(new_n548), .C2(new_n227), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n597), .B(new_n710), .C1(new_n712), .C2(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n715), .A2(new_n493), .A3(new_n694), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT97), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n670), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n316), .A2(new_n232), .A3(new_n317), .A4(KEYINPUT97), .ZN(new_n719));
  AND4_X1   g533(.A1(KEYINPUT98), .A2(new_n718), .A3(new_n488), .A4(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n487), .B1(new_n670), .B2(new_n717), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT98), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n716), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT99), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT99), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n716), .B(new_n725), .C1(new_n720), .C2(new_n722), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  OAI211_X1 g542(.A(new_n634), .B(new_n710), .C1(new_n712), .C2(new_n714), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n488), .A2(new_n319), .A3(new_n640), .A4(new_n693), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n685), .B(KEYINPUT100), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT101), .B(G125), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G27));
  AOI21_X1  g549(.A(new_n410), .B1(new_n418), .B2(new_n409), .ZN(new_n736));
  INV_X1    g550(.A(new_n422), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT102), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n422), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(G469), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n320), .B1(new_n741), .B2(new_n415), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n485), .B1(new_n643), .B2(new_n644), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT103), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(KEYINPUT103), .B(new_n485), .C1(new_n643), .C2(new_n644), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT104), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n742), .A2(new_n745), .A3(new_n749), .A4(new_n746), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n689), .A3(new_n732), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n683), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n681), .A2(KEYINPUT105), .A3(new_n682), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n538), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n597), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n610), .A2(KEYINPUT100), .A3(new_n620), .A4(new_n675), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT100), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n685), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n748), .B2(new_n750), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n752), .A2(new_n753), .B1(new_n758), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n264), .ZN(G33));
  NAND3_X1  g579(.A1(new_n751), .A2(new_n689), .A3(new_n650), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT106), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n598), .B1(new_n748), .B2(new_n750), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT106), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n650), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND3_X1  g586(.A1(new_n738), .A2(KEYINPUT45), .A3(new_n740), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n420), .B2(new_n422), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n321), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n641), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n640), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT108), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n779), .B2(new_n641), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n781), .B2(KEYINPUT108), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n320), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n316), .A2(new_n317), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n620), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT43), .Z(new_n788));
  NOR2_X1   g602(.A1(new_n603), .A2(new_n679), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT44), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n745), .A2(new_n746), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n790), .B2(KEYINPUT44), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n785), .A2(new_n791), .A3(new_n666), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT109), .B(G137), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G39));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n785), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n785), .B1(new_n801), .B2(new_n799), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OR4_X1    g617(.A1(new_n553), .A2(new_n793), .A3(new_n597), .A4(new_n685), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n249), .ZN(G42));
  NOR2_X1   g620(.A1(G952), .A2(G953), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT117), .Z(new_n808));
  NAND2_X1  g622(.A1(new_n788), .A2(new_n490), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n715), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n792), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n693), .A2(new_n640), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(KEYINPUT113), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n320), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n812), .B1(new_n803), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n715), .A2(new_n669), .A3(new_n485), .A4(new_n694), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n810), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT50), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n793), .A2(new_n694), .ZN(new_n822));
  INV_X1    g636(.A(new_n665), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n597), .A4(new_n490), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT114), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n610), .A2(new_n620), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n809), .A2(new_n694), .A3(new_n793), .ZN(new_n828));
  INV_X1    g642(.A(new_n729), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n821), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  OR3_X1    g645(.A1(new_n817), .A2(new_n818), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n818), .B1(new_n817), .B2(new_n831), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n810), .A2(new_n702), .A3(new_n811), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT115), .Z(new_n835));
  AND2_X1   g649(.A1(new_n757), .A2(new_n597), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n489), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n835), .B(new_n841), .C1(new_n690), .C2(new_n825), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n832), .A2(new_n833), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n696), .A2(new_n700), .A3(new_n703), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n724), .B2(new_n726), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n752), .A2(new_n753), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n758), .A2(new_n763), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n786), .A2(new_n620), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n605), .A2(new_n318), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n495), .B1(new_n635), .B2(new_n598), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n751), .A2(new_n732), .A3(new_n829), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n232), .A2(new_n314), .A3(new_n649), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n684), .A2(new_n792), .A3(new_n424), .A4(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n846), .A2(new_n849), .A3(new_n771), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n711), .A2(G472), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n713), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n602), .A2(KEYINPUT96), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n634), .A3(new_n702), .A4(new_n710), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n651), .B1(new_n863), .B2(new_n762), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n424), .A2(new_n678), .A3(new_n684), .A4(new_n686), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n742), .A2(new_n679), .A3(new_n675), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n663), .B2(new_n664), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n720), .B2(new_n722), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT52), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n650), .A2(new_n488), .A3(new_n424), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n731), .A2(new_n732), .B1(new_n684), .B2(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(KEYINPUT52), .A2(new_n869), .A3(new_n872), .A4(new_n687), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT53), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n844), .B1(new_n858), .B2(new_n874), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n769), .A2(new_n751), .A3(new_n689), .A4(new_n650), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n769), .B1(new_n768), .B2(new_n650), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n878), .A2(new_n764), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  INV_X1    g696(.A(new_n869), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n733), .A2(new_n651), .A3(new_n687), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n866), .A2(KEYINPUT52), .A3(new_n869), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n880), .A2(new_n887), .A3(KEYINPUT111), .A4(new_n846), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n870), .A2(new_n873), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n881), .B1(new_n858), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n875), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT112), .B1(new_n858), .B2(new_n874), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT112), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n880), .A2(new_n887), .A3(new_n894), .A4(new_n846), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n897), .A3(new_n890), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n808), .B1(new_n843), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n813), .B(KEYINPUT49), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n320), .A2(new_n671), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n597), .A2(new_n786), .A3(new_n620), .A4(new_n902), .ZN(new_n903));
  OR3_X1    g717(.A1(new_n901), .A2(new_n903), .A3(new_n669), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n665), .B2(new_n904), .ZN(G75));
  NOR2_X1   g719(.A1(new_n241), .A2(G952), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n896), .A2(new_n890), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(G902), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(new_n483), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n445), .A2(new_n447), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT118), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT55), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT119), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(new_n456), .Z(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n907), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n911), .A2(new_n917), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n911), .A2(new_n921), .A3(new_n917), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(G51));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n898), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n896), .A2(KEYINPUT121), .A3(new_n897), .A4(new_n890), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n322), .B(KEYINPUT57), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n691), .B(KEYINPUT122), .Z(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n910), .A2(new_n779), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n906), .B1(new_n932), .B2(new_n933), .ZN(G54));
  INV_X1    g748(.A(KEYINPUT58), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n910), .A2(new_n935), .A3(new_n233), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n907), .B1(new_n936), .B2(new_n300), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n300), .B2(new_n936), .ZN(G60));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n892), .B2(new_n898), .ZN(new_n941));
  INV_X1    g755(.A(new_n616), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n907), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n616), .A2(new_n940), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n928), .B2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n896), .B2(new_n890), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n907), .B1(new_n948), .B2(new_n595), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n631), .B(new_n947), .C1(new_n896), .C2(new_n890), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(G66));
  NAND2_X1  g768(.A1(new_n846), .A2(new_n853), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n241), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT124), .Z(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n492), .B2(new_n448), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(G898), .ZN(new_n960));
  INV_X1    g774(.A(new_n241), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n913), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n959), .B(new_n962), .Z(G69));
  OR2_X1    g777(.A1(new_n673), .A2(new_n884), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n689), .A2(new_n667), .ZN(new_n966));
  NOR4_X1   g780(.A1(new_n966), .A2(new_n793), .A3(new_n318), .A4(new_n850), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n795), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n241), .B1(new_n970), .B2(new_n805), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n531), .A2(new_n533), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(new_n294), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n971), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n973), .B1(G900), .B2(new_n961), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n803), .A2(new_n804), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n785), .A2(new_n666), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n980), .B(new_n836), .C1(new_n722), .C2(new_n720), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n795), .A2(new_n866), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n878), .A2(new_n764), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT127), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n979), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n978), .B1(new_n985), .B2(new_n961), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n975), .A2(new_n977), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n241), .B1(G227), .B2(G900), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n988), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n975), .A2(new_n986), .A3(new_n990), .A4(new_n977), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  INV_X1    g808(.A(new_n970), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n979), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n996), .B2(new_n955), .ZN(new_n997));
  INV_X1    g811(.A(new_n655), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n906), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n891), .A2(new_n536), .A3(new_n655), .A4(new_n994), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n994), .B1(new_n985), .B2(new_n955), .ZN(new_n1001));
  INV_X1    g815(.A(new_n536), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .ZN(G57));
endmodule


