//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n198), .A2(G128), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(new_n199), .B2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n196), .A2(KEYINPUT65), .A3(G143), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .A4(new_n200), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(KEYINPUT68), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(KEYINPUT68), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n202), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT70), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n205), .A2(new_n200), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n204), .A4(new_n207), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n208), .A2(KEYINPUT68), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n201), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT70), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G134), .ZN(new_n221));
  INV_X1    g035(.A(G134), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G137), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n225), .B(G131), .C1(new_n224), .C2(new_n221), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT11), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n222), .B2(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n220), .A2(KEYINPUT11), .A3(G134), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n230), .A4(new_n223), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n213), .A2(new_n219), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(new_n229), .A3(new_n223), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n197), .A2(new_n200), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n239), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n204), .A2(new_n205), .A3(new_n200), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(new_n244), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n237), .B(new_n241), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G116), .B(G119), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT2), .B(G113), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n250), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n248), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT69), .ZN(new_n254));
  OR3_X1    g068(.A1(new_n252), .A2(KEYINPUT69), .A3(new_n248), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n247), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n247), .B1(new_n218), .B2(new_n232), .ZN(new_n259));
  INV_X1    g073(.A(new_n256), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n234), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n195), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n216), .A2(new_n217), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT70), .B1(new_n264), .B2(new_n202), .ZN(new_n265));
  AOI211_X1 g079(.A(new_n212), .B(new_n201), .C1(new_n216), .C2(new_n217), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n257), .B1(new_n267), .B2(new_n233), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n259), .A2(new_n260), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n234), .A2(new_n247), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n260), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n234), .A2(KEYINPUT73), .A3(new_n247), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT28), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(KEYINPUT74), .B(new_n194), .C1(new_n271), .C2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n234), .A2(KEYINPUT30), .A3(new_n247), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n279));
  NAND2_X1  g093(.A1(new_n259), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n260), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n268), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n193), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n281), .A2(KEYINPUT31), .A3(new_n193), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n234), .A2(KEYINPUT73), .A3(new_n247), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT73), .B1(new_n234), .B2(new_n247), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n289), .A2(new_n290), .A3(new_n260), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n263), .B(new_n270), .C1(new_n291), .C2(KEYINPUT28), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT74), .B1(new_n292), .B2(new_n194), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n187), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n187), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(new_n295), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n288), .B2(new_n293), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n193), .B1(new_n281), .B2(new_n282), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(KEYINPUT29), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(new_n292), .B2(new_n194), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n256), .B1(new_n234), .B2(new_n247), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n305), .B(KEYINPUT28), .C1(new_n306), .C2(new_n268), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT28), .B1(new_n306), .B2(new_n268), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT75), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n309), .B2(new_n276), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n193), .A2(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n304), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G472), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n194), .B1(new_n271), .B2(new_n276), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n287), .A3(new_n277), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT76), .A3(new_n298), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n296), .A2(new_n301), .A3(new_n315), .A4(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n211), .A2(G125), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G953), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G224), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n325), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT80), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G104), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G107), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G107), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G104), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(G104), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n330), .ZN(new_n340));
  INV_X1    g154(.A(G101), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(G101), .B1(new_n335), .B2(new_n338), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n248), .A2(KEYINPUT5), .ZN(new_n346));
  INV_X1    g160(.A(G116), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n347), .A2(KEYINPUT5), .A3(G119), .ZN(new_n348));
  INV_X1    g162(.A(G113), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n346), .A2(new_n350), .B1(new_n252), .B2(new_n248), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n339), .A2(new_n330), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n334), .A2(G107), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n353), .B(new_n354), .C1(new_n355), .C2(new_n339), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G101), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n342), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT81), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n354), .B1(new_n335), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n339), .B1(new_n330), .B2(new_n332), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n364), .B2(new_n341), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n357), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n356), .A2(new_n360), .A3(G101), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n254), .A2(new_n369), .A3(new_n255), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n352), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G122), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n370), .B1(new_n359), .B2(new_n367), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(new_n352), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(KEYINPUT6), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(new_n375), .C1(new_n376), .C2(new_n352), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n380), .A2(new_n381), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n328), .B(new_n378), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n373), .B(KEYINPUT8), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n345), .A2(new_n351), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n352), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT7), .ZN(new_n388));
  AOI22_X1  g202(.A1(KEYINPUT86), .A2(new_n388), .B1(new_n326), .B2(G224), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(KEYINPUT86), .B2(new_n388), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n323), .B2(new_n324), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n372), .B2(new_n373), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n325), .A2(KEYINPUT7), .A3(new_n327), .ZN(new_n394));
  AOI21_X1  g208(.A(G902), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n384), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G210), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n384), .A2(new_n395), .A3(new_n397), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G214), .B1(G237), .B2(G902), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G478), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT15), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT92), .B1(new_n347), .B2(G122), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n408));
  INV_X1    g222(.A(G122), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(G116), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n347), .A2(G122), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G107), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n337), .A3(new_n412), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(KEYINPUT93), .A3(new_n415), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT13), .B1(new_n206), .B2(G143), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(new_n222), .ZN(new_n421));
  XNOR2_X1  g235(.A(G128), .B(G143), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n412), .B(KEYINPUT14), .ZN(new_n425));
  INV_X1    g239(.A(new_n411), .ZN(new_n426));
  OAI21_X1  g240(.A(G107), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n422), .B(new_n222), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n415), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT9), .B(G234), .ZN(new_n430));
  INV_X1    g244(.A(G217), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n430), .A2(new_n431), .A3(G953), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n424), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n424), .B2(new_n429), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n313), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT94), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(KEYINPUT94), .B(new_n313), .C1(new_n434), .C2(new_n435), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n406), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n435), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n433), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT94), .B1(new_n442), .B2(new_n313), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n405), .ZN(new_n444));
  AOI211_X1 g258(.A(new_n313), .B(new_n326), .C1(G234), .C2(G237), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(G898), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g261(.A1(KEYINPUT95), .A2(G952), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT95), .A2(G952), .ZN(new_n449));
  AOI21_X1  g263(.A(G953), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G234), .ZN(new_n451));
  INV_X1    g265(.A(G237), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n440), .A2(new_n444), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n326), .A3(G214), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n199), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT18), .A3(G131), .ZN(new_n461));
  XNOR2_X1  g275(.A(G125), .B(G140), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n196), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT18), .A2(G131), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n458), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G140), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT16), .ZN(new_n469));
  INV_X1    g283(.A(G125), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G140), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n471), .A3(KEYINPUT16), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT77), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n468), .A2(KEYINPUT77), .A3(KEYINPUT16), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n474), .A2(new_n196), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT88), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n462), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT19), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n462), .A2(new_n477), .A3(KEYINPUT19), .ZN(new_n481));
  AOI21_X1  g295(.A(G146), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n460), .B2(G131), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n460), .A2(G131), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n458), .A2(KEYINPUT87), .A3(new_n230), .A4(new_n459), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n466), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n334), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n456), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n493));
  INV_X1    g307(.A(new_n475), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT77), .B1(new_n462), .B2(KEYINPUT16), .ZN(new_n495));
  OAI211_X1 g309(.A(G146), .B(new_n494), .C1(new_n495), .C2(new_n469), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n480), .A2(new_n481), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(G146), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n491), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(KEYINPUT89), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n488), .A2(KEYINPUT17), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n196), .B1(new_n474), .B2(new_n475), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n496), .C1(new_n505), .C2(new_n486), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n491), .B(new_n493), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n492), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(G475), .A2(G902), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n508), .A2(KEYINPUT90), .A3(new_n509), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(KEYINPUT20), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT90), .B1(new_n508), .B2(new_n509), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n493), .B1(new_n503), .B2(new_n506), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT91), .A3(new_n501), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n517), .A2(new_n501), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n507), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n313), .B(new_n518), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n515), .A2(new_n516), .B1(new_n522), .B2(G475), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n455), .A2(KEYINPUT96), .A3(new_n514), .A4(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT96), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n514), .A2(new_n523), .ZN(new_n526));
  INV_X1    g340(.A(new_n439), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n405), .B1(new_n443), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n454), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n438), .A2(new_n406), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n525), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n403), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n431), .B1(G234), .B2(new_n313), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n206), .A2(G119), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT23), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n539));
  INV_X1    g353(.A(G110), .ZN(new_n540));
  INV_X1    g354(.A(G119), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G128), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n536), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT24), .B(G110), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n543), .A2(new_n546), .B1(new_n196), .B2(new_n462), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n496), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT22), .B(G137), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n326), .A2(G221), .A3(G234), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n549), .A2(G221), .A3(G234), .A4(new_n326), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n504), .A2(new_n496), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n538), .A2(new_n542), .A3(new_n539), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G110), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n544), .A2(new_n545), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n548), .B(new_n554), .C1(new_n555), .C2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n553), .B(KEYINPUT78), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n504), .B2(new_n496), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n496), .A2(new_n547), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(new_n564), .A3(new_n313), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT25), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n560), .A2(new_n564), .A3(KEYINPUT25), .A4(new_n313), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n535), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n560), .A2(new_n564), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n534), .A2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT79), .ZN(new_n576));
  INV_X1    g390(.A(G469), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n313), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G140), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n326), .A2(G227), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n237), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n344), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n369), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n322), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n267), .A2(new_n584), .B1(new_n368), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n216), .A2(KEYINPUT82), .A3(new_n217), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n214), .A2(new_n204), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n198), .A2(G128), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT82), .B1(new_n216), .B2(new_n217), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n345), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n583), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n582), .B1(new_n587), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n366), .B1(new_n365), .B2(new_n357), .ZN(new_n597));
  AND4_X1   g411(.A1(new_n366), .A2(new_n357), .A3(KEYINPUT4), .A4(new_n342), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n586), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n213), .A2(new_n219), .A3(new_n584), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n595), .A2(new_n582), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n581), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n581), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n218), .A2(new_n344), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n594), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT12), .B1(new_n606), .B2(new_n237), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n608), .B(new_n582), .C1(new_n594), .C2(new_n605), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n601), .B(new_n604), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n603), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n578), .B1(new_n611), .B2(new_n577), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n601), .B1(new_n607), .B2(new_n609), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(KEYINPUT83), .B(new_n601), .C1(new_n607), .C2(new_n609), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n581), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n601), .A2(new_n604), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT84), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n595), .A2(new_n599), .A3(new_n600), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n237), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT84), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n601), .A2(new_n622), .A3(new_n604), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n617), .A2(G469), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n576), .B1(new_n612), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n321), .A2(new_n533), .A3(new_n574), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT97), .B(G101), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G3));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n433), .B2(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n442), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n441), .B(new_n433), .C1(KEYINPUT99), .C2(new_n630), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n404), .A2(G902), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT100), .B(G478), .Z(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n634), .A2(new_n635), .B1(new_n436), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n526), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n403), .A2(new_n454), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n626), .A2(new_n294), .A3(new_n574), .ZN(new_n642));
  INV_X1    g456(.A(G472), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n313), .B1(new_n288), .B2(new_n293), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n319), .A2(KEYINPUT98), .A3(new_n313), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n641), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT34), .B(G104), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  AND2_X1   g465(.A1(new_n642), .A2(new_n648), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n440), .A2(new_n444), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n514), .A3(new_n523), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n403), .A2(new_n655), .A3(new_n454), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NAND2_X1  g475(.A1(new_n524), .A2(new_n532), .ZN(new_n662));
  INV_X1    g476(.A(new_n402), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n399), .B2(new_n400), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n567), .A2(new_n568), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n534), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n561), .A2(KEYINPUT36), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n562), .A2(new_n563), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n667), .B(new_n668), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n571), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n666), .A2(KEYINPUT103), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n667), .B(new_n668), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n572), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n672), .B1(new_n569), .B2(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n671), .A2(KEYINPUT104), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT104), .B1(new_n671), .B2(new_n675), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n626), .A2(new_n662), .A3(new_n664), .A4(new_n678), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n646), .A2(new_n647), .B1(new_n187), .B2(new_n319), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  AND4_X1   g497(.A1(new_n296), .A2(new_n301), .A3(new_n315), .A4(new_n320), .ZN(new_n684));
  INV_X1    g498(.A(new_n445), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n453), .B1(new_n685), .B2(G900), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT105), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n526), .A2(new_n653), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n626), .A2(new_n678), .A3(new_n664), .A4(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n626), .A2(new_n678), .A3(new_n664), .A4(new_n688), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(new_n321), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  INV_X1    g509(.A(new_n400), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n397), .B1(new_n384), .B2(new_n395), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT38), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT38), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n401), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n671), .A2(new_n675), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n654), .A2(new_n402), .A3(new_n526), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n687), .B(KEYINPUT39), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n626), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n194), .B1(new_n306), .B2(new_n268), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n283), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n313), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G472), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n296), .A2(new_n301), .A3(new_n320), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n705), .A2(new_n708), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  AND2_X1   g530(.A1(new_n626), .A2(new_n678), .ZN(new_n717));
  INV_X1    g531(.A(new_n687), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n526), .A2(new_n639), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n321), .A2(new_n717), .A3(new_n664), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT107), .B(G146), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G48));
  NAND2_X1  g536(.A1(new_n603), .A2(new_n610), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n313), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  INV_X1    g539(.A(new_n610), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n604), .B1(new_n621), .B2(new_n601), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n577), .B(new_n313), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n728), .A3(new_n575), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n321), .A2(new_n641), .A3(new_n574), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  NAND4_X1  g547(.A1(new_n321), .A2(new_n656), .A3(new_n574), .A4(new_n730), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  NOR2_X1   g549(.A1(new_n403), .A2(new_n729), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n321), .A2(new_n662), .A3(new_n678), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  OR2_X1    g552(.A1(new_n310), .A2(new_n193), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n297), .B1(new_n739), .B2(new_n287), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(G472), .B2(new_n644), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n704), .A2(new_n698), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n729), .A2(new_n454), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n741), .A2(new_n574), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  NAND4_X1  g559(.A1(new_n741), .A2(new_n736), .A3(new_n703), .A4(new_n719), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  INV_X1    g561(.A(new_n575), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n612), .B2(new_n625), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n696), .A2(new_n697), .A3(new_n663), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n321), .A2(new_n574), .A3(new_n719), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n574), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n294), .A2(new_n295), .B1(new_n314), .B2(G472), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(new_n299), .ZN(new_n757));
  AND4_X1   g571(.A1(KEYINPUT42), .A2(new_n749), .A3(new_n719), .A4(new_n750), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(KEYINPUT108), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT108), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n754), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND4_X1  g576(.A1(new_n321), .A2(new_n574), .A3(new_n688), .A4(new_n751), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n526), .A2(new_n638), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT43), .B1(new_n526), .B2(new_n638), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n703), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n648), .B2(new_n294), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n765), .B1(new_n771), .B2(KEYINPUT44), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n680), .A2(KEYINPUT109), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n578), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n623), .A2(new_n621), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n777), .A2(new_n616), .B1(new_n778), .B2(new_n619), .ZN(new_n779));
  OAI21_X1  g593(.A(G469), .B1(new_n779), .B2(KEYINPUT45), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n617), .A2(KEYINPUT45), .A3(new_n624), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n776), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n617), .A2(new_n624), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(G469), .A3(new_n781), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n728), .A2(new_n789), .A3(new_n776), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n748), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n784), .A2(new_n706), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n750), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(KEYINPUT44), .B2(new_n771), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n775), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT110), .B(G137), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(G39));
  NAND3_X1  g612(.A1(new_n750), .A2(new_n719), .A3(new_n755), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n321), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n790), .B1(new_n780), .B2(new_n782), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n575), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n789), .B1(new_n788), .B2(new_n776), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT47), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT47), .B1(new_n784), .B2(new_n791), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  NAND4_X1  g622(.A1(new_n731), .A2(new_n734), .A3(new_n737), .A4(new_n744), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n654), .A2(new_n526), .A3(new_n687), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n321), .A2(new_n717), .A3(new_n750), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n751), .A2(new_n741), .A3(new_n703), .A4(new_n719), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n763), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n761), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n627), .A2(new_n649), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT111), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT111), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n627), .A2(new_n818), .A3(new_n649), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n652), .A2(new_n656), .B1(new_n679), .B2(new_n680), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n746), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n690), .B2(new_n693), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n569), .A2(new_n674), .A3(new_n687), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n713), .A2(new_n742), .A3(new_n749), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n824), .A2(new_n825), .A3(new_n720), .A4(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n691), .A2(new_n321), .A3(new_n692), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n692), .B1(new_n691), .B2(new_n321), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n746), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n720), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT52), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n822), .A2(new_n834), .A3(KEYINPUT53), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n820), .A2(new_n819), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n814), .A3(new_n761), .A4(new_n817), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n828), .A2(new_n833), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT54), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n702), .A2(new_n663), .A3(new_n730), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT112), .ZN(new_n844));
  INV_X1    g658(.A(new_n453), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n768), .A2(new_n845), .A3(new_n769), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n846), .A2(new_n574), .A3(new_n741), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n844), .B(new_n847), .C1(KEYINPUT113), .C2(KEYINPUT50), .ZN(new_n848));
  AND2_X1   g662(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n804), .B1(new_n802), .B2(new_n803), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n791), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n725), .A2(new_n728), .ZN(new_n854));
  INV_X1    g668(.A(new_n576), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n847), .B(new_n750), .C1(new_n853), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n848), .A2(new_n849), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n793), .A2(new_n729), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n574), .A3(new_n845), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n713), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n526), .A2(new_n639), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n846), .A2(new_n859), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n741), .A2(new_n703), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n861), .A2(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n850), .A2(new_n857), .A3(new_n858), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  INV_X1    g684(.A(new_n861), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n450), .B1(new_n871), .B2(new_n640), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n864), .A2(new_n757), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT48), .Z(new_n874));
  AOI211_X1 g688(.A(new_n872), .B(new_n874), .C1(new_n736), .C2(new_n847), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n842), .A2(new_n869), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(G952), .A2(G953), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n854), .A2(KEYINPUT49), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n766), .A2(new_n574), .A3(new_n855), .A4(new_n402), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n881), .B(new_n702), .C1(KEYINPUT49), .C2(new_n854), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n877), .A2(new_n878), .B1(new_n713), .B2(new_n882), .ZN(G75));
  NAND3_X1  g697(.A1(new_n841), .A2(G210), .A3(G902), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n328), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n888), .B1(new_n884), .B2(new_n885), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n326), .A2(G952), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(G51));
  XNOR2_X1  g706(.A(new_n578), .B(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n842), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n723), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n788), .B(KEYINPUT114), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n841), .A2(G902), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n891), .B1(new_n895), .B2(new_n897), .ZN(G54));
  INV_X1    g712(.A(new_n508), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n841), .A2(G902), .ZN(new_n900));
  NAND2_X1  g714(.A1(KEYINPUT58), .A2(G475), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT115), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n891), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n900), .A2(new_n899), .A3(new_n902), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(G60));
  NAND2_X1  g721(.A1(G478), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT59), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n842), .A2(new_n634), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n634), .B1(new_n842), .B2(new_n909), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n910), .A2(new_n911), .A3(new_n891), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n841), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n570), .B(KEYINPUT118), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n891), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n835), .B2(new_n840), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n673), .B(KEYINPUT116), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n917), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n904), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n841), .A2(new_n915), .A3(new_n921), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT119), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n925), .B2(KEYINPUT117), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n930), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n927), .A3(new_n923), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(G66));
  INV_X1    g748(.A(G224), .ZN(new_n935));
  OAI21_X1  g749(.A(G953), .B1(new_n446), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n821), .A2(new_n809), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n886), .B1(G898), .B2(new_n326), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  NAND2_X1  g754(.A1(new_n278), .A2(new_n280), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n497), .B(KEYINPUT120), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n296), .A2(new_n315), .A3(new_n299), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n944), .A2(new_n574), .A3(new_n742), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n802), .A2(new_n803), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n706), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n944), .A2(new_n574), .A3(new_n742), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT123), .B1(new_n792), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n720), .A3(new_n824), .ZN(new_n952));
  AND4_X1   g766(.A1(new_n321), .A2(new_n574), .A3(new_n688), .A4(new_n751), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n853), .B2(new_n800), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n761), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n796), .ZN(new_n957));
  AOI21_X1  g771(.A(G953), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n326), .A2(G900), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT122), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n943), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT121), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n720), .B(new_n746), .C1(new_n829), .C2(new_n830), .ZN(new_n965));
  INV_X1    g779(.A(new_n715), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n824), .A2(KEYINPUT62), .A3(new_n715), .A4(new_n720), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n793), .B(new_n707), .C1(new_n640), .C2(new_n655), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n684), .A2(new_n755), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n807), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n774), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n771), .A2(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n771), .A2(KEYINPUT44), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n978), .A2(new_n793), .A3(new_n792), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n973), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(G953), .B1(new_n969), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n963), .B1(new_n981), .B2(new_n943), .ZN(new_n982));
  INV_X1    g796(.A(new_n943), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n853), .A2(new_n800), .B1(new_n970), .B2(new_n971), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n775), .B2(new_n795), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n967), .B2(new_n968), .ZN(new_n986));
  OAI211_X1 g800(.A(KEYINPUT121), .B(new_n983), .C1(new_n986), .C2(G953), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n326), .B1(G227), .B2(G900), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n962), .A2(new_n982), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  INV_X1    g805(.A(new_n965), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(new_n761), .A3(new_n954), .A4(new_n951), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n326), .B1(new_n993), .B2(new_n796), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n983), .B1(new_n994), .B2(new_n960), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(new_n988), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT124), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n996), .A2(new_n997), .A3(new_n982), .A4(new_n987), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n991), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n981), .A2(new_n943), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n988), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT125), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n999), .A2(KEYINPUT125), .A3(new_n1001), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  XNOR2_X1  g820(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n643), .A2(new_n313), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n283), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n841), .B(new_n1009), .C1(new_n1010), .C2(new_n302), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n986), .A2(new_n937), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n1009), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n281), .A2(new_n282), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT127), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1013), .A2(new_n193), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n956), .A2(new_n957), .A3(new_n937), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n1009), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1015), .A2(new_n193), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n891), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1011), .A2(new_n1016), .A3(new_n1020), .ZN(G57));
endmodule


