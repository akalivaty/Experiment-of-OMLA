//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n191), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G125), .B(G140), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n199), .B1(new_n201), .B2(KEYINPUT16), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT72), .B1(new_n206), .B2(G128), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G110), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT24), .B(G110), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT71), .B1(new_n206), .B2(G128), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT71), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G119), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n212), .B(new_n215), .C1(G119), .C2(new_n214), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n204), .B(new_n210), .C1(new_n211), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n211), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n209), .B2(G110), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT65), .B(G146), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n202), .A2(G146), .B1(new_n201), .B2(new_n220), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n219), .A2(KEYINPUT73), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT73), .B1(new_n219), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n217), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G137), .ZN(new_n225));
  INV_X1    g039(.A(G221), .ZN(new_n226));
  INV_X1    g040(.A(G234), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n226), .A2(new_n227), .A3(G953), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n225), .B(new_n228), .Z(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n217), .B(new_n229), .C1(new_n222), .C2(new_n223), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n188), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n232), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n190), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n189), .A2(G902), .ZN(new_n238));
  XOR2_X1   g052(.A(new_n238), .B(KEYINPUT75), .Z(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n231), .A2(new_n232), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT74), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n237), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G472), .ZN(new_n246));
  NOR2_X1   g060(.A1(G237), .A2(G953), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G210), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n248), .B(KEYINPUT27), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G101), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT70), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G119), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n206), .A2(G116), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT68), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT2), .B(G113), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n206), .A2(G116), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(G119), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT2), .B(G113), .Z(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n260), .A3(new_n261), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n191), .A2(KEYINPUT65), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n271), .A3(G143), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n273));
  INV_X1    g087(.A(G143), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(G146), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT66), .B1(new_n191), .B2(G143), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n272), .A2(new_n275), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n214), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n274), .A2(G146), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n269), .A2(new_n271), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(new_n274), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n278), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT67), .B1(new_n284), .B2(G137), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n286));
  INV_X1    g100(.A(G137), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G134), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(G137), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G131), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT11), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n284), .B2(G137), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n287), .A2(KEYINPUT11), .A3(G134), .ZN(new_n294));
  INV_X1    g108(.A(G131), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .A4(new_n289), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n293), .A2(new_n294), .A3(new_n289), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G131), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n296), .ZN(new_n301));
  AND2_X1   g115(.A1(KEYINPUT0), .A2(G128), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n272), .A2(new_n275), .A3(new_n276), .A4(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n305));
  NOR2_X1   g119(.A1(KEYINPUT0), .A2(G128), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(G143), .B1(new_n269), .B2(new_n271), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n280), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n301), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n268), .B1(new_n298), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n298), .A2(new_n268), .A3(new_n310), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n254), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n254), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n253), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n291), .A2(new_n296), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n220), .B2(G143), .ZN(new_n321));
  OAI22_X1  g135(.A1(new_n321), .A2(new_n214), .B1(new_n280), .B2(new_n308), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n319), .B1(new_n322), .B2(new_n278), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n301), .A2(new_n303), .A3(new_n309), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n318), .B(KEYINPUT30), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT30), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT69), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n318), .A2(KEYINPUT30), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n298), .A2(new_n310), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n268), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n251), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n298), .A2(new_n268), .A3(new_n310), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n317), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g149(.A(KEYINPUT69), .B(new_n326), .C1(new_n298), .C2(new_n310), .ZN(new_n336));
  AND4_X1   g150(.A1(new_n298), .A2(new_n310), .A3(new_n327), .A4(new_n328), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n267), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n251), .A3(new_n313), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(KEYINPUT31), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n246), .B(new_n188), .C1(new_n335), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT32), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT28), .B1(new_n332), .B2(new_n311), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n252), .B1(new_n343), .B2(new_n315), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n339), .B2(KEYINPUT31), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n325), .A2(new_n329), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n332), .B1(new_n346), .B2(new_n267), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n334), .A3(new_n251), .ZN(new_n348));
  AOI21_X1  g162(.A(G902), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n246), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n342), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n314), .A2(new_n316), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n252), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n251), .B2(new_n347), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n354), .B1(new_n353), .B2(new_n251), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n188), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G472), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n245), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT19), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT19), .B1(new_n193), .B2(new_n195), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n220), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G237), .ZN(new_n364));
  INV_X1    g178(.A(G953), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G214), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT84), .A3(new_n274), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n274), .A2(KEYINPUT84), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G214), .A3(new_n247), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n295), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n295), .B1(new_n367), .B2(new_n369), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n203), .B(new_n363), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT18), .A3(G131), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n196), .A2(G146), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n196), .B2(new_n281), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n367), .A2(new_n378), .A3(new_n369), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT17), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n374), .A2(KEYINPUT17), .A3(G131), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n200), .A3(new_n203), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n384), .B(new_n380), .C1(new_n387), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n392));
  NOR2_X1   g206(.A1(G475), .A2(G902), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n395));
  INV_X1    g209(.A(new_n393), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n386), .B2(new_n390), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n365), .A2(G952), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n227), .B2(new_n364), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n188), .B(new_n365), .C1(G234), .C2(G237), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT21), .B(G898), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n372), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT17), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n370), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n408), .A2(new_n203), .A3(new_n200), .A4(new_n388), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n384), .B1(new_n409), .B2(new_n380), .ZN(new_n410));
  INV_X1    g224(.A(new_n390), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n188), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G475), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n398), .A2(new_n405), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n415));
  INV_X1    g229(.A(G107), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT85), .B(G122), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G116), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n416), .B1(new_n418), .B2(KEYINPUT14), .ZN(new_n419));
  INV_X1    g233(.A(G122), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(G116), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n214), .A2(G143), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n214), .A3(G143), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT86), .B1(new_n274), .B2(G128), .ZN(new_n428));
  AOI211_X1 g242(.A(new_n424), .B(new_n425), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n427), .ZN(new_n430));
  INV_X1    g244(.A(new_n425), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT88), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n429), .A2(new_n432), .A3(new_n284), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n426), .B1(new_n214), .B2(G143), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n274), .A2(KEYINPUT86), .A3(G128), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n424), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n430), .A2(KEYINPUT88), .A3(new_n431), .ZN(new_n438));
  AOI21_X1  g252(.A(G134), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n423), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n284), .B1(new_n429), .B2(new_n432), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(G134), .A3(new_n438), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT89), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n422), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n421), .B(G107), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n425), .A2(KEYINPUT13), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT87), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n430), .B1(KEYINPUT13), .B2(new_n425), .ZN(new_n448));
  OAI21_X1  g262(.A(G134), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n445), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(new_n187), .A3(G953), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n444), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n422), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT89), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT89), .B1(new_n441), .B2(new_n442), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n445), .A2(new_n441), .A3(new_n449), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n415), .B(new_n188), .C1(new_n454), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(KEYINPUT15), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n453), .B1(new_n444), .B2(new_n450), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(new_n459), .A3(new_n452), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n463), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n415), .A3(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n414), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G140), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n365), .A2(G227), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT10), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT76), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT3), .B1(new_n383), .B2(G107), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n416), .A3(G104), .ZN(new_n479));
  INV_X1    g293(.A(G101), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n383), .A2(G107), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n477), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n383), .A2(G107), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n416), .A2(G104), .ZN(new_n484));
  OAI21_X1  g298(.A(G101), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT1), .B1(new_n274), .B2(G146), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G128), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n269), .A2(new_n271), .A3(G143), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n276), .A2(new_n275), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n476), .B(new_n486), .C1(new_n278), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n278), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n482), .A2(new_n485), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT76), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n475), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n301), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(G101), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n309), .A2(new_n303), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(G101), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(KEYINPUT4), .A3(new_n482), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n486), .A2(new_n475), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n501), .A2(new_n503), .B1(new_n283), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n496), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n486), .B(new_n278), .C1(new_n279), .C2(new_n282), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n276), .A2(new_n275), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n509), .A2(new_n272), .B1(G128), .B2(new_n487), .ZN(new_n510));
  AND4_X1   g324(.A1(new_n272), .A2(new_n275), .A3(new_n276), .A4(new_n277), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n494), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n476), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n493), .A2(KEYINPUT76), .A3(new_n494), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT77), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT12), .B1(new_n301), .B2(new_n516), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n515), .A2(new_n497), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n507), .B1(new_n492), .B2(new_n495), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n520), .B2(new_n301), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n474), .B(new_n506), .C1(new_n518), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT10), .B1(new_n513), .B2(new_n514), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n501), .A2(new_n503), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n283), .A2(new_n504), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n523), .A2(new_n526), .A3(new_n301), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n497), .B1(new_n496), .B2(new_n505), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n473), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G469), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n188), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n527), .A2(new_n473), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n301), .B1(new_n523), .B2(new_n526), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n520), .A2(new_n301), .A3(new_n519), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n517), .B1(new_n515), .B2(new_n497), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n527), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n535), .B(G469), .C1(new_n538), .C2(new_n474), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n531), .A2(new_n188), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n532), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n451), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n226), .B1(new_n543), .B2(new_n188), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G214), .B1(G237), .B2(G902), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n267), .A2(new_n503), .A3(new_n500), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT5), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n258), .B2(new_n263), .ZN(new_n550));
  OAI21_X1  g364(.A(G113), .B1(new_n260), .B2(KEYINPUT5), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n494), .B(new_n266), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT6), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n548), .A2(new_n552), .A3(new_n555), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT6), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n555), .B1(new_n548), .B2(new_n552), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT78), .B(new_n557), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n560), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT78), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT6), .A4(new_n558), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n194), .B1(new_n309), .B2(new_n303), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n566), .A2(KEYINPUT79), .B1(new_n283), .B2(G125), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT79), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n568), .B(new_n194), .C1(new_n309), .C2(new_n303), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n365), .A2(G224), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT80), .Z(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n309), .A2(new_n303), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n568), .B1(new_n574), .B2(new_n194), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n566), .A2(KEYINPUT79), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n322), .A2(new_n194), .A3(new_n278), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n572), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n565), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n266), .B(new_n486), .C1(new_n550), .C2(new_n551), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n256), .A2(new_n257), .A3(new_n549), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n266), .B1(new_n584), .B2(new_n551), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n494), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n555), .B(KEYINPUT8), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n558), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT81), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n571), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n571), .A2(KEYINPUT7), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n591), .B(new_n592), .C1(new_n567), .C2(new_n569), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT7), .B(new_n571), .C1(new_n570), .C2(new_n590), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G210), .B1(G237), .B2(G902), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT82), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n582), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n599), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n561), .A2(new_n564), .B1(new_n573), .B2(new_n580), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n589), .A2(new_n593), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n592), .B1(new_n578), .B2(new_n591), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n188), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n601), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n547), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n470), .A2(new_n542), .A3(new_n545), .A4(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n360), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  AOI211_X1 g425(.A(G472), .B(G902), .C1(new_n345), .C2(new_n348), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n339), .A2(KEYINPUT31), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n348), .A3(new_n317), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n246), .B1(new_n614), .B2(new_n188), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n522), .B2(new_n529), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n540), .B1(new_n617), .B2(new_n531), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n544), .B1(new_n618), .B2(new_n539), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n619), .A3(new_n244), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT91), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n582), .A2(new_n596), .A3(new_n598), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n597), .B1(new_n602), .B2(new_n605), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n546), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT92), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n622), .A2(new_n623), .A3(KEYINPUT92), .A4(new_n546), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n465), .A2(new_n466), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n465), .A2(KEYINPUT93), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n630), .A3(KEYINPUT33), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n465), .B(new_n466), .C1(KEYINPUT93), .C2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(G478), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n462), .A2(new_n188), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n467), .B2(new_n462), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n398), .A2(new_n413), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n405), .A3(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n621), .A2(new_n628), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT34), .B(G104), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  INV_X1    g456(.A(new_n628), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n464), .A2(new_n469), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n397), .A2(new_n395), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n397), .A2(new_n395), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n413), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n645), .A2(new_n404), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n621), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT35), .B(G107), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  AND2_X1   g468(.A1(new_n470), .A2(new_n607), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n224), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n224), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n657), .A2(new_n240), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n237), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n655), .A2(new_n619), .A3(new_n616), .A4(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  AOI21_X1  g478(.A(new_n660), .B1(new_n352), .B2(new_n359), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n626), .A2(new_n545), .A3(new_n542), .A4(new_n627), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n402), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n400), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n645), .A2(new_n648), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n665), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  INV_X1    g488(.A(new_n600), .ZN(new_n675));
  INV_X1    g489(.A(new_n606), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT38), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n638), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n464), .B2(new_n469), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n546), .A2(new_n679), .A3(new_n660), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n312), .A2(new_n313), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n333), .B1(new_n683), .B2(new_n253), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n684), .A2(G902), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n352), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n542), .A2(new_n545), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n670), .B(KEYINPUT39), .Z(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT40), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT40), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n682), .A2(new_n687), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND4_X1  g509(.A1(new_n634), .A2(new_n638), .A3(new_n636), .A4(new_n670), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT94), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n665), .A2(new_n697), .A3(new_n667), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NOR2_X1   g513(.A1(new_n639), .A2(new_n628), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n537), .A2(new_n536), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n534), .A2(new_n506), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n533), .A2(new_n701), .B1(new_n702), .B2(new_n473), .ZN(new_n703));
  OAI21_X1  g517(.A(G469), .B1(new_n703), .B2(G902), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n545), .A3(new_n532), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n700), .A2(new_n360), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND3_X1  g523(.A1(new_n650), .A2(new_n360), .A3(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NAND2_X1  g525(.A1(new_n582), .A2(new_n596), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n547), .B1(new_n712), .B2(new_n597), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT92), .B1(new_n713), .B2(new_n622), .ZN(new_n714));
  INV_X1    g528(.A(new_n627), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n714), .A2(new_n715), .A3(new_n705), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n665), .A2(new_n470), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  INV_X1    g532(.A(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n341), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n614), .A2(new_n188), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G472), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n349), .A2(KEYINPUT95), .A3(new_n246), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n244), .A2(new_n720), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n626), .A2(new_n627), .A3(new_n681), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n724), .A2(new_n726), .A3(new_n405), .A4(new_n706), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  AND4_X1   g542(.A1(new_n722), .A2(new_n720), .A3(new_n661), .A4(new_n723), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n697), .A2(new_n729), .A3(new_n716), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n600), .A2(new_n606), .A3(new_n546), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n542), .A2(new_n733), .A3(new_n545), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT96), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n352), .A2(new_n359), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n619), .A2(KEYINPUT96), .A3(new_n733), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n244), .ZN(new_n739));
  INV_X1    g553(.A(new_n697), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n732), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n736), .A2(new_n738), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT42), .A3(new_n360), .A4(new_n697), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT97), .B(G131), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G33));
  NAND4_X1  g560(.A1(new_n360), .A2(new_n672), .A3(new_n736), .A4(new_n738), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  NAND2_X1  g562(.A1(new_n637), .A2(new_n680), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(KEYINPUT43), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(KEYINPUT43), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n722), .A2(new_n341), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n661), .ZN(new_n755));
  OR3_X1    g569(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n753), .B1(new_n752), .B2(new_n755), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n733), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(KEYINPUT98), .A3(new_n733), .A4(new_n757), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n535), .B1(new_n474), .B2(new_n538), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n531), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n541), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n532), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n545), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n689), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n760), .A2(new_n761), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n771), .A2(new_n775), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n342), .A2(new_n351), .B1(new_n358), .B2(G472), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n697), .A2(new_n245), .A3(new_n778), .A4(new_n733), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n776), .A2(new_n777), .B1(KEYINPUT99), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n780), .A2(KEYINPUT99), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  NAND4_X1  g598(.A1(new_n710), .A2(new_n707), .A3(new_n717), .A4(new_n727), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT103), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n547), .B(new_n404), .C1(new_n600), .C2(new_n606), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT102), .B1(new_n644), .B2(new_n680), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT102), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n789), .B(new_n638), .C1(new_n464), .C2(new_n469), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n620), .A2(new_n791), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n608), .A2(new_n754), .A3(new_n660), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n786), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n607), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n639), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n542), .A2(new_n244), .A3(new_n545), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n754), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n609), .A2(new_n360), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n662), .B(KEYINPUT103), .C1(new_n620), .C2(new_n791), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n794), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT104), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT104), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n794), .A2(new_n799), .A3(new_n803), .A4(new_n800), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n785), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT108), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n673), .A2(new_n730), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n778), .A2(new_n666), .A3(new_n660), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n670), .B(KEYINPUT107), .Z(new_n809));
  NAND4_X1  g623(.A1(new_n542), .A2(new_n545), .A3(new_n660), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n725), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n808), .A2(new_n697), .B1(new_n687), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n806), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n687), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n698), .A2(new_n673), .A3(new_n730), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(KEYINPUT108), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT52), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n807), .A2(new_n812), .A3(new_n806), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(KEYINPUT108), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n697), .A2(new_n729), .A3(new_n736), .A4(new_n738), .ZN(new_n822));
  INV_X1    g636(.A(new_n734), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n644), .A2(new_n648), .A3(new_n671), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n665), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n747), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT105), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT105), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n747), .A2(new_n822), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n827), .A2(new_n744), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n805), .A2(new_n817), .A3(new_n821), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n802), .A2(new_n804), .ZN(new_n837));
  INV_X1    g651(.A(new_n785), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n830), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n807), .A2(KEYINPUT106), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n673), .A2(new_n730), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT106), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n840), .A2(new_n698), .A3(new_n814), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n839), .A2(KEYINPUT53), .A3(new_n845), .A4(new_n821), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n831), .A2(KEYINPUT109), .A3(new_n832), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n835), .A2(new_n836), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(new_n805), .A3(new_n821), .A4(new_n830), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(new_n832), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n831), .A2(new_n832), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT54), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n706), .A2(new_n733), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n245), .A3(new_n400), .ZN(new_n855));
  INV_X1    g669(.A(new_n687), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n637), .A2(new_n638), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n752), .A2(new_n400), .A3(new_n854), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n729), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n679), .A2(new_n546), .A3(new_n705), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n752), .A2(new_n400), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n864), .A3(new_n724), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT50), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n704), .A2(new_n532), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT101), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n544), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n776), .A2(new_n777), .A3(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n724), .A3(new_n733), .A4(new_n864), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n869), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n871), .A2(new_n877), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n737), .A2(new_n244), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT48), .B1(new_n860), .B2(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n881), .A2(KEYINPUT113), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(KEYINPUT113), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT48), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n859), .A2(new_n884), .A3(new_n360), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT112), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n885), .A2(KEYINPUT112), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n882), .A2(new_n883), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n864), .A2(new_n716), .A3(new_n724), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n637), .A2(new_n638), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n855), .A2(new_n891), .A3(new_n856), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n399), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT111), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n888), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n889), .B1(new_n888), .B2(new_n894), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n878), .B(new_n879), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n853), .A2(new_n897), .B1(G952), .B2(G953), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n873), .B(KEYINPUT49), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n749), .A2(new_n245), .A3(new_n544), .A4(new_n547), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n679), .B1(KEYINPUT100), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n900), .A2(KEYINPUT100), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n899), .A2(new_n856), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT115), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT115), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n898), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(G75));
  NAND3_X1  g722(.A1(new_n835), .A2(new_n846), .A3(new_n847), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(G902), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G210), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n565), .A2(new_n581), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n602), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n365), .A2(G952), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G51));
  NAND2_X1  g733(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(new_n921), .A3(new_n848), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n909), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n540), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n530), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n765), .B(KEYINPUT118), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n910), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n918), .B1(new_n927), .B2(new_n929), .ZN(G54));
  NAND3_X1  g744(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n386), .A3(new_n390), .ZN(new_n932));
  INV_X1    g746(.A(new_n918), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .A4(new_n391), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G60));
  XOR2_X1   g749(.A(new_n635), .B(KEYINPUT59), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n631), .A2(new_n633), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT119), .Z(new_n938));
  AND4_X1   g752(.A1(new_n923), .A2(new_n922), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n853), .B2(new_n936), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n918), .ZN(G63));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n243), .B1(new_n909), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n942), .B1(new_n946), .B2(new_n918), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n846), .A2(new_n847), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT109), .B1(new_n831), .B2(new_n832), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n243), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(KEYINPUT121), .A3(new_n933), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n909), .A2(new_n657), .A3(new_n658), .A4(new_n945), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n947), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XOR2_X1   g769(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT61), .A4(new_n933), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(G66));
  INV_X1    g773(.A(G224), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n403), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n805), .B2(G953), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n561), .B(new_n564), .C1(G898), .C2(new_n365), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  NAND2_X1  g778(.A1(new_n668), .A2(G953), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT123), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n772), .A2(new_n360), .A3(new_n726), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n968), .A2(new_n744), .A3(new_n747), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n840), .A2(new_n698), .A3(new_n843), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n783), .A2(new_n969), .A3(new_n773), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n967), .B1(new_n971), .B2(new_n365), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n361), .A2(new_n362), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n346), .B(new_n973), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n972), .A2(KEYINPUT124), .A3(new_n974), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n891), .A2(new_n788), .A3(new_n790), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n976), .A2(new_n360), .A3(new_n690), .A4(new_n733), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n783), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n970), .A2(new_n694), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n978), .A2(new_n980), .A3(new_n773), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n365), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n974), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT124), .B1(new_n972), .B2(new_n974), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n975), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n365), .B1(G227), .B2(G900), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT125), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT122), .B1(new_n983), .B2(new_n974), .ZN(new_n992));
  INV_X1    g806(.A(new_n987), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n972), .B2(new_n974), .ZN(new_n994));
  OR3_X1    g808(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n986), .A2(new_n996), .A3(new_n987), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n989), .A2(new_n995), .A3(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  INV_X1    g814(.A(new_n805), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n971), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n347), .B(KEYINPUT127), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1003), .A2(new_n251), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n918), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n347), .A2(new_n251), .ZN(new_n1006));
  OAI221_X1 g820(.A(new_n1000), .B1(new_n1006), .B2(new_n333), .C1(new_n850), .C2(new_n851), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1000), .B1(new_n982), .B2(new_n1001), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT126), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1003), .A2(new_n251), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(G57));
endmodule


