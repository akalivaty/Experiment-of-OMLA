//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n462), .B1(new_n467), .B2(G2105), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n460), .C1(new_n463), .C2(new_n464), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G137), .A4(new_n460), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n468), .A2(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n460), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n478), .B(new_n483), .C1(G124), .C2(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(G126), .A2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n479), .B2(new_n480), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n460), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT69), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n460), .C1(new_n463), .C2(new_n464), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n471), .A2(new_n501), .A3(G138), .A4(new_n460), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n491), .A2(new_n498), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT5), .B(G543), .Z(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n510), .A2(KEYINPUT70), .A3(G63), .A4(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(new_n522), .B1(G51), .B2(new_n507), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n509), .A2(new_n510), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n525), .A2(G89), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n507), .A2(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n511), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n515), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n525), .A2(G81), .B1(G43), .B2(new_n507), .ZN(new_n539));
  XOR2_X1   g114(.A(new_n539), .B(KEYINPUT72), .Z(new_n540));
  AOI22_X1  g115(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n515), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  NAND2_X1  g123(.A1(new_n507), .A2(G53), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(KEYINPUT9), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(KEYINPUT9), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n550), .A2(new_n551), .B1(G91), .B2(new_n525), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n519), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND2_X1  g137(.A1(new_n525), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n507), .A2(G49), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  NAND2_X1  g141(.A1(G73), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G61), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n519), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(G48), .B2(new_n507), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n511), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n511), .A2(new_n572), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n573), .A3(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(new_n507), .A2(G47), .ZN(new_n577));
  XOR2_X1   g152(.A(KEYINPUT75), .B(G85), .Z(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n511), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n515), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G290));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NOR2_X1   g159(.A1(G301), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n525), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  NAND2_X1  g162(.A1(new_n510), .A2(G66), .ZN(new_n588));
  INV_X1    g163(.A(G79), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT76), .B1(new_n589), .B2(new_n504), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n589), .A2(new_n504), .A3(KEYINPUT76), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n507), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT77), .Z(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n585), .B1(new_n596), .B2(new_n584), .ZN(G284));
  AOI21_X1  g172(.A(new_n585), .B1(new_n596), .B2(new_n584), .ZN(G321));
  NOR2_X1   g173(.A1(G168), .A2(new_n584), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n584), .B2(G299), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT78), .ZN(G297));
  XNOR2_X1  g176(.A(new_n600), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n540), .A2(new_n542), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n584), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n595), .A2(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n584), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n471), .A2(new_n461), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(G2100), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT80), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n481), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n484), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n460), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2096), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n613), .B2(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n629), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT17), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT81), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n641), .ZN(new_n646));
  INV_X1    g221(.A(new_n639), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n646), .B(new_n643), .C1(new_n647), .C2(new_n641), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n641), .A3(new_n642), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2096), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n655), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G229));
  XNOR2_X1  g246(.A(KEYINPUT30), .B(G28), .ZN(new_n672));
  INV_X1    g247(.A(G29), .ZN(new_n673));
  OR2_X1    g248(.A1(KEYINPUT31), .A2(G11), .ZN(new_n674));
  NAND2_X1  g249(.A1(KEYINPUT31), .A2(G11), .ZN(new_n675));
  AOI22_X1  g250(.A1(new_n672), .A2(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n620), .B2(new_n673), .ZN(new_n677));
  NOR2_X1   g252(.A1(G162), .A2(new_n673), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n673), .B2(G35), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT29), .B(G2090), .Z(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NOR2_X1   g257(.A1(G171), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G5), .B2(new_n682), .ZN(new_n684));
  INV_X1    g259(.A(G1961), .ZN(new_n685));
  OAI221_X1 g260(.A(new_n681), .B1(new_n679), .B2(new_n680), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(G164), .A2(new_n673), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G27), .B2(new_n673), .ZN(new_n688));
  INV_X1    g263(.A(G2078), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(G160), .A2(G29), .ZN(new_n692));
  INV_X1    g267(.A(G34), .ZN(new_n693));
  AOI21_X1  g268(.A(G29), .B1(new_n693), .B2(KEYINPUT24), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(KEYINPUT24), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G2084), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n690), .A2(new_n691), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT25), .ZN(new_n700));
  NAND2_X1  g275(.A1(G103), .A2(G2104), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(G2105), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n481), .A2(G139), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n460), .B2(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G33), .B(new_n706), .S(G29), .Z(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G2072), .Z(new_n708));
  INV_X1    g283(.A(new_n684), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(G1961), .B2(new_n709), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n686), .A2(new_n699), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n673), .A2(G32), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT26), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n461), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n714), .B(new_n716), .C1(G129), .C2(new_n484), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n712), .B1(new_n717), .B2(new_n673), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT93), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT27), .B(G1996), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G168), .A2(new_n682), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n682), .B2(G21), .ZN(new_n723));
  INV_X1    g298(.A(G1966), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n696), .A2(new_n697), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT92), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n711), .A2(new_n721), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n723), .A2(new_n724), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT94), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n682), .A2(G20), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT95), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT23), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G299), .B2(G16), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT96), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1956), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n682), .A2(G4), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n596), .B2(new_n682), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT86), .B(G1348), .Z(new_n740));
  XOR2_X1   g315(.A(new_n739), .B(new_n740), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n682), .A2(G19), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT87), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n543), .B2(new_n682), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT89), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT88), .B(G1341), .Z(new_n746));
  XOR2_X1   g321(.A(new_n745), .B(new_n746), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n673), .A2(G26), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT28), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n484), .A2(G128), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT90), .Z(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(G116), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G2105), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G140), .B2(new_n481), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n749), .B1(new_n756), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n741), .A2(new_n747), .A3(new_n759), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n728), .B(new_n737), .C1(new_n760), .C2(KEYINPUT91), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n682), .A2(G23), .ZN(new_n762));
  INV_X1    g337(.A(G288), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n682), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT33), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1976), .ZN(new_n766));
  MUX2_X1   g341(.A(G6), .B(G305), .S(G16), .Z(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT32), .B(G1981), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G22), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G166), .B2(G16), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT84), .B(G1971), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n766), .A2(new_n769), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT34), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(KEYINPUT34), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n481), .A2(G131), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n484), .A2(G119), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n460), .A2(G107), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G25), .B(new_n782), .S(G29), .Z(new_n783));
  XOR2_X1   g358(.A(KEYINPUT35), .B(G1991), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G16), .A2(G24), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n582), .B(KEYINPUT82), .Z(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT83), .B(G1986), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n776), .A2(new_n777), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(KEYINPUT85), .A2(KEYINPUT36), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n791), .B(new_n792), .Z(new_n793));
  OR2_X1    g368(.A1(new_n760), .A2(KEYINPUT91), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n761), .A2(new_n793), .A3(new_n794), .ZN(G150));
  INV_X1    g370(.A(G150), .ZN(G311));
  AOI22_X1  g371(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(new_n515), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n525), .A2(G93), .B1(G55), .B2(new_n507), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G860), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT37), .Z(new_n803));
  OAI21_X1  g378(.A(new_n801), .B1(new_n543), .B2(KEYINPUT97), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n540), .A2(KEYINPUT97), .A3(new_n542), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n596), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT98), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G860), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n803), .B1(new_n814), .B2(new_n816), .ZN(G145));
  XNOR2_X1  g392(.A(new_n756), .B(new_n706), .ZN(new_n818));
  AOI22_X1  g393(.A1(G130), .A2(new_n484), .B1(new_n481), .B2(G142), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n820), .A2(new_n460), .A3(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n460), .B2(G118), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n819), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n818), .B(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n782), .B(KEYINPUT100), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n611), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n487), .A2(new_n490), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n501), .B1(new_n481), .B2(G138), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n828), .B(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT101), .B1(new_n833), .B2(new_n717), .ZN(new_n834));
  XOR2_X1   g409(.A(G162), .B(new_n620), .Z(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(G160), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n837), .C1(new_n717), .C2(new_n833), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n492), .A2(new_n497), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n500), .B2(new_n502), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n828), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n828), .A2(new_n840), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n717), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n833), .A2(new_n717), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n836), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n838), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g425(.A(new_n808), .B(new_n607), .Z(new_n851));
  XOR2_X1   g426(.A(new_n594), .B(G299), .Z(new_n852));
  INV_X1    g427(.A(KEYINPUT41), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(KEYINPUT102), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n853), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(KEYINPUT102), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n851), .A2(new_n852), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n861));
  XOR2_X1   g436(.A(G288), .B(KEYINPUT104), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G305), .ZN(new_n863));
  XOR2_X1   g438(.A(G166), .B(new_n582), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(KEYINPUT42), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n865), .B(KEYINPUT105), .Z(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n868), .B2(KEYINPUT42), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n860), .A2(new_n861), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n860), .B2(new_n861), .ZN(new_n871));
  OAI21_X1  g446(.A(G868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n801), .A2(new_n584), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(G295));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n873), .ZN(G331));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n876));
  XNOR2_X1  g451(.A(G168), .B(G301), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n808), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n806), .A2(new_n807), .A3(new_n877), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n852), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n855), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n884), .B2(new_n867), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI211_X1 g461(.A(KEYINPUT106), .B(new_n881), .C1(new_n882), .C2(new_n856), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n881), .A2(KEYINPUT106), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n867), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n868), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n867), .A3(new_n888), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n848), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n876), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n848), .A3(new_n894), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n897), .A2(KEYINPUT43), .B1(new_n898), .B2(new_n885), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n896), .B1(new_n876), .B2(new_n899), .ZN(G397));
  NOR2_X1   g475(.A1(new_n840), .A2(G1384), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(KEYINPUT45), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n717), .B(G1996), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n756), .B(new_n758), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n782), .B(new_n784), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n582), .B(G1986), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n500), .A2(new_n502), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n487), .A2(new_n490), .A3(KEYINPUT69), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n493), .B1(new_n492), .B2(new_n497), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT50), .ZN(new_n916));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n918), .B(new_n903), .C1(new_n916), .C2(new_n901), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(G2090), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(G1384), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n832), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(G164), .B2(G1384), .ZN(new_n925));
  AOI21_X1  g500(.A(G1971), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(G8), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G303), .A2(G8), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n832), .A2(new_n916), .A3(new_n917), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n903), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT107), .B1(new_n933), .B2(G2090), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n924), .A2(new_n925), .ZN(new_n935));
  INV_X1    g510(.A(G1971), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n921), .B1(new_n901), .B2(new_n916), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n939));
  INV_X1    g514(.A(G2090), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n931), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n934), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n928), .B(KEYINPUT55), .Z(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(G8), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n903), .A2(new_n901), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n945), .A2(G8), .ZN(new_n946));
  INV_X1    g521(.A(G1981), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n570), .A2(new_n575), .A3(new_n947), .A4(new_n573), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n507), .A2(G48), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n950), .B2(new_n515), .ZN(new_n951));
  OAI21_X1  g526(.A(G1981), .B1(new_n951), .B2(new_n574), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(KEYINPUT108), .A2(KEYINPUT49), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n948), .B(new_n952), .C1(KEYINPUT108), .C2(KEYINPUT49), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n946), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n763), .A2(G1976), .ZN(new_n958));
  INV_X1    g533(.A(G1976), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT52), .B1(G288), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n946), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n945), .A2(new_n958), .A3(G8), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT52), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n957), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n930), .A2(new_n944), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n932), .A2(new_n903), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n931), .A2(KEYINPUT115), .A3(new_n903), .A4(new_n932), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n685), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n832), .A2(new_n923), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n925), .A2(new_n689), .A3(new_n903), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n903), .B1(new_n901), .B2(KEYINPUT45), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  INV_X1    g553(.A(new_n923), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n978), .B1(G164), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n915), .A2(KEYINPUT109), .A3(new_n923), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n974), .A2(G2078), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n977), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n971), .A2(new_n975), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT119), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(G171), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(G171), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT119), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n965), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n938), .A2(new_n697), .A3(new_n931), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n980), .A2(new_n981), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n976), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n990), .B1(new_n992), .B2(G1966), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(G8), .A3(G286), .ZN(new_n994));
  OAI211_X1 g569(.A(G168), .B(new_n990), .C1(new_n992), .C2(G1966), .ZN(new_n995));
  AND2_X1   g570(.A1(KEYINPUT118), .A2(G8), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n995), .A2(KEYINPUT51), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT51), .B1(new_n995), .B2(new_n996), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n989), .B(KEYINPUT123), .C1(KEYINPUT62), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT123), .B1(new_n1003), .B2(new_n989), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n992), .A2(new_n982), .B1(new_n974), .B2(new_n973), .ZN(new_n1006));
  AOI211_X1 g581(.A(KEYINPUT119), .B(G301), .C1(new_n1006), .C2(new_n971), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n985), .B1(new_n984), .B2(G171), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n689), .A2(KEYINPUT120), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n974), .B1(KEYINPUT120), .B2(new_n689), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n977), .A2(new_n972), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n971), .A2(new_n975), .A3(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(G171), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT54), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n930), .A2(new_n944), .A3(new_n964), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(G171), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(KEYINPUT54), .C1(G171), .C2(new_n984), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n999), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT121), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n988), .A2(new_n986), .A3(new_n1014), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n995), .A2(new_n996), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n995), .A2(KEYINPUT51), .A3(new_n996), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n965), .B1(new_n1029), .B2(new_n994), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1023), .A2(new_n1024), .A3(new_n1030), .A4(new_n1018), .ZN(new_n1031));
  XNOR2_X1  g606(.A(G299), .B(KEYINPUT57), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT56), .B(G2072), .Z(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT113), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n925), .A2(new_n903), .A3(new_n972), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n924), .A2(KEYINPUT114), .A3(new_n925), .A4(new_n1034), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT112), .B(G1956), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1037), .A2(new_n1038), .B1(new_n919), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1032), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n919), .A2(new_n1039), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1043), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(G299), .B(KEYINPUT57), .Z(new_n1047));
  AND2_X1   g622(.A1(new_n1047), .A2(new_n1040), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n594), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n969), .A2(new_n740), .A3(new_n970), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n903), .A2(new_n901), .A3(new_n758), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1046), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1047), .A2(new_n1040), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT61), .B(new_n1054), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1047), .A2(new_n1040), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(new_n1048), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1996), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n924), .A2(new_n1059), .A3(new_n925), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  NAND2_X1  g636(.A1(new_n945), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n605), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1055), .A2(new_n1058), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT60), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n587), .B(new_n593), .C1(new_n1052), .C2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1050), .A2(KEYINPUT60), .A3(new_n594), .A4(new_n1051), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1068), .A2(new_n1069), .B1(new_n1067), .B2(new_n1052), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1053), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1020), .A2(new_n1031), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n957), .A2(new_n959), .A3(new_n763), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n948), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n946), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n961), .A2(new_n957), .A3(new_n963), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n944), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n993), .A2(G8), .A3(G168), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT63), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n942), .A2(G8), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1076), .B1(new_n1081), .B2(new_n929), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n944), .B(new_n1080), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT110), .B(KEYINPUT63), .Z(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n965), .B2(new_n1078), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1077), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1072), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1005), .B1(new_n1090), .B2(KEYINPUT122), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1072), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n911), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n784), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n782), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n907), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(G2067), .B2(new_n756), .ZN(new_n1098));
  INV_X1    g673(.A(new_n904), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT124), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1059), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT46), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n906), .A2(new_n717), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1103), .B1(new_n904), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1106));
  XNOR2_X1  g681(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  OR3_X1    g682(.A1(new_n904), .A2(G1986), .A3(G290), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT48), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1110), .B(new_n1111), .C1(new_n909), .C2(new_n904), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1101), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT126), .B1(new_n1094), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1113), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1072), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1092), .B1(new_n1072), .B2(new_n1089), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n1005), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1115), .B(new_n1116), .C1(new_n1119), .C2(new_n911), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(new_n1120), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g696(.A(G319), .ZN(new_n1123));
  NOR3_X1   g697(.A1(G227), .A2(new_n1123), .A3(G401), .ZN(new_n1124));
  NAND2_X1  g698(.A1(new_n670), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g699(.A(new_n1125), .B(KEYINPUT127), .ZN(new_n1126));
  NAND2_X1  g700(.A1(new_n849), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g701(.A1(new_n1127), .A2(new_n899), .ZN(G308));
  OR2_X1    g702(.A1(new_n1127), .A2(new_n899), .ZN(G225));
endmodule


