//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n589, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n451), .B(new_n452), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT70), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(new_n461), .B(G125), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n461), .B1(new_n466), .B2(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n469), .C1(new_n462), .C2(new_n463), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n466), .A2(KEYINPUT71), .A3(G137), .A4(new_n469), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n469), .A2(G2104), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n472), .A2(new_n473), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n462), .A2(new_n463), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n469), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND3_X1  g061(.A1(new_n466), .A2(G126), .A3(G2105), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n491), .B(new_n492), .C1(new_n463), .C2(new_n462), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n466), .B2(new_n491), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n487), .B(new_n489), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(G543), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n506), .A2(new_n512), .ZN(G166));
  AOI22_X1  g088(.A1(new_n507), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(new_n503), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n511), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(G51), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT73), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n505), .ZN(new_n528));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n508), .A2(new_n529), .B1(new_n530), .B2(new_n511), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G171));
  INV_X1    g107(.A(new_n508), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n533), .A2(G81), .B1(new_n517), .B2(G43), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n505), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND4_X1  g116(.A1(G319), .A2(G483), .A3(G661), .A4(new_n541), .ZN(G188));
  NAND2_X1  g117(.A1(G78), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G65), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n515), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(new_n533), .B2(G91), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT9), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(G299));
  INV_X1    g124(.A(G171), .ZN(G301));
  INV_X1    g125(.A(G168), .ZN(G286));
  INV_X1    g126(.A(G166), .ZN(G303));
  OAI21_X1  g127(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n553));
  INV_X1    g128(.A(G49), .ZN(new_n554));
  INV_X1    g129(.A(G87), .ZN(new_n555));
  OAI221_X1 g130(.A(new_n553), .B1(new_n554), .B2(new_n511), .C1(new_n555), .C2(new_n508), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(G288));
  NAND3_X1  g133(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n507), .A2(new_n561), .A3(G48), .A4(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G61), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n501), .B2(new_n502), .ZN(new_n565));
  AND2_X1   g140(.A1(G73), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n503), .A2(G86), .A3(new_n507), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(G305));
  AOI22_X1  g144(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n505), .ZN(new_n571));
  XNOR2_X1  g146(.A(KEYINPUT77), .B(G85), .ZN(new_n572));
  INV_X1    g147(.A(G47), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n508), .A2(new_n572), .B1(new_n573), .B2(new_n511), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n503), .A2(G92), .A3(new_n507), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G66), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n515), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G284));
  OAI21_X1  g161(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G321));
  XOR2_X1   g162(.A(G299), .B(KEYINPUT78), .Z(new_n588));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  MUX2_X1   g164(.A(G286), .B(new_n588), .S(new_n589), .Z(G297));
  MUX2_X1   g165(.A(G286), .B(new_n588), .S(new_n589), .Z(G280));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n585), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G868), .B2(new_n537), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g172(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n598));
  INV_X1    g173(.A(G111), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G2105), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n481), .A2(G123), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AOI211_X1 g178(.A(new_n600), .B(new_n603), .C1(G135), .C2(new_n479), .ZN(new_n604));
  INV_X1    g179(.A(G2096), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n466), .A2(new_n474), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n606), .A2(new_n607), .A3(new_n613), .A4(new_n614), .ZN(G156));
  INV_X1    g190(.A(G14), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT14), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2427), .B(G2430), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT82), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n619), .B2(new_n620), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n623), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n627), .B(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n616), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n632), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n635), .A2(KEYINPUT83), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n630), .B2(new_n632), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n634), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(G401));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(new_n612), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n644), .B2(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(new_n605), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT85), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n656), .A2(new_n657), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(new_n658), .ZN(new_n665));
  MUX2_X1   g240(.A(new_n665), .B(new_n664), .S(new_n655), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n673), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n673), .B2(new_n674), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(G229));
  XNOR2_X1  g256(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G34), .ZN(new_n683));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(new_n476), .B2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(G2084), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n585), .A2(G16), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G4), .B2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G1348), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n688), .B(new_n693), .C1(new_n692), .C2(new_n691), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G19), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n537), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1341), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT31), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(G11), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(G11), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n701), .A2(G28), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n684), .B1(new_n701), .B2(G28), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n699), .B(new_n700), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n604), .B2(G29), .ZN(new_n705));
  INV_X1    g280(.A(G2072), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n684), .A2(G33), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n708));
  NAND2_X1  g283(.A1(G103), .A2(G2104), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G2105), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n469), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n479), .A2(G139), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n469), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n707), .B1(new_n714), .B2(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n705), .B1(new_n706), .B2(new_n715), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n697), .B(new_n716), .C1(new_n706), .C2(new_n715), .ZN(new_n717));
  NOR2_X1   g292(.A1(G5), .A2(G16), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT96), .Z(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(G301), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT97), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n684), .A2(G32), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n479), .A2(G141), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n481), .A2(G129), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n729), .B(new_n730), .Z(new_n731));
  AOI211_X1 g306(.A(new_n728), .B(new_n731), .C1(G105), .C2(new_n474), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n684), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT95), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n684), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n684), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G2090), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n684), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n684), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2078), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n736), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n694), .A2(new_n717), .A3(new_n724), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n720), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n720), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G1966), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n720), .A2(G20), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT23), .Z(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G299), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1956), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n748), .A2(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n684), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT92), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n479), .A2(G140), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT90), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n481), .A2(G128), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT91), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n469), .A2(G116), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n760), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n758), .B1(new_n765), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n746), .A2(new_n754), .A3(new_n755), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n684), .A2(G25), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n479), .A2(G131), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(G107), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G2105), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n481), .B2(G119), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n770), .B1(new_n779), .B2(new_n684), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT89), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT35), .B(G1991), .Z(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n720), .A2(G24), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n575), .B2(new_n720), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1986), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n720), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(new_n556), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n720), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT33), .B(G1976), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n720), .A2(G22), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G166), .B2(new_n720), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G6), .B(G305), .S(G16), .Z(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT32), .B(G1981), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT34), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n798), .A2(KEYINPUT34), .A3(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n781), .A2(new_n783), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n788), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT36), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n769), .A2(new_n806), .ZN(G150));
  XOR2_X1   g382(.A(G150), .B(KEYINPUT99), .Z(G311));
  NAND2_X1  g383(.A1(new_n585), .A2(G559), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n505), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  INV_X1    g388(.A(G55), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n508), .A2(new_n813), .B1(new_n814), .B2(new_n511), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n537), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n810), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT101), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT100), .B(G860), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n818), .B2(new_n819), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n816), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n822), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(G145));
  INV_X1    g403(.A(G37), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n778), .B(new_n609), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  INV_X1    g406(.A(G118), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(G2105), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n481), .A2(G130), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT104), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n833), .B(new_n835), .C1(G142), .C2(new_n479), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n830), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n487), .A2(new_n489), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n491), .B1(new_n462), .B2(new_n463), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT4), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n841), .A2(KEYINPUT103), .A3(new_n493), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT103), .B1(new_n841), .B2(new_n493), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n765), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n714), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(new_n732), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n732), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n837), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n837), .ZN(new_n850));
  XNOR2_X1  g425(.A(G162), .B(new_n476), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT102), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n604), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n847), .A2(new_n848), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n837), .A2(KEYINPUT105), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n847), .B(new_n848), .C1(KEYINPUT105), .C2(new_n837), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI221_X1 g434(.A(new_n829), .B1(new_n849), .B2(new_n854), .C1(new_n859), .C2(new_n853), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g436(.A1(new_n825), .A2(new_n589), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n575), .B(G305), .ZN(new_n863));
  XNOR2_X1  g438(.A(G166), .B(new_n556), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n863), .B(new_n864), .Z(new_n865));
  XOR2_X1   g440(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n817), .B(new_n594), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n584), .B(G299), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n869), .A2(KEYINPUT41), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(KEYINPUT41), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT107), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n870), .B1(new_n876), .B2(new_n868), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n867), .B1(new_n877), .B2(KEYINPUT109), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(KEYINPUT109), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n867), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n862), .B1(new_n880), .B2(new_n589), .ZN(G295));
  OAI21_X1  g456(.A(new_n862), .B1(new_n880), .B2(new_n589), .ZN(G331));
  XNOR2_X1  g457(.A(G168), .B(G171), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n817), .ZN(new_n884));
  XNOR2_X1  g459(.A(G168), .B(G301), .ZN(new_n885));
  INV_X1    g460(.A(new_n817), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n888), .A2(new_n869), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n876), .B2(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(new_n865), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n888), .A2(KEYINPUT110), .A3(new_n869), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n884), .A2(new_n887), .B1(new_n871), .B2(new_n874), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT110), .B1(new_n888), .B2(new_n869), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n893), .B(new_n865), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n892), .A2(KEYINPUT43), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n890), .A2(new_n891), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT43), .B1(new_n898), .B2(new_n892), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT44), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n901), .A3(new_n896), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n898), .B2(new_n892), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n905), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g481(.A(G1384), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT45), .B1(new_n844), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n468), .A2(new_n475), .A3(G40), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n910), .B(KEYINPUT111), .Z(new_n911));
  INV_X1    g486(.A(G1996), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT46), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n765), .B(new_n767), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n732), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(KEYINPUT47), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n732), .B(G1996), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n779), .A2(new_n782), .ZN(new_n922));
  OAI22_X1  g497(.A1(new_n921), .A2(new_n922), .B1(G2067), .B2(new_n765), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n911), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n778), .A2(new_n783), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n920), .A2(new_n915), .A3(new_n922), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n911), .ZN(new_n927));
  NOR2_X1   g502(.A1(G290), .A2(G1986), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n911), .A2(KEYINPUT48), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT48), .B1(new_n911), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n924), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT125), .ZN(new_n934));
  INV_X1    g509(.A(G1976), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT52), .B1(G288), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n790), .A2(G1976), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n938));
  INV_X1    g513(.A(G8), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n494), .B2(new_n495), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n841), .A2(KEYINPUT103), .A3(new_n493), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G1384), .B1(new_n943), .B2(new_n839), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n938), .B(new_n939), .C1(new_n944), .C2(new_n909), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n909), .A2(new_n907), .A3(new_n844), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT113), .B1(new_n946), .B2(G8), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n936), .B(new_n937), .C1(new_n945), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(G305), .A2(G1981), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n563), .A2(new_n668), .A3(new_n567), .A4(new_n568), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT49), .B1(new_n951), .B2(KEYINPUT114), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT49), .ZN(new_n954));
  AOI211_X1 g529(.A(new_n953), .B(new_n954), .C1(new_n949), .C2(new_n950), .ZN(new_n955));
  OAI22_X1  g530(.A1(new_n945), .A2(new_n947), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n946), .A2(G8), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n938), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n946), .A2(KEYINPUT113), .A3(G8), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n958), .B1(new_n962), .B2(new_n937), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(G166), .A2(new_n939), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT55), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n496), .B2(new_n907), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n468), .A2(new_n475), .A3(G40), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n844), .A2(new_n967), .A3(new_n907), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(G2090), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT45), .B1(new_n496), .B2(new_n907), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(new_n969), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n844), .A2(KEYINPUT45), .A3(new_n907), .ZN(new_n976));
  AOI21_X1  g551(.A(G1971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n966), .B(G8), .C1(new_n973), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n975), .A2(new_n976), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n981), .A2(G1971), .B1(G2090), .B2(new_n972), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(KEYINPUT112), .A3(G8), .A4(new_n966), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n967), .B1(new_n844), .B2(new_n907), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n496), .A2(new_n967), .A3(new_n907), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n909), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n985), .A2(new_n987), .A3(G2090), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n988), .B2(new_n977), .ZN(new_n989));
  INV_X1    g564(.A(new_n966), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n964), .A2(new_n984), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n908), .B2(new_n969), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NOR3_X1   g570(.A1(G164), .A2(new_n995), .A3(G1384), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT116), .B(new_n909), .C1(new_n944), .C2(KEYINPUT45), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2078), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n994), .A2(new_n997), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G2078), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n975), .A2(new_n976), .A3(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1003), .A2(new_n999), .B1(new_n972), .B2(new_n723), .ZN(new_n1004));
  AOI21_X1  g579(.A(G301), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n992), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G286), .A2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(new_n1011));
  INV_X1    g586(.A(G1966), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT117), .B(G2084), .Z(new_n1014));
  AND3_X1   g589(.A1(new_n970), .A2(new_n971), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1010), .B1(new_n1017), .B2(G8), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT122), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1021), .B(new_n1015), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1020), .A2(new_n1022), .A3(G286), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1009), .A2(new_n939), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1019), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n844), .A2(new_n907), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n969), .B1(new_n1027), .B2(new_n995), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n996), .B1(new_n1028), .B2(KEYINPUT116), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1966), .B1(new_n1029), .B2(new_n994), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1021), .B1(new_n1030), .B2(new_n1015), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1015), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT122), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1008), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT62), .B1(new_n1026), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1031), .A2(G168), .A3(new_n1033), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1018), .B1(new_n1037), .B2(new_n1024), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT62), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1034), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1007), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1042));
  AOI22_X1  g617(.A1(new_n944), .A2(KEYINPUT45), .B1(KEYINPUT124), .B2(new_n969), .ZN(new_n1043));
  INV_X1    g618(.A(new_n908), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n969), .A2(KEYINPUT124), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1000), .A4(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1004), .A2(G301), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1042), .B1(new_n1047), .B2(new_n1005), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1001), .A2(new_n1004), .A3(G301), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1004), .A2(new_n1046), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT54), .B(new_n1049), .C1(new_n1050), .C2(G301), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n992), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n975), .A2(new_n976), .A3(new_n912), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT58), .B(G1341), .Z(new_n1055));
  NAND2_X1  g630(.A1(new_n946), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n537), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1057), .B(new_n537), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1348), .B1(new_n970), .B2(new_n971), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n946), .A2(G2067), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT60), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1070), .A3(new_n585), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  INV_X1    g647(.A(G1956), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n985), .B2(new_n987), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n975), .A2(new_n976), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n548), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G299), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n546), .B(new_n548), .C1(new_n1077), .C2(KEYINPUT57), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1074), .A2(new_n1076), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1072), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1067), .A2(KEYINPUT60), .A3(new_n584), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1064), .A2(new_n1071), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1074), .A2(new_n1076), .A3(new_n1081), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1083), .B2(KEYINPUT120), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1074), .A2(new_n1076), .A3(new_n1089), .A4(new_n1081), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(KEYINPUT61), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT121), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1088), .A2(new_n1093), .A3(KEYINPUT61), .A4(new_n1090), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1086), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1083), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n585), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1082), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g673(.A(new_n1053), .B1(new_n1038), .B2(new_n1034), .C1(new_n1095), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n964), .ZN(new_n1100));
  INV_X1    g675(.A(new_n950), .ZN(new_n1101));
  NOR2_X1   g676(.A1(G288), .A2(G1976), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT115), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n952), .A2(new_n955), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n962), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1100), .A2(new_n984), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1032), .A2(new_n939), .A3(G286), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n964), .A2(new_n1108), .A3(new_n984), .A4(new_n991), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n982), .A2(G8), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1112), .B2(new_n990), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n964), .A2(new_n1108), .A3(new_n984), .A4(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1107), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1041), .A2(new_n1099), .A3(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n575), .B(new_n670), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n911), .B1(new_n926), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n934), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1053), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1038), .A2(new_n1034), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1115), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1007), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1026), .A2(KEYINPUT62), .A3(new_n1035), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1039), .B1(new_n1038), .B2(new_n1034), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n934), .B(new_n1118), .C1(new_n1122), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n933), .B1(new_n1119), .B2(new_n1128), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g704(.A(G227), .ZN(new_n1131));
  NAND2_X1  g705(.A1(new_n1131), .A2(G319), .ZN(new_n1132));
  XNOR2_X1  g706(.A(new_n1132), .B(KEYINPUT126), .ZN(new_n1133));
  NAND4_X1  g707(.A1(new_n639), .A2(new_n679), .A3(new_n680), .A4(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g708(.A(new_n1134), .B(KEYINPUT127), .ZN(new_n1135));
  OAI21_X1  g709(.A(new_n860), .B1(new_n903), .B2(new_n904), .ZN(new_n1136));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n1136), .ZN(G308));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n1138));
  XNOR2_X1  g712(.A(new_n1134), .B(new_n1138), .ZN(new_n1139));
  OR2_X1    g713(.A1(new_n903), .A2(new_n904), .ZN(new_n1140));
  NAND3_X1  g714(.A1(new_n1139), .A2(new_n1140), .A3(new_n860), .ZN(G225));
endmodule


