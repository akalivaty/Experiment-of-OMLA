

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  NOR2_X2 U322 ( .A1(n553), .A2(n494), .ZN(n495) );
  XNOR2_X2 U323 ( .A(n296), .B(n295), .ZN(n434) );
  XNOR2_X1 U324 ( .A(n351), .B(n378), .ZN(n356) );
  XOR2_X1 U325 ( .A(n392), .B(n391), .Z(n545) );
  XOR2_X1 U326 ( .A(n344), .B(n377), .Z(n542) );
  INV_X1 U327 ( .A(n373), .ZN(n355) );
  XNOR2_X1 U328 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U329 ( .A(n361), .B(n360), .Z(n537) );
  XOR2_X1 U330 ( .A(KEYINPUT38), .B(n457), .Z(n466) );
  XNOR2_X1 U331 ( .A(G71GAT), .B(G57GAT), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n290), .B(KEYINPUT13), .ZN(n411) );
  XOR2_X1 U333 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n292) );
  NAND2_X1 U334 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U336 ( .A(n293), .B(KEYINPUT32), .Z(n298) );
  XNOR2_X1 U337 ( .A(G78GAT), .B(G204GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n294), .B(G148GAT), .ZN(n368) );
  XOR2_X1 U339 ( .A(G85GAT), .B(G92GAT), .Z(n296) );
  XNOR2_X1 U340 ( .A(G99GAT), .B(G106GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n368), .B(n434), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U343 ( .A(n299), .B(KEYINPUT33), .Z(n301) );
  XOR2_X1 U344 ( .A(G176GAT), .B(G64GAT), .Z(n359) );
  XNOR2_X1 U345 ( .A(G120GAT), .B(n359), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n411), .B(n302), .ZN(n570) );
  XOR2_X1 U348 ( .A(G113GAT), .B(G22GAT), .Z(n304) );
  XNOR2_X1 U349 ( .A(G141GAT), .B(G197GAT), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n305), .B(G50GAT), .Z(n307) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G1GAT), .ZN(n408) );
  XOR2_X1 U353 ( .A(n408), .B(G36GAT), .Z(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n313) );
  XOR2_X1 U355 ( .A(G29GAT), .B(G43GAT), .Z(n309) );
  XNOR2_X1 U356 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n435) );
  XOR2_X1 U358 ( .A(n435), .B(KEYINPUT66), .Z(n311) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U361 ( .A(n313), .B(n312), .Z(n321) );
  XOR2_X1 U362 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n315) );
  XNOR2_X1 U363 ( .A(G169GAT), .B(G8GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U365 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n317) );
  XNOR2_X1 U366 ( .A(KEYINPUT65), .B(KEYINPUT64), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(n321), .B(n320), .Z(n507) );
  INV_X1 U370 ( .A(n507), .ZN(n567) );
  NOR2_X1 U371 ( .A1(n570), .A2(n567), .ZN(n322) );
  XOR2_X1 U372 ( .A(n322), .B(KEYINPUT70), .Z(n452) );
  XOR2_X1 U373 ( .A(KEYINPUT1), .B(G57GAT), .Z(n324) );
  XNOR2_X1 U374 ( .A(G1GAT), .B(G148GAT), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U376 ( .A(KEYINPUT85), .B(KEYINPUT6), .Z(n326) );
  XNOR2_X1 U377 ( .A(KEYINPUT4), .B(KEYINPUT84), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U379 ( .A(n328), .B(n327), .Z(n339) );
  XOR2_X1 U380 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n330) );
  XNOR2_X1 U381 ( .A(KEYINPUT3), .B(KEYINPUT83), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U383 ( .A(G141GAT), .B(n331), .Z(n374) );
  XOR2_X1 U384 ( .A(G85GAT), .B(G155GAT), .Z(n333) );
  XNOR2_X1 U385 ( .A(G29GAT), .B(G162GAT), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U387 ( .A(KEYINPUT5), .B(n334), .Z(n336) );
  NAND2_X1 U388 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n374), .B(n337), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n344) );
  XOR2_X1 U392 ( .A(KEYINPUT0), .B(G120GAT), .Z(n341) );
  XNOR2_X1 U393 ( .A(G113GAT), .B(G127GAT), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n343) );
  XOR2_X1 U395 ( .A(G134GAT), .B(KEYINPUT75), .Z(n342) );
  XOR2_X1 U396 ( .A(n343), .B(n342), .Z(n377) );
  XOR2_X1 U397 ( .A(G92GAT), .B(KEYINPUT86), .Z(n346) );
  NAND2_X1 U398 ( .A1(G226GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U400 ( .A(n347), .B(G204GAT), .Z(n351) );
  XOR2_X1 U401 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n349) );
  XNOR2_X1 U402 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(n350), .ZN(n378) );
  XOR2_X1 U405 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n353) );
  XNOR2_X1 U406 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U408 ( .A(G197GAT), .B(n354), .Z(n373) );
  XOR2_X1 U409 ( .A(G8GAT), .B(G183GAT), .Z(n418) );
  XOR2_X1 U410 ( .A(n357), .B(n418), .Z(n361) );
  XNOR2_X1 U411 ( .A(G36GAT), .B(G190GAT), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n358), .B(G218GAT), .ZN(n427) );
  XNOR2_X1 U413 ( .A(n427), .B(n359), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n537), .B(KEYINPUT87), .ZN(n362) );
  XOR2_X1 U415 ( .A(KEYINPUT27), .B(n362), .Z(n401) );
  XOR2_X1 U416 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n364) );
  XNOR2_X1 U417 ( .A(KEYINPUT79), .B(KEYINPUT22), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U419 ( .A(n365), .B(G106GAT), .Z(n367) );
  XOR2_X1 U420 ( .A(G22GAT), .B(G155GAT), .Z(n419) );
  XNOR2_X1 U421 ( .A(n419), .B(G218GAT), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n372) );
  XNOR2_X1 U423 ( .A(G50GAT), .B(G162GAT), .ZN(n424) );
  XNOR2_X1 U424 ( .A(n368), .B(n424), .ZN(n370) );
  NAND2_X1 U425 ( .A1(G228GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U427 ( .A(n372), .B(n371), .Z(n376) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n543) );
  INV_X1 U430 ( .A(n377), .ZN(n392) );
  INV_X1 U431 ( .A(n378), .ZN(n386) );
  NAND2_X1 U432 ( .A1(G227GAT), .A2(G233GAT), .ZN(n384) );
  XOR2_X1 U433 ( .A(G176GAT), .B(G183GAT), .Z(n380) );
  XNOR2_X1 U434 ( .A(G43GAT), .B(G71GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U436 ( .A(G190GAT), .B(G99GAT), .Z(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U439 ( .A(n386), .B(n385), .Z(n390) );
  XOR2_X1 U440 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n388) );
  XNOR2_X1 U441 ( .A(G15GAT), .B(KEYINPUT76), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n391) );
  NOR2_X1 U444 ( .A1(n543), .A2(n545), .ZN(n394) );
  XNOR2_X1 U445 ( .A(KEYINPUT26), .B(KEYINPUT88), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n565) );
  NAND2_X1 U447 ( .A1(n401), .A2(n565), .ZN(n522) );
  XNOR2_X1 U448 ( .A(n522), .B(KEYINPUT89), .ZN(n395) );
  NOR2_X1 U449 ( .A1(n542), .A2(n395), .ZN(n400) );
  NAND2_X1 U450 ( .A1(n545), .A2(n537), .ZN(n396) );
  NAND2_X1 U451 ( .A1(n396), .A2(n543), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n397), .B(KEYINPUT90), .ZN(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT25), .B(n398), .Z(n399) );
  NAND2_X1 U454 ( .A1(n400), .A2(n399), .ZN(n406) );
  INV_X1 U455 ( .A(n545), .ZN(n403) );
  XOR2_X1 U456 ( .A(n543), .B(KEYINPUT28), .Z(n487) );
  INV_X1 U457 ( .A(n401), .ZN(n402) );
  NOR2_X1 U458 ( .A1(n487), .A2(n402), .ZN(n505) );
  NAND2_X1 U459 ( .A1(n403), .A2(n505), .ZN(n404) );
  NAND2_X1 U460 ( .A1(n404), .A2(n542), .ZN(n405) );
  NAND2_X1 U461 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U462 ( .A(KEYINPUT91), .B(n407), .ZN(n454) );
  XNOR2_X1 U463 ( .A(G211GAT), .B(G78GAT), .ZN(n410) );
  INV_X1 U464 ( .A(n408), .ZN(n409) );
  XOR2_X1 U465 ( .A(n410), .B(n409), .Z(n423) );
  XOR2_X1 U466 ( .A(n411), .B(KEYINPUT15), .Z(n413) );
  NAND2_X1 U467 ( .A1(G231GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U469 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n415) );
  XNOR2_X1 U470 ( .A(G127GAT), .B(G64GAT), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U472 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U475 ( .A(n423), .B(n422), .Z(n530) );
  INV_X1 U476 ( .A(n530), .ZN(n574) );
  XNOR2_X1 U477 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n426) );
  INV_X1 U478 ( .A(n424), .ZN(n425) );
  XOR2_X1 U479 ( .A(n426), .B(n425), .Z(n439) );
  XOR2_X1 U480 ( .A(n427), .B(KEYINPUT11), .Z(n429) );
  NAND2_X1 U481 ( .A1(G232GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U483 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n431) );
  XNOR2_X1 U484 ( .A(G134GAT), .B(KEYINPUT73), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U486 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U489 ( .A(n439), .B(n438), .ZN(n535) );
  XNOR2_X1 U490 ( .A(n535), .B(KEYINPUT74), .ZN(n558) );
  NAND2_X1 U491 ( .A1(n574), .A2(n558), .ZN(n440) );
  XOR2_X1 U492 ( .A(KEYINPUT16), .B(n440), .Z(n441) );
  NAND2_X1 U493 ( .A1(n454), .A2(n441), .ZN(n469) );
  NOR2_X1 U494 ( .A1(n452), .A2(n469), .ZN(n450) );
  NAND2_X1 U495 ( .A1(n450), .A2(n542), .ZN(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n443) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(G1324GAT) );
  NAND2_X1 U500 ( .A1(n537), .A2(n450), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n446), .B(KEYINPUT94), .ZN(n447) );
  XNOR2_X1 U502 ( .A(G8GAT), .B(n447), .ZN(G1325GAT) );
  XOR2_X1 U503 ( .A(G15GAT), .B(KEYINPUT35), .Z(n449) );
  NAND2_X1 U504 ( .A1(n450), .A2(n545), .ZN(n448) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(G1326GAT) );
  NAND2_X1 U506 ( .A1(n450), .A2(n487), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n451), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U508 ( .A(G29GAT), .B(KEYINPUT95), .Z(n459) );
  INV_X1 U509 ( .A(n452), .ZN(n456) );
  XNOR2_X1 U510 ( .A(KEYINPUT36), .B(n558), .ZN(n581) );
  NOR2_X1 U511 ( .A1(n574), .A2(n581), .ZN(n453) );
  NAND2_X1 U512 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(KEYINPUT37), .B(n455), .ZN(n482) );
  NAND2_X1 U514 ( .A1(n456), .A2(n482), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n542), .A2(n466), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n461) );
  XOR2_X1 U517 ( .A(KEYINPUT39), .B(KEYINPUT96), .Z(n460) );
  XNOR2_X1 U518 ( .A(n461), .B(n460), .ZN(G1328GAT) );
  NAND2_X1 U519 ( .A1(n466), .A2(n537), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n462), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U521 ( .A(KEYINPUT97), .B(KEYINPUT40), .Z(n464) );
  NAND2_X1 U522 ( .A1(n466), .A2(n545), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U524 ( .A(G43GAT), .B(n465), .ZN(G1330GAT) );
  NAND2_X1 U525 ( .A1(n466), .A2(n487), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT98), .ZN(n468) );
  XNOR2_X1 U527 ( .A(G50GAT), .B(n468), .ZN(G1331GAT) );
  XNOR2_X1 U528 ( .A(KEYINPUT41), .B(n570), .ZN(n527) );
  XOR2_X1 U529 ( .A(n527), .B(KEYINPUT99), .Z(n548) );
  NOR2_X1 U530 ( .A1(n548), .A2(n507), .ZN(n481) );
  INV_X1 U531 ( .A(n481), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n470), .A2(n469), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n542), .A2(n476), .ZN(n471) );
  XNOR2_X1 U534 ( .A(KEYINPUT42), .B(n471), .ZN(n472) );
  XNOR2_X1 U535 ( .A(G57GAT), .B(n472), .ZN(G1332GAT) );
  NAND2_X1 U536 ( .A1(n537), .A2(n476), .ZN(n473) );
  XNOR2_X1 U537 ( .A(n473), .B(KEYINPUT100), .ZN(n474) );
  XNOR2_X1 U538 ( .A(G64GAT), .B(n474), .ZN(G1333GAT) );
  NAND2_X1 U539 ( .A1(n545), .A2(n476), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n475), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n478) );
  NAND2_X1 U542 ( .A1(n476), .A2(n487), .ZN(n477) );
  XNOR2_X1 U543 ( .A(n478), .B(n477), .ZN(n480) );
  XOR2_X1 U544 ( .A(G78GAT), .B(KEYINPUT102), .Z(n479) );
  XNOR2_X1 U545 ( .A(n480), .B(n479), .ZN(G1335GAT) );
  AND2_X1 U546 ( .A1(n482), .A2(n481), .ZN(n488) );
  NAND2_X1 U547 ( .A1(n488), .A2(n542), .ZN(n483) );
  XNOR2_X1 U548 ( .A(n483), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U549 ( .A(G92GAT), .B(KEYINPUT103), .Z(n485) );
  NAND2_X1 U550 ( .A1(n488), .A2(n537), .ZN(n484) );
  XNOR2_X1 U551 ( .A(n485), .B(n484), .ZN(G1337GAT) );
  NAND2_X1 U552 ( .A1(n545), .A2(n488), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n486), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U554 ( .A(G106GAT), .B(KEYINPUT104), .ZN(n492) );
  XOR2_X1 U555 ( .A(KEYINPUT105), .B(KEYINPUT44), .Z(n490) );
  NAND2_X1 U556 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U557 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U558 ( .A(n492), .B(n491), .ZN(G1339GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n509) );
  XOR2_X1 U560 ( .A(KEYINPUT107), .B(KEYINPUT47), .Z(n497) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(n530), .Z(n553) );
  NOR2_X1 U562 ( .A1(n567), .A2(n527), .ZN(n493) );
  XNOR2_X1 U563 ( .A(n493), .B(KEYINPUT46), .ZN(n494) );
  NAND2_X1 U564 ( .A1(n495), .A2(n535), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n497), .B(n496), .ZN(n503) );
  NOR2_X1 U566 ( .A1(n581), .A2(n530), .ZN(n499) );
  XNOR2_X1 U567 ( .A(KEYINPUT45), .B(KEYINPUT108), .ZN(n498) );
  XNOR2_X1 U568 ( .A(n499), .B(n498), .ZN(n501) );
  NOR2_X1 U569 ( .A1(n507), .A2(n570), .ZN(n500) );
  AND2_X1 U570 ( .A1(n501), .A2(n500), .ZN(n502) );
  NOR2_X1 U571 ( .A1(n503), .A2(n502), .ZN(n504) );
  XOR2_X1 U572 ( .A(KEYINPUT48), .B(n504), .Z(n538) );
  NAND2_X1 U573 ( .A1(n538), .A2(n542), .ZN(n521) );
  NAND2_X1 U574 ( .A1(n505), .A2(n545), .ZN(n506) );
  NOR2_X1 U575 ( .A1(n521), .A2(n506), .ZN(n514) );
  NAND2_X1 U576 ( .A1(n514), .A2(n507), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U578 ( .A(G113GAT), .B(n510), .ZN(G1340GAT) );
  INV_X1 U579 ( .A(n514), .ZN(n517) );
  NOR2_X1 U580 ( .A1(n548), .A2(n517), .ZN(n512) );
  XNOR2_X1 U581 ( .A(KEYINPUT111), .B(KEYINPUT49), .ZN(n511) );
  XNOR2_X1 U582 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U583 ( .A(G120GAT), .B(n513), .Z(G1341GAT) );
  NAND2_X1 U584 ( .A1(n553), .A2(n514), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n515), .B(KEYINPUT50), .ZN(n516) );
  XNOR2_X1 U586 ( .A(G127GAT), .B(n516), .ZN(G1342GAT) );
  NOR2_X1 U587 ( .A1(n558), .A2(n517), .ZN(n519) );
  XNOR2_X1 U588 ( .A(KEYINPUT51), .B(KEYINPUT112), .ZN(n518) );
  XNOR2_X1 U589 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U590 ( .A(G134GAT), .B(n520), .ZN(G1343GAT) );
  NOR2_X1 U591 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U592 ( .A(KEYINPUT113), .B(n523), .ZN(n534) );
  NOR2_X1 U593 ( .A1(n567), .A2(n534), .ZN(n524) );
  XOR2_X1 U594 ( .A(G141GAT), .B(n524), .Z(G1344GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT52), .B(KEYINPUT114), .Z(n526) );
  XNOR2_X1 U596 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n525) );
  XNOR2_X1 U597 ( .A(n526), .B(n525), .ZN(n529) );
  NOR2_X1 U598 ( .A1(n527), .A2(n534), .ZN(n528) );
  XOR2_X1 U599 ( .A(n529), .B(n528), .Z(G1345GAT) );
  NOR2_X1 U600 ( .A1(n530), .A2(n534), .ZN(n532) );
  XNOR2_X1 U601 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U603 ( .A(G155GAT), .B(n533), .ZN(G1346GAT) );
  NOR2_X1 U604 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U605 ( .A(G162GAT), .B(n536), .Z(G1347GAT) );
  AND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n539), .B(KEYINPUT54), .ZN(n540) );
  XNOR2_X1 U608 ( .A(KEYINPUT117), .B(n540), .ZN(n541) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n564) );
  NAND2_X1 U610 ( .A1(n564), .A2(n543), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n544), .B(KEYINPUT55), .ZN(n546) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n559) );
  NOR2_X1 U613 ( .A1(n567), .A2(n559), .ZN(n547) );
  XOR2_X1 U614 ( .A(G169GAT), .B(n547), .Z(G1348GAT) );
  NOR2_X1 U615 ( .A1(n548), .A2(n559), .ZN(n550) );
  XNOR2_X1 U616 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G176GAT), .ZN(G1349GAT) );
  INV_X1 U619 ( .A(n559), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G183GAT), .B(n555), .ZN(G1350GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT119), .B(KEYINPUT58), .Z(n557) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(n561), .B(n560), .Z(G1351GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n563) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT121), .B(n566), .ZN(n575) );
  INV_X1 U633 ( .A(n575), .ZN(n580) );
  NOR2_X1 U634 ( .A1(n567), .A2(n580), .ZN(n568) );
  XOR2_X1 U635 ( .A(n569), .B(n568), .Z(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U637 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT124), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n579) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1355GAT) );
endmodule

