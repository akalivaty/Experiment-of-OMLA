

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  XOR2_X1 U325 ( .A(G85GAT), .B(KEYINPUT74), .Z(n387) );
  XNOR2_X1 U326 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U327 ( .A(n399), .B(n398), .ZN(n405) );
  XNOR2_X1 U328 ( .A(KEYINPUT123), .B(n454), .ZN(n566) );
  XNOR2_X1 U329 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U330 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(G78GAT), .B(G148GAT), .Z(n294) );
  XNOR2_X1 U332 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n294), .B(n293), .ZN(n383) );
  XOR2_X1 U334 ( .A(n383), .B(G197GAT), .Z(n296) );
  XOR2_X1 U335 ( .A(G141GAT), .B(G22GAT), .Z(n369) );
  XNOR2_X1 U336 ( .A(G50GAT), .B(n369), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n302) );
  XOR2_X1 U338 ( .A(G155GAT), .B(KEYINPUT2), .Z(n298) );
  XNOR2_X1 U339 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n322) );
  XOR2_X1 U341 ( .A(n322), .B(KEYINPUT23), .Z(n300) );
  NAND2_X1 U342 ( .A1(G228GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U344 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U345 ( .A(KEYINPUT21), .B(G218GAT), .Z(n304) );
  XNOR2_X1 U346 ( .A(G211GAT), .B(G204GAT), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U348 ( .A(KEYINPUT92), .B(n305), .Z(n432) );
  XOR2_X1 U349 ( .A(KEYINPUT22), .B(KEYINPUT94), .Z(n307) );
  XNOR2_X1 U350 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n432), .B(n308), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n466) );
  XOR2_X1 U354 ( .A(G57GAT), .B(G120GAT), .Z(n312) );
  XNOR2_X1 U355 ( .A(G113GAT), .B(G1GAT), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U357 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n314) );
  XNOR2_X1 U358 ( .A(KEYINPUT96), .B(KEYINPUT6), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U360 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U361 ( .A(KEYINPUT4), .B(KEYINPUT97), .Z(n318) );
  NAND2_X1 U362 ( .A1(G225GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U364 ( .A(KEYINPUT95), .B(n319), .ZN(n320) );
  XNOR2_X1 U365 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U366 ( .A(G85GAT), .B(G148GAT), .Z(n324) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(n322), .ZN(n323) );
  XNOR2_X1 U368 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U369 ( .A(n326), .B(n325), .Z(n332) );
  XOR2_X1 U370 ( .A(KEYINPUT86), .B(G134GAT), .Z(n328) );
  XNOR2_X1 U371 ( .A(KEYINPUT85), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U372 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U373 ( .A(KEYINPUT0), .B(n329), .ZN(n451) );
  INV_X1 U374 ( .A(n451), .ZN(n330) );
  XNOR2_X1 U375 ( .A(G141GAT), .B(n330), .ZN(n331) );
  XNOR2_X1 U376 ( .A(n332), .B(n331), .ZN(n522) );
  INV_X1 U377 ( .A(n522), .ZN(n506) );
  INV_X1 U378 ( .A(KEYINPUT47), .ZN(n409) );
  XOR2_X1 U379 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n334) );
  XNOR2_X1 U380 ( .A(KEYINPUT82), .B(KEYINPUT84), .ZN(n333) );
  XNOR2_X1 U381 ( .A(n334), .B(n333), .ZN(n354) );
  XOR2_X1 U382 ( .A(G64GAT), .B(KEYINPUT79), .Z(n336) );
  XNOR2_X1 U383 ( .A(G15GAT), .B(G71GAT), .ZN(n335) );
  XNOR2_X1 U384 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U385 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n338) );
  XNOR2_X1 U386 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U388 ( .A(n340), .B(n339), .Z(n352) );
  XNOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n341) );
  XNOR2_X1 U390 ( .A(n341), .B(KEYINPUT72), .ZN(n372) );
  XOR2_X1 U391 ( .A(n372), .B(KEYINPUT83), .Z(n343) );
  NAND2_X1 U392 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n350) );
  XOR2_X1 U394 ( .A(G78GAT), .B(G155GAT), .Z(n345) );
  XNOR2_X1 U395 ( .A(G127GAT), .B(G183GAT), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U397 ( .A(n346), .B(G211GAT), .Z(n348) );
  XOR2_X1 U398 ( .A(G1GAT), .B(KEYINPUT70), .Z(n361) );
  XNOR2_X1 U399 ( .A(G22GAT), .B(n361), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U402 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U403 ( .A(n354), .B(n353), .ZN(n580) );
  XOR2_X1 U404 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n360) );
  XOR2_X1 U405 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n356) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(KEYINPUT67), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n358) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(G15GAT), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n357), .B(G113GAT), .ZN(n448) );
  XNOR2_X1 U410 ( .A(n358), .B(n448), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n365) );
  XOR2_X1 U412 ( .A(G197GAT), .B(G8GAT), .Z(n433) );
  XOR2_X1 U413 ( .A(n433), .B(n361), .Z(n363) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U416 ( .A(n365), .B(n364), .Z(n371) );
  XOR2_X1 U417 ( .A(KEYINPUT7), .B(G50GAT), .Z(n367) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G29GAT), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U420 ( .A(KEYINPUT8), .B(n368), .Z(n403) );
  XNOR2_X1 U421 ( .A(n403), .B(n369), .ZN(n370) );
  XNOR2_X1 U422 ( .A(n371), .B(n370), .ZN(n573) );
  XNOR2_X1 U423 ( .A(n372), .B(n387), .ZN(n374) );
  NAND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U426 ( .A(G92GAT), .B(G64GAT), .Z(n425) );
  XNOR2_X1 U427 ( .A(n375), .B(n425), .ZN(n377) );
  XNOR2_X1 U428 ( .A(G176GAT), .B(G204GAT), .ZN(n376) );
  XNOR2_X1 U429 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U430 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n379) );
  XNOR2_X1 U431 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n378) );
  XOR2_X1 U432 ( .A(n379), .B(n378), .Z(n380) );
  XNOR2_X1 U433 ( .A(n381), .B(n380), .ZN(n385) );
  XNOR2_X1 U434 ( .A(G99GAT), .B(G71GAT), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n382), .B(G120GAT), .ZN(n442) );
  XNOR2_X1 U436 ( .A(n442), .B(n383), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n576) );
  XNOR2_X1 U438 ( .A(KEYINPUT41), .B(n576), .ZN(n554) );
  NAND2_X1 U439 ( .A1(n573), .A2(n554), .ZN(n386) );
  XNOR2_X1 U440 ( .A(KEYINPUT46), .B(n386), .ZN(n406) );
  XNOR2_X1 U441 ( .A(n387), .B(G162GAT), .ZN(n389) );
  XOR2_X1 U442 ( .A(G43GAT), .B(G218GAT), .Z(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U444 ( .A(G92GAT), .B(G106GAT), .Z(n391) );
  XNOR2_X1 U445 ( .A(G190GAT), .B(G99GAT), .ZN(n390) );
  XOR2_X1 U446 ( .A(n391), .B(n390), .Z(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n399) );
  XOR2_X1 U448 ( .A(KEYINPUT65), .B(KEYINPUT78), .Z(n395) );
  XNOR2_X1 U449 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n394) );
  XOR2_X1 U450 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U451 ( .A1(G232GAT), .A2(G233GAT), .ZN(n396) );
  XOR2_X1 U452 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n401) );
  XNOR2_X1 U453 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n400) );
  XNOR2_X1 U454 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U456 ( .A(n405), .B(n404), .ZN(n540) );
  NAND2_X1 U457 ( .A1(n406), .A2(n540), .ZN(n407) );
  NOR2_X1 U458 ( .A1(n580), .A2(n407), .ZN(n408) );
  XNOR2_X1 U459 ( .A(n409), .B(n408), .ZN(n418) );
  XOR2_X1 U460 ( .A(n573), .B(KEYINPUT71), .Z(n561) );
  INV_X1 U461 ( .A(KEYINPUT36), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n540), .B(n410), .ZN(n583) );
  NAND2_X1 U463 ( .A1(n583), .A2(n580), .ZN(n412) );
  XOR2_X1 U464 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n413) );
  NAND2_X1 U466 ( .A1(n576), .A2(n413), .ZN(n414) );
  XOR2_X1 U467 ( .A(KEYINPUT115), .B(n414), .Z(n415) );
  NOR2_X1 U468 ( .A1(n561), .A2(n415), .ZN(n416) );
  XNOR2_X1 U469 ( .A(KEYINPUT116), .B(n416), .ZN(n417) );
  NOR2_X1 U470 ( .A1(n418), .A2(n417), .ZN(n419) );
  XNOR2_X1 U471 ( .A(n419), .B(KEYINPUT48), .ZN(n544) );
  XOR2_X1 U472 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n421) );
  XNOR2_X1 U473 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n420) );
  XNOR2_X1 U474 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U475 ( .A(n422), .B(G183GAT), .Z(n424) );
  XNOR2_X1 U476 ( .A(G169GAT), .B(G176GAT), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n447) );
  XOR2_X1 U478 ( .A(KEYINPUT79), .B(n425), .Z(n427) );
  NAND2_X1 U479 ( .A1(G226GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U481 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n429) );
  XNOR2_X1 U482 ( .A(G36GAT), .B(KEYINPUT77), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U484 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U487 ( .A(n447), .B(n436), .Z(n510) );
  NOR2_X1 U488 ( .A1(n544), .A2(n510), .ZN(n437) );
  XNOR2_X1 U489 ( .A(KEYINPUT54), .B(n437), .ZN(n438) );
  AND2_X1 U490 ( .A1(n506), .A2(n438), .ZN(n572) );
  NAND2_X1 U491 ( .A1(n466), .A2(n572), .ZN(n439) );
  XNOR2_X1 U492 ( .A(KEYINPUT55), .B(n439), .ZN(n453) );
  XOR2_X1 U493 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n441) );
  XNOR2_X1 U494 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U496 ( .A(n442), .B(KEYINPUT87), .Z(n444) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U499 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U502 ( .A(n452), .B(n451), .Z(n512) );
  INV_X1 U503 ( .A(n512), .ZN(n532) );
  NAND2_X1 U504 ( .A1(n453), .A2(n532), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n566), .A2(n554), .ZN(n458) );
  XOR2_X1 U506 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n456) );
  XNOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n455) );
  NAND2_X1 U508 ( .A1(n540), .A2(n580), .ZN(n459) );
  XOR2_X1 U509 ( .A(KEYINPUT16), .B(n459), .Z(n474) );
  XNOR2_X1 U510 ( .A(n532), .B(KEYINPUT91), .ZN(n461) );
  XOR2_X1 U511 ( .A(n510), .B(KEYINPUT27), .Z(n464) );
  NAND2_X1 U512 ( .A1(n522), .A2(n464), .ZN(n547) );
  XOR2_X1 U513 ( .A(n466), .B(KEYINPUT66), .Z(n460) );
  XNOR2_X1 U514 ( .A(KEYINPUT28), .B(n460), .ZN(n528) );
  NOR2_X1 U515 ( .A1(n547), .A2(n528), .ZN(n531) );
  NAND2_X1 U516 ( .A1(n461), .A2(n531), .ZN(n473) );
  XNOR2_X1 U517 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n532), .A2(n466), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n463), .B(n462), .ZN(n571) );
  NAND2_X1 U520 ( .A1(n571), .A2(n464), .ZN(n469) );
  INV_X1 U521 ( .A(n510), .ZN(n524) );
  NAND2_X1 U522 ( .A1(n532), .A2(n524), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT25), .B(n467), .Z(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U526 ( .A1(n470), .A2(n506), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT101), .B(n471), .Z(n472) );
  NAND2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n487) );
  NAND2_X1 U529 ( .A1(n474), .A2(n487), .ZN(n504) );
  NAND2_X1 U530 ( .A1(n561), .A2(n576), .ZN(n490) );
  NOR2_X1 U531 ( .A1(n504), .A2(n490), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n475), .B(KEYINPUT102), .ZN(n485) );
  NAND2_X1 U533 ( .A1(n485), .A2(n522), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT34), .B(KEYINPUT104), .Z(n477) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(KEYINPUT103), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(G1324GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n481) );
  NAND2_X1 U539 ( .A1(n485), .A2(n524), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U543 ( .A1(n532), .A2(n485), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NAND2_X1 U545 ( .A1(n485), .A2(n528), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n493) );
  NAND2_X1 U548 ( .A1(n583), .A2(n487), .ZN(n488) );
  NOR2_X1 U549 ( .A1(n580), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT37), .B(n489), .ZN(n521) );
  NOR2_X1 U551 ( .A1(n521), .A2(n490), .ZN(n491) );
  XNOR2_X1 U552 ( .A(KEYINPUT38), .B(n491), .ZN(n501) );
  NAND2_X1 U553 ( .A1(n522), .A2(n501), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U555 ( .A(G29GAT), .B(n494), .Z(G1328GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n496) );
  NAND2_X1 U557 ( .A1(n501), .A2(n524), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n499) );
  NAND2_X1 U561 ( .A1(n532), .A2(n501), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U563 ( .A(G43GAT), .B(n500), .Z(G1330GAT) );
  NAND2_X1 U564 ( .A1(n501), .A2(n528), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U566 ( .A(n573), .ZN(n503) );
  NAND2_X1 U567 ( .A1(n503), .A2(n554), .ZN(n520) );
  NOR2_X1 U568 ( .A1(n520), .A2(n504), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT111), .ZN(n515) );
  NOR2_X1 U570 ( .A1(n506), .A2(n515), .ZN(n508) );
  XNOR2_X1 U571 ( .A(KEYINPUT42), .B(KEYINPUT112), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n509), .Z(G1332GAT) );
  NOR2_X1 U574 ( .A1(n510), .A2(n515), .ZN(n511) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n512), .A2(n515), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT113), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  INV_X1 U579 ( .A(n528), .ZN(n516) );
  NOR2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X1 U581 ( .A(KEYINPUT114), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n522), .A2(n527), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n524), .A2(n527), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n527), .A2(n532), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n529), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT117), .Z(n535) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U596 ( .A1(n544), .A2(n533), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n541), .A2(n561), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U600 ( .A1(n541), .A2(n554), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U602 ( .A1(n580), .A2(n541), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  INV_X1 U606 ( .A(n540), .ZN(n565) );
  NAND2_X1 U607 ( .A1(n541), .A2(n565), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n549) );
  INV_X1 U610 ( .A(n544), .ZN(n545) );
  NAND2_X1 U611 ( .A1(n545), .A2(n571), .ZN(n546) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n558), .A2(n573), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n552) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U619 ( .A(KEYINPUT120), .B(n553), .Z(n556) );
  NAND2_X1 U620 ( .A1(n558), .A2(n554), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n580), .A2(n558), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n565), .A2(n558), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT122), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n566), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT125), .Z(n564) );
  NAND2_X1 U630 ( .A1(n566), .A2(n580), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(KEYINPUT60), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT126), .B(n570), .Z(n575) );
  AND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U639 ( .A1(n584), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U642 ( .A(n576), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n584), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  XOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT127), .Z(n582) );
  NAND2_X1 U646 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1354GAT) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

