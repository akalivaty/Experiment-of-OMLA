

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786;

  XOR2_X1 U362 ( .A(G101), .B(KEYINPUT71), .Z(n340) );
  NOR2_X2 U363 ( .A1(n709), .A2(n708), .ZN(n647) );
  NAND2_X2 U364 ( .A1(n398), .A2(n397), .ZN(n455) );
  XNOR2_X2 U365 ( .A(n669), .B(n351), .ZN(n410) );
  NOR2_X2 U366 ( .A1(n619), .A2(n618), .ZN(n688) );
  NOR2_X2 U367 ( .A1(n656), .A2(n642), .ZN(n671) );
  XNOR2_X2 U368 ( .A(n440), .B(n439), .ZN(n786) );
  NAND2_X1 U369 ( .A1(n470), .A2(n473), .ZN(n716) );
  NOR2_X1 U370 ( .A1(n697), .A2(n615), .ZN(n598) );
  NOR2_X2 U371 ( .A1(n596), .A2(n708), .ZN(n643) );
  AND2_X1 U372 ( .A1(n358), .A2(n341), .ZN(n357) );
  AND2_X1 U373 ( .A1(n487), .A2(n485), .ZN(n484) );
  NAND2_X1 U374 ( .A1(n352), .A2(n438), .ZN(n669) );
  XNOR2_X1 U375 ( .A(n456), .B(n621), .ZN(n352) );
  AND2_X1 U376 ( .A1(n344), .A2(n343), .ZN(n623) );
  NAND2_X1 U377 ( .A1(n344), .A2(n688), .ZN(n599) );
  XNOR2_X1 U378 ( .A(n598), .B(n345), .ZN(n344) );
  NAND2_X1 U379 ( .A1(n342), .A2(n713), .ZN(n708) );
  INV_X1 U380 ( .A(n446), .ZN(n342) );
  BUF_X1 U381 ( .A(n659), .Z(n446) );
  AND2_X1 U382 ( .A1(n390), .A2(n592), .ZN(n358) );
  INV_X1 U383 ( .A(KEYINPUT86), .ZN(n351) );
  INV_X1 U384 ( .A(G953), .ZN(n776) );
  INV_X1 U385 ( .A(KEYINPUT39), .ZN(n345) );
  INV_X1 U386 ( .A(n383), .ZN(n341) );
  XNOR2_X1 U387 ( .A(n667), .B(n666), .ZN(n760) );
  NAND2_X1 U388 ( .A1(n484), .A2(n483), .ZN(n667) );
  AND2_X1 U389 ( .A1(n410), .A2(n668), .ZN(n409) );
  AND2_X1 U390 ( .A1(n486), .A2(n665), .ZN(n485) );
  AND2_X1 U391 ( .A1(n657), .A2(n658), .ZN(n440) );
  NOR2_X1 U392 ( .A1(n673), .A2(n691), .ZN(n649) );
  AND2_X1 U393 ( .A1(n510), .A2(n509), .ZN(n693) );
  NOR2_X1 U394 ( .A1(n685), .A2(n703), .ZN(n620) );
  XNOR2_X1 U395 ( .A(n599), .B(n600), .ZN(n783) );
  XNOR2_X1 U396 ( .A(n424), .B(n646), .ZN(n673) );
  XNOR2_X1 U397 ( .A(n365), .B(n364), .ZN(n645) );
  XNOR2_X1 U398 ( .A(n607), .B(n606), .ZN(n729) );
  AND2_X1 U399 ( .A1(n355), .A2(n353), .ZN(n361) );
  NOR2_X1 U400 ( .A1(n697), .A2(n605), .ZN(n607) );
  NAND2_X1 U401 ( .A1(n367), .A2(n366), .ZN(n365) );
  INV_X1 U402 ( .A(n622), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n495), .B(n341), .ZN(n367) );
  XNOR2_X1 U404 ( .A(n612), .B(n443), .ZN(n697) );
  AND2_X1 U405 ( .A1(n362), .A2(n383), .ZN(n360) );
  AND2_X1 U406 ( .A1(n467), .A2(n464), .ZN(n463) );
  AND2_X1 U407 ( .A1(n659), .A2(n475), .ZN(n561) );
  XOR2_X1 U408 ( .A(n740), .B(n739), .Z(n742) );
  OR2_X1 U409 ( .A1(n470), .A2(n468), .ZN(n467) );
  NAND2_X1 U410 ( .A1(n736), .A2(n356), .ZN(n362) );
  NAND2_X1 U411 ( .A1(n416), .A2(n358), .ZN(n363) );
  AND2_X1 U412 ( .A1(n385), .A2(n390), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n348), .B(n381), .ZN(n659) );
  NOR2_X2 U414 ( .A1(n471), .A2(n387), .ZN(n470) );
  INV_X1 U415 ( .A(n627), .ZN(n366) );
  XNOR2_X1 U416 ( .A(n346), .B(n560), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n437), .B(n523), .ZN(n430) );
  XNOR2_X1 U418 ( .A(n453), .B(n435), .ZN(n437) );
  XNOR2_X1 U419 ( .A(n516), .B(n515), .ZN(n435) );
  XNOR2_X1 U420 ( .A(n490), .B(n628), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n434), .B(G104), .ZN(n568) );
  INV_X1 U422 ( .A(KEYINPUT23), .ZN(n347) );
  NAND2_X1 U423 ( .A1(G234), .A2(G237), .ZN(n543) );
  XNOR2_X1 U424 ( .A(KEYINPUT80), .B(G110), .ZN(n481) );
  XOR2_X1 U425 ( .A(G902), .B(KEYINPUT15), .Z(n668) );
  XNOR2_X1 U426 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n433) );
  INV_X1 U427 ( .A(G122), .ZN(n434) );
  XNOR2_X1 U428 ( .A(KEYINPUT99), .B(KEYINPUT12), .ZN(n564) );
  NOR2_X1 U429 ( .A1(G953), .A2(G237), .ZN(n520) );
  BUF_X1 U430 ( .A(KEYINPUT95), .Z(n490) );
  INV_X2 U431 ( .A(G128), .ZN(n429) );
  XOR2_X1 U432 ( .A(G110), .B(G107), .Z(n533) );
  XNOR2_X1 U433 ( .A(n770), .B(n347), .ZN(n346) );
  NAND2_X1 U434 ( .A1(n350), .A2(n349), .ZN(n348) );
  INV_X1 U435 ( .A(n350), .ZN(n757) );
  INV_X1 U436 ( .A(G902), .ZN(n349) );
  INV_X1 U437 ( .A(n410), .ZN(n774) );
  NAND2_X1 U438 ( .A1(n354), .A2(n341), .ZN(n353) );
  INV_X1 U439 ( .A(n362), .ZN(n354) );
  NAND2_X1 U440 ( .A1(n357), .A2(n416), .ZN(n355) );
  AND2_X1 U441 ( .A1(n363), .A2(n362), .ZN(n495) );
  NAND2_X1 U442 ( .A1(n361), .A2(n359), .ZN(n371) );
  NAND2_X1 U443 ( .A1(n363), .A2(n360), .ZN(n359) );
  BUF_X1 U444 ( .A(n728), .Z(n368) );
  INV_X1 U445 ( .A(n641), .ZN(n369) );
  NAND2_X1 U446 ( .A1(n663), .A2(n370), .ZN(n486) );
  AND2_X1 U447 ( .A1(KEYINPUT44), .A2(KEYINPUT88), .ZN(n370) );
  XNOR2_X1 U448 ( .A(n497), .B(n496), .ZN(n782) );
  NOR2_X1 U449 ( .A1(n371), .A2(n627), .ZN(n372) );
  XNOR2_X1 U450 ( .A(n372), .B(n628), .ZN(n373) );
  XNOR2_X1 U451 ( .A(n637), .B(KEYINPUT35), .ZN(n374) );
  XNOR2_X1 U452 ( .A(n637), .B(KEYINPUT35), .ZN(n781) );
  NAND2_X1 U453 ( .A1(n409), .A2(n411), .ZN(n375) );
  NAND2_X1 U454 ( .A1(n409), .A2(n411), .ZN(n406) );
  XNOR2_X1 U455 ( .A(n432), .B(n431), .ZN(n453) );
  BUF_X1 U456 ( .A(n769), .Z(n376) );
  XNOR2_X1 U457 ( .A(n429), .B(G143), .ZN(n377) );
  NAND2_X1 U458 ( .A1(n398), .A2(n397), .ZN(n378) );
  INV_X1 U459 ( .A(n411), .ZN(n379) );
  INV_X1 U460 ( .A(n596), .ZN(n380) );
  NAND2_X1 U461 ( .A1(n405), .A2(KEYINPUT64), .ZN(n404) );
  NAND2_X1 U462 ( .A1(n396), .A2(n395), .ZN(n400) );
  OR2_X2 U463 ( .A1(n760), .A2(n441), .ZN(n732) );
  NAND2_X1 U464 ( .A1(n457), .A2(n505), .ZN(n456) );
  AND2_X1 U465 ( .A1(n507), .A2(n458), .ZN(n457) );
  XNOR2_X1 U466 ( .A(n448), .B(n506), .ZN(n505) );
  NOR2_X1 U467 ( .A1(n747), .A2(G902), .ZN(n538) );
  NOR2_X1 U468 ( .A1(n562), .A2(n472), .ZN(n471) );
  NAND2_X1 U469 ( .A1(n563), .A2(n349), .ZN(n472) );
  XNOR2_X1 U470 ( .A(n640), .B(n639), .ZN(n655) );
  INV_X1 U471 ( .A(KEYINPUT22), .ZN(n639) );
  NAND2_X1 U472 ( .A1(n604), .A2(n713), .ZN(n451) );
  NAND2_X1 U473 ( .A1(n404), .A2(n401), .ZN(n397) );
  NAND2_X1 U474 ( .A1(n400), .A2(n399), .ZN(n398) );
  XOR2_X1 U475 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n552) );
  XNOR2_X1 U476 ( .A(KEYINPUT4), .B(G131), .ZN(n522) );
  NAND2_X1 U477 ( .A1(n732), .A2(KEYINPUT64), .ZN(n395) );
  INV_X1 U478 ( .A(n406), .ZN(n396) );
  INV_X1 U479 ( .A(n732), .ZN(n405) );
  AND2_X1 U480 ( .A1(n482), .A2(n780), .ZN(n438) );
  XOR2_X1 U481 ( .A(KEYINPUT83), .B(KEYINPUT93), .Z(n532) );
  XNOR2_X1 U482 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n539) );
  NOR2_X1 U483 ( .A1(n462), .A2(n469), .ZN(n461) );
  INV_X1 U484 ( .A(n473), .ZN(n462) );
  NOR2_X1 U485 ( .A1(n466), .A2(n465), .ZN(n464) );
  NOR2_X1 U486 ( .A1(n700), .A2(n469), .ZN(n465) );
  INV_X1 U487 ( .A(n533), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n568), .B(n433), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n481), .B(KEYINPUT24), .ZN(n480) );
  XNOR2_X1 U490 ( .A(G119), .B(G128), .ZN(n479) );
  XNOR2_X1 U491 ( .A(n576), .B(n575), .ZN(n750) );
  XNOR2_X1 U492 ( .A(n574), .B(n512), .ZN(n575) );
  XNOR2_X1 U493 ( .A(KEYINPUT41), .B(KEYINPUT112), .ZN(n606) );
  NOR2_X1 U494 ( .A1(n626), .A2(n625), .ZN(n627) );
  INV_X1 U495 ( .A(KEYINPUT28), .ZN(n477) );
  XNOR2_X1 U496 ( .A(n586), .B(n449), .ZN(n618) );
  XNOR2_X1 U497 ( .A(KEYINPUT101), .B(G478), .ZN(n449) );
  XNOR2_X1 U498 ( .A(KEYINPUT6), .B(KEYINPUT103), .ZN(n511) );
  XNOR2_X1 U499 ( .A(n504), .B(n391), .ZN(n503) );
  INV_X1 U500 ( .A(n684), .ZN(n508) );
  INV_X1 U501 ( .A(KEYINPUT46), .ZN(n506) );
  AND2_X1 U502 ( .A1(n661), .A2(n662), .ZN(n488) );
  AND2_X1 U503 ( .A1(G953), .A2(G902), .ZN(n545) );
  INV_X1 U504 ( .A(KEYINPUT30), .ZN(n469) );
  NAND2_X1 U505 ( .A1(n700), .A2(n469), .ZN(n468) );
  NOR2_X1 U506 ( .A1(G237), .A2(G902), .ZN(n530) );
  XOR2_X1 U507 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n565) );
  XNOR2_X1 U508 ( .A(G113), .B(G143), .ZN(n572) );
  XOR2_X1 U509 ( .A(G140), .B(G131), .Z(n573) );
  XNOR2_X1 U510 ( .A(n526), .B(n525), .ZN(n528) );
  XNOR2_X1 U511 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n525) );
  NAND2_X1 U512 ( .A1(n403), .A2(KEYINPUT64), .ZN(n402) );
  INV_X1 U513 ( .A(n408), .ZN(n403) );
  XNOR2_X1 U514 ( .A(n593), .B(n444), .ZN(n443) );
  INV_X1 U515 ( .A(KEYINPUT38), .ZN(n444) );
  XNOR2_X1 U516 ( .A(n445), .B(KEYINPUT69), .ZN(n601) );
  INV_X1 U517 ( .A(n595), .ZN(n475) );
  NAND2_X1 U518 ( .A1(n418), .A2(n668), .ZN(n417) );
  XNOR2_X1 U519 ( .A(n521), .B(n519), .ZN(n500) );
  XNOR2_X1 U520 ( .A(n537), .B(n412), .ZN(n747) );
  XNOR2_X1 U521 ( .A(n415), .B(G101), .ZN(n412) );
  NAND2_X1 U522 ( .A1(n442), .A2(KEYINPUT2), .ZN(n441) );
  INV_X1 U523 ( .A(n669), .ZN(n442) );
  XNOR2_X1 U524 ( .A(KEYINPUT34), .B(KEYINPUT82), .ZN(n632) );
  XNOR2_X1 U525 ( .A(n559), .B(n513), .ZN(n560) );
  XNOR2_X1 U526 ( .A(n480), .B(n479), .ZN(n559) );
  XNOR2_X1 U527 ( .A(n584), .B(n450), .ZN(n752) );
  XNOR2_X1 U528 ( .A(n583), .B(n585), .ZN(n450) );
  XOR2_X1 U529 ( .A(G122), .B(KEYINPUT7), .Z(n585) );
  NAND2_X1 U530 ( .A1(n609), .A2(n608), .ZN(n610) );
  INV_X1 U531 ( .A(n654), .ZN(n509) );
  INV_X1 U532 ( .A(KEYINPUT32), .ZN(n439) );
  INV_X1 U533 ( .A(KEYINPUT105), .ZN(n496) );
  NAND2_X1 U534 ( .A1(n660), .A2(n498), .ZN(n497) );
  NOR2_X1 U535 ( .A1(n716), .A2(n342), .ZN(n498) );
  NAND2_X1 U536 ( .A1(n503), .A2(n502), .ZN(n501) );
  INV_X1 U537 ( .A(n436), .ZN(n766) );
  INV_X1 U538 ( .A(KEYINPUT60), .ZN(n491) );
  NAND2_X1 U539 ( .A1(n493), .A2(n502), .ZN(n492) );
  XNOR2_X1 U540 ( .A(n494), .B(n392), .ZN(n493) );
  XNOR2_X1 U541 ( .A(n420), .B(n419), .ZN(G75) );
  XNOR2_X1 U542 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n419) );
  NAND2_X1 U543 ( .A1(n734), .A2(n421), .ZN(n420) );
  AND2_X1 U544 ( .A1(n735), .A2(n776), .ZN(n421) );
  XOR2_X1 U545 ( .A(n552), .B(n551), .Z(n381) );
  XOR2_X1 U546 ( .A(KEYINPUT70), .B(G469), .Z(n382) );
  XNOR2_X1 U547 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n383) );
  AND2_X1 U548 ( .A1(n407), .A2(n414), .ZN(n384) );
  OR2_X1 U549 ( .A1(n418), .A2(n668), .ZN(n385) );
  AND2_X1 U550 ( .A1(n786), .A2(n782), .ZN(n386) );
  AND2_X1 U551 ( .A1(n474), .A2(G902), .ZN(n387) );
  NAND2_X1 U552 ( .A1(n588), .A2(G214), .ZN(n700) );
  AND2_X1 U553 ( .A1(n601), .A2(n688), .ZN(n388) );
  INV_X1 U554 ( .A(n482), .ZN(n696) );
  OR2_X1 U555 ( .A1(n644), .A2(n716), .ZN(n389) );
  AND2_X1 U556 ( .A1(n417), .A2(n700), .ZN(n390) );
  XOR2_X1 U557 ( .A(n562), .B(KEYINPUT62), .Z(n391) );
  XOR2_X1 U558 ( .A(n750), .B(n749), .Z(n392) );
  NAND2_X1 U559 ( .A1(n408), .A2(n413), .ZN(n393) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n413) );
  XOR2_X1 U561 ( .A(n670), .B(KEYINPUT92), .Z(n394) );
  NOR2_X1 U562 ( .A1(G952), .A2(n776), .ZN(n759) );
  INV_X1 U563 ( .A(n759), .ZN(n502) );
  NAND2_X1 U564 ( .A1(n375), .A2(n393), .ZN(n399) );
  NAND2_X1 U565 ( .A1(n732), .A2(n402), .ZN(n401) );
  NAND2_X1 U566 ( .A1(n411), .A2(n410), .ZN(n407) );
  NAND2_X1 U567 ( .A1(n668), .A2(KEYINPUT2), .ZN(n408) );
  INV_X1 U568 ( .A(n760), .ZN(n411) );
  XNOR2_X2 U569 ( .A(n769), .B(G146), .ZN(n415) );
  XNOR2_X2 U570 ( .A(n581), .B(n522), .ZN(n769) );
  INV_X1 U571 ( .A(KEYINPUT2), .ZN(n414) );
  XNOR2_X1 U572 ( .A(n499), .B(n415), .ZN(n562) );
  INV_X1 U573 ( .A(n736), .ZN(n416) );
  XNOR2_X2 U574 ( .A(n430), .B(n529), .ZN(n736) );
  INV_X1 U575 ( .A(n592), .ZN(n418) );
  BUF_X1 U576 ( .A(n378), .Z(n422) );
  NAND2_X1 U577 ( .A1(n736), .A2(n540), .ZN(n423) );
  NOR2_X1 U578 ( .A1(n645), .A2(n389), .ZN(n424) );
  BUF_X1 U579 ( .A(n747), .Z(n425) );
  BUF_X1 U580 ( .A(n581), .Z(n426) );
  NOR2_X2 U581 ( .A1(n655), .A2(n641), .ZN(n660) );
  XNOR2_X1 U582 ( .A(n631), .B(n630), .ZN(n728) );
  NOR2_X1 U583 ( .A1(n645), .A2(n728), .ZN(n633) );
  NOR2_X1 U584 ( .A1(n709), .A2(n708), .ZN(n427) );
  NAND2_X1 U585 ( .A1(n786), .A2(n782), .ZN(n663) );
  INV_X1 U586 ( .A(n612), .ZN(n428) );
  XNOR2_X1 U587 ( .A(n620), .B(KEYINPUT47), .ZN(n458) );
  XNOR2_X2 U588 ( .A(n429), .B(G143), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n435), .B(n500), .ZN(n499) );
  OR2_X1 U590 ( .A1(n437), .A2(n765), .ZN(n436) );
  NOR2_X1 U591 ( .A1(n655), .A2(n656), .ZN(n657) );
  NAND2_X1 U592 ( .A1(n656), .A2(n388), .ZN(n587) );
  NAND2_X1 U593 ( .A1(n663), .A2(KEYINPUT44), .ZN(n661) );
  OR2_X1 U594 ( .A1(n489), .A2(n662), .ZN(n483) );
  NAND2_X1 U595 ( .A1(n783), .A2(n784), .ZN(n448) );
  XNOR2_X1 U596 ( .A(n578), .B(n577), .ZN(n614) );
  INV_X1 U597 ( .A(n614), .ZN(n619) );
  NOR2_X1 U598 ( .A1(n373), .A2(n451), .ZN(n640) );
  XNOR2_X2 U599 ( .A(n602), .B(n539), .ZN(n709) );
  XNOR2_X2 U600 ( .A(n538), .B(n382), .ZN(n602) );
  NAND2_X1 U601 ( .A1(n561), .A2(n713), .ZN(n445) );
  INV_X1 U602 ( .A(n447), .ZN(n567) );
  XNOR2_X1 U603 ( .A(n553), .B(n554), .ZN(n447) );
  XNOR2_X2 U604 ( .A(G146), .B(G125), .ZN(n553) );
  XNOR2_X1 U605 ( .A(n478), .B(n477), .ZN(n476) );
  INV_X1 U606 ( .A(n729), .ZN(n608) );
  XNOR2_X1 U607 ( .A(n653), .B(KEYINPUT89), .ZN(n489) );
  XNOR2_X1 U608 ( .A(n745), .B(n452), .ZN(n748) );
  XNOR2_X1 U609 ( .A(n425), .B(n746), .ZN(n452) );
  XNOR2_X1 U610 ( .A(n454), .B(KEYINPUT124), .ZN(G63) );
  NOR2_X2 U611 ( .A1(n755), .A2(n759), .ZN(n454) );
  NAND2_X1 U612 ( .A1(n455), .A2(G478), .ZN(n754) );
  NAND2_X1 U613 ( .A1(n455), .A2(G210), .ZN(n741) );
  NAND2_X1 U614 ( .A1(n422), .A2(G469), .ZN(n745) );
  NAND2_X1 U615 ( .A1(n378), .A2(G475), .ZN(n494) );
  NAND2_X1 U616 ( .A1(n378), .A2(G472), .ZN(n504) );
  NAND2_X1 U617 ( .A1(n422), .A2(G217), .ZN(n756) );
  NAND2_X1 U618 ( .A1(n562), .A2(n474), .ZN(n473) );
  AND2_X1 U619 ( .A1(n562), .A2(n459), .ZN(n466) );
  NOR2_X1 U620 ( .A1(n468), .A2(n563), .ZN(n459) );
  NAND2_X1 U621 ( .A1(n463), .A2(n460), .ZN(n594) );
  NAND2_X1 U622 ( .A1(n470), .A2(n461), .ZN(n460) );
  INV_X1 U623 ( .A(n563), .ZN(n474) );
  NAND2_X1 U624 ( .A1(n476), .A2(n380), .ZN(n603) );
  NAND2_X1 U625 ( .A1(n601), .A2(n716), .ZN(n478) );
  NAND2_X1 U626 ( .A1(n616), .A2(n428), .ZN(n684) );
  OR2_X1 U627 ( .A1(n591), .A2(n428), .ZN(n482) );
  NAND2_X1 U628 ( .A1(n489), .A2(n488), .ZN(n487) );
  XNOR2_X1 U629 ( .A(n492), .B(n491), .ZN(G60) );
  XNOR2_X2 U630 ( .A(n524), .B(G134), .ZN(n581) );
  XNOR2_X1 U631 ( .A(n501), .B(n394), .ZN(G57) );
  NOR2_X1 U632 ( .A1(n693), .A2(n508), .ZN(n507) );
  XNOR2_X1 U633 ( .A(n613), .B(KEYINPUT36), .ZN(n510) );
  XNOR2_X2 U634 ( .A(n716), .B(n511), .ZN(n656) );
  NOR2_X2 U635 ( .A1(n743), .A2(n759), .ZN(n744) );
  XNOR2_X1 U636 ( .A(n754), .B(n753), .ZN(n755) );
  XOR2_X1 U637 ( .A(n573), .B(n572), .Z(n512) );
  AND2_X1 U638 ( .A1(n582), .A2(G221), .ZN(n513) );
  INV_X1 U639 ( .A(KEYINPUT48), .ZN(n621) );
  INV_X1 U640 ( .A(KEYINPUT88), .ZN(n662) );
  XNOR2_X1 U641 ( .A(n629), .B(KEYINPUT33), .ZN(n630) );
  INV_X1 U642 ( .A(n555), .ZN(n556) );
  XNOR2_X1 U643 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U644 ( .A(n610), .B(KEYINPUT42), .ZN(n784) );
  XNOR2_X1 U645 ( .A(G116), .B(G113), .ZN(n514) );
  XNOR2_X1 U646 ( .A(n340), .B(n514), .ZN(n516) );
  XOR2_X1 U647 ( .A(G119), .B(KEYINPUT3), .Z(n515) );
  XOR2_X1 U648 ( .A(KEYINPUT5), .B(KEYINPUT77), .Z(n518) );
  XNOR2_X1 U649 ( .A(G137), .B(KEYINPUT78), .ZN(n517) );
  XNOR2_X1 U650 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U651 ( .A(KEYINPUT79), .B(n520), .Z(n571) );
  NAND2_X1 U652 ( .A1(G210), .A2(n571), .ZN(n521) );
  INV_X1 U653 ( .A(n668), .ZN(n540) );
  INV_X1 U654 ( .A(KEYINPUT18), .ZN(n523) );
  XOR2_X1 U655 ( .A(n377), .B(n553), .Z(n526) );
  NAND2_X1 U656 ( .A1(G224), .A2(n776), .ZN(n527) );
  XOR2_X1 U657 ( .A(KEYINPUT76), .B(n530), .Z(n588) );
  NAND2_X1 U658 ( .A1(n588), .A2(G210), .ZN(n531) );
  XNOR2_X1 U659 ( .A(n532), .B(n531), .ZN(n592) );
  XOR2_X1 U660 ( .A(G137), .B(G140), .Z(n555) );
  XOR2_X1 U661 ( .A(n533), .B(n555), .Z(n535) );
  NAND2_X1 U662 ( .A1(G227), .A2(n776), .ZN(n534) );
  XNOR2_X1 U663 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U664 ( .A(n536), .B(G104), .Z(n537) );
  INV_X1 U665 ( .A(n709), .ZN(n641) );
  NAND2_X1 U666 ( .A1(G234), .A2(n540), .ZN(n541) );
  XNOR2_X1 U667 ( .A(KEYINPUT20), .B(n541), .ZN(n550) );
  NAND2_X1 U668 ( .A1(n550), .A2(G221), .ZN(n542) );
  XNOR2_X1 U669 ( .A(KEYINPUT21), .B(n542), .ZN(n638) );
  INV_X1 U670 ( .A(n638), .ZN(n713) );
  XNOR2_X1 U671 ( .A(n543), .B(KEYINPUT14), .ZN(n546) );
  NAND2_X1 U672 ( .A1(n546), .A2(G952), .ZN(n544) );
  XNOR2_X1 U673 ( .A(n544), .B(KEYINPUT94), .ZN(n727) );
  NOR2_X1 U674 ( .A1(G953), .A2(n727), .ZN(n626) );
  NAND2_X1 U675 ( .A1(n546), .A2(n545), .ZN(n624) );
  XOR2_X1 U676 ( .A(KEYINPUT107), .B(n624), .Z(n547) );
  NOR2_X1 U677 ( .A1(G900), .A2(n547), .ZN(n548) );
  XNOR2_X1 U678 ( .A(n548), .B(KEYINPUT108), .ZN(n549) );
  NOR2_X1 U679 ( .A1(n626), .A2(n549), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n550), .A2(G217), .ZN(n551) );
  XNOR2_X1 U681 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n554) );
  XNOR2_X2 U682 ( .A(n567), .B(n556), .ZN(n770) );
  NAND2_X1 U683 ( .A1(n776), .A2(G234), .ZN(n558) );
  XNOR2_X1 U684 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n557) );
  XNOR2_X1 U685 ( .A(n558), .B(n557), .ZN(n582) );
  XNOR2_X1 U686 ( .A(G472), .B(KEYINPUT73), .ZN(n563) );
  XNOR2_X1 U687 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U688 ( .A(KEYINPUT100), .B(n566), .Z(n570) );
  XOR2_X1 U689 ( .A(n568), .B(n447), .Z(n569) );
  XNOR2_X1 U690 ( .A(n570), .B(n569), .ZN(n576) );
  NAND2_X1 U691 ( .A1(G214), .A2(n571), .ZN(n574) );
  NOR2_X1 U692 ( .A1(G902), .A2(n750), .ZN(n578) );
  XNOR2_X1 U693 ( .A(KEYINPUT13), .B(G475), .ZN(n577) );
  XNOR2_X1 U694 ( .A(G116), .B(G107), .ZN(n579) );
  XNOR2_X1 U695 ( .A(n579), .B(KEYINPUT9), .ZN(n580) );
  XNOR2_X1 U696 ( .A(n426), .B(n580), .ZN(n584) );
  NAND2_X1 U697 ( .A1(n582), .A2(G217), .ZN(n583) );
  NOR2_X1 U698 ( .A1(G902), .A2(n752), .ZN(n586) );
  XNOR2_X1 U699 ( .A(n587), .B(KEYINPUT109), .ZN(n589) );
  NAND2_X1 U700 ( .A1(n589), .A2(n700), .ZN(n611) );
  NOR2_X1 U701 ( .A1(n641), .A2(n611), .ZN(n590) );
  XNOR2_X1 U702 ( .A(n590), .B(KEYINPUT43), .ZN(n591) );
  XOR2_X1 U703 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n600) );
  INV_X1 U704 ( .A(n688), .ZN(n686) );
  XOR2_X1 U705 ( .A(n423), .B(n592), .Z(n612) );
  INV_X1 U706 ( .A(KEYINPUT75), .ZN(n593) );
  NOR2_X1 U707 ( .A1(n595), .A2(n594), .ZN(n597) );
  INV_X1 U708 ( .A(n602), .ZN(n596) );
  NAND2_X1 U709 ( .A1(n597), .A2(n643), .ZN(n615) );
  XNOR2_X1 U710 ( .A(KEYINPUT110), .B(n603), .ZN(n617) );
  INV_X1 U711 ( .A(n617), .ZN(n609) );
  OR2_X1 U712 ( .A1(n618), .A2(n614), .ZN(n699) );
  INV_X1 U713 ( .A(n699), .ZN(n604) );
  NAND2_X1 U714 ( .A1(n700), .A2(n604), .ZN(n605) );
  XOR2_X1 U715 ( .A(n709), .B(KEYINPUT91), .Z(n654) );
  NOR2_X1 U716 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U717 ( .A1(n618), .A2(n614), .ZN(n634) );
  NOR2_X1 U718 ( .A1(n615), .A2(n634), .ZN(n616) );
  OR2_X1 U719 ( .A1(n617), .A2(n371), .ZN(n685) );
  NAND2_X1 U720 ( .A1(n619), .A2(n618), .ZN(n680) );
  XNOR2_X1 U721 ( .A(KEYINPUT102), .B(n680), .ZN(n622) );
  AND2_X1 U722 ( .A1(n686), .A2(n622), .ZN(n703) );
  XNOR2_X1 U723 ( .A(n623), .B(KEYINPUT113), .ZN(n780) );
  NOR2_X1 U724 ( .A1(G898), .A2(n624), .ZN(n625) );
  INV_X1 U725 ( .A(KEYINPUT0), .ZN(n628) );
  NAND2_X1 U726 ( .A1(n647), .A2(n656), .ZN(n631) );
  XOR2_X1 U727 ( .A(KEYINPUT72), .B(KEYINPUT106), .Z(n629) );
  XNOR2_X1 U728 ( .A(n633), .B(n632), .ZN(n636) );
  XNOR2_X1 U729 ( .A(n634), .B(KEYINPUT81), .ZN(n635) );
  NAND2_X1 U730 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U731 ( .A1(n781), .A2(KEYINPUT44), .ZN(n652) );
  XOR2_X1 U732 ( .A(n446), .B(KEYINPUT104), .Z(n712) );
  NAND2_X1 U733 ( .A1(n660), .A2(n712), .ZN(n642) );
  INV_X1 U734 ( .A(n643), .ZN(n644) );
  INV_X1 U735 ( .A(KEYINPUT97), .ZN(n646) );
  NAND2_X1 U736 ( .A1(n716), .A2(n427), .ZN(n719) );
  NOR2_X1 U737 ( .A1(n373), .A2(n719), .ZN(n648) );
  XOR2_X1 U738 ( .A(KEYINPUT31), .B(n648), .Z(n691) );
  NOR2_X1 U739 ( .A1(n649), .A2(n703), .ZN(n650) );
  NOR2_X1 U740 ( .A1(n671), .A2(n650), .ZN(n651) );
  NAND2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U742 ( .A1(n654), .A2(n712), .ZN(n658) );
  NOR2_X1 U743 ( .A1(n374), .A2(KEYINPUT44), .ZN(n664) );
  NAND2_X1 U744 ( .A1(n386), .A2(n664), .ZN(n665) );
  XNOR2_X1 U745 ( .A(KEYINPUT87), .B(KEYINPUT45), .ZN(n666) );
  INV_X1 U746 ( .A(KEYINPUT63), .ZN(n670) );
  XOR2_X1 U747 ( .A(G101), .B(n671), .Z(G3) );
  NAND2_X1 U748 ( .A1(n673), .A2(n688), .ZN(n672) );
  XNOR2_X1 U749 ( .A(n672), .B(G104), .ZN(G6) );
  INV_X1 U750 ( .A(n680), .ZN(n690) );
  NAND2_X1 U751 ( .A1(n673), .A2(n690), .ZN(n679) );
  XOR2_X1 U752 ( .A(KEYINPUT116), .B(KEYINPUT27), .Z(n675) );
  XNOR2_X1 U753 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n674) );
  XNOR2_X1 U754 ( .A(n675), .B(n674), .ZN(n677) );
  XOR2_X1 U755 ( .A(G107), .B(KEYINPUT26), .Z(n676) );
  XNOR2_X1 U756 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U757 ( .A(n679), .B(n678), .ZN(G9) );
  NOR2_X1 U758 ( .A1(n680), .A2(n685), .ZN(n682) );
  XNOR2_X1 U759 ( .A(KEYINPUT117), .B(KEYINPUT29), .ZN(n681) );
  XNOR2_X1 U760 ( .A(n682), .B(n681), .ZN(n683) );
  XOR2_X1 U761 ( .A(G128), .B(n683), .Z(G30) );
  XNOR2_X1 U762 ( .A(G143), .B(n684), .ZN(G45) );
  NOR2_X1 U763 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U764 ( .A(G146), .B(n687), .Z(G48) );
  NAND2_X1 U765 ( .A1(n691), .A2(n688), .ZN(n689) );
  XNOR2_X1 U766 ( .A(n689), .B(G113), .ZN(G15) );
  NAND2_X1 U767 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U768 ( .A(n692), .B(G116), .ZN(G18) );
  XNOR2_X1 U769 ( .A(n693), .B(KEYINPUT37), .ZN(n694) );
  XNOR2_X1 U770 ( .A(n694), .B(KEYINPUT118), .ZN(n695) );
  XNOR2_X1 U771 ( .A(G125), .B(n695), .ZN(G27) );
  XOR2_X1 U772 ( .A(G140), .B(n696), .Z(G42) );
  INV_X1 U773 ( .A(n697), .ZN(n701) );
  NOR2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n698) );
  NOR2_X1 U775 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U777 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U778 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U779 ( .A(n706), .B(KEYINPUT120), .ZN(n707) );
  NOR2_X1 U780 ( .A1(n368), .A2(n707), .ZN(n724) );
  NAND2_X1 U781 ( .A1(n369), .A2(n708), .ZN(n710) );
  XOR2_X1 U782 ( .A(KEYINPUT50), .B(n710), .Z(n711) );
  XNOR2_X1 U783 ( .A(n711), .B(KEYINPUT119), .ZN(n718) );
  NOR2_X1 U784 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U785 ( .A(KEYINPUT49), .B(n714), .Z(n715) );
  NOR2_X1 U786 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U789 ( .A(KEYINPUT51), .B(n721), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n729), .A2(n722), .ZN(n723) );
  NOR2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U792 ( .A(n725), .B(KEYINPUT52), .ZN(n726) );
  NOR2_X1 U793 ( .A1(n727), .A2(n726), .ZN(n731) );
  NOR2_X1 U794 ( .A1(n729), .A2(n368), .ZN(n730) );
  NOR2_X1 U795 ( .A1(n731), .A2(n730), .ZN(n735) );
  XOR2_X1 U796 ( .A(n384), .B(KEYINPUT84), .Z(n733) );
  NAND2_X1 U797 ( .A1(n733), .A2(n732), .ZN(n734) );
  BUF_X1 U798 ( .A(n736), .Z(n740) );
  XOR2_X1 U799 ( .A(KEYINPUT55), .B(KEYINPUT90), .Z(n738) );
  XNOR2_X1 U800 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n737) );
  XNOR2_X1 U801 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U802 ( .A(n741), .B(n742), .ZN(n743) );
  XNOR2_X1 U803 ( .A(n744), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U804 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n746) );
  NOR2_X1 U805 ( .A1(n759), .A2(n748), .ZN(G54) );
  XOR2_X1 U806 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n749) );
  INV_X1 U807 ( .A(KEYINPUT123), .ZN(n751) );
  XNOR2_X1 U808 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U809 ( .A(n757), .B(n756), .ZN(n758) );
  NOR2_X1 U810 ( .A1(n759), .A2(n758), .ZN(G66) );
  OR2_X1 U811 ( .A1(G953), .A2(n379), .ZN(n764) );
  NAND2_X1 U812 ( .A1(G953), .A2(G224), .ZN(n761) );
  XNOR2_X1 U813 ( .A(KEYINPUT61), .B(n761), .ZN(n762) );
  NAND2_X1 U814 ( .A1(n762), .A2(G898), .ZN(n763) );
  NAND2_X1 U815 ( .A1(n764), .A2(n763), .ZN(n767) );
  NOR2_X1 U816 ( .A1(G898), .A2(n776), .ZN(n765) );
  XNOR2_X1 U817 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U818 ( .A(KEYINPUT125), .B(n768), .Z(G69) );
  XOR2_X1 U819 ( .A(n376), .B(n770), .Z(n775) );
  XNOR2_X1 U820 ( .A(G227), .B(n775), .ZN(n771) );
  NAND2_X1 U821 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U822 ( .A1(G953), .A2(n772), .ZN(n773) );
  XNOR2_X1 U823 ( .A(n773), .B(KEYINPUT126), .ZN(n779) );
  XNOR2_X1 U824 ( .A(n775), .B(n774), .ZN(n777) );
  NAND2_X1 U825 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U826 ( .A1(n779), .A2(n778), .ZN(G72) );
  XNOR2_X1 U827 ( .A(G134), .B(n780), .ZN(G36) );
  XOR2_X1 U828 ( .A(n374), .B(G122), .Z(G24) );
  XNOR2_X1 U829 ( .A(n782), .B(G110), .ZN(G12) );
  XNOR2_X1 U830 ( .A(G131), .B(n783), .ZN(G33) );
  XOR2_X1 U831 ( .A(n784), .B(G137), .Z(n785) );
  XNOR2_X1 U832 ( .A(KEYINPUT127), .B(n785), .ZN(G39) );
  XNOR2_X1 U833 ( .A(n786), .B(G119), .ZN(G21) );
endmodule

