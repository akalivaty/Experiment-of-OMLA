//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT64), .Z(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n459), .A2(G2104), .ZN(new_n469));
  OAI22_X1  g044(.A1(new_n466), .A2(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT65), .Z(G160));
  INV_X1    g047(.A(new_n466), .ZN(new_n473));
  MUX2_X1   g048(.A(G100), .B(G112), .S(G2105), .Z(new_n474));
  AOI22_X1  g049(.A1(new_n473), .A2(G136), .B1(G2104), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n460), .ZN(new_n476));
  OR3_X1    g051(.A1(new_n476), .A2(KEYINPUT66), .A3(new_n459), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT66), .B1(new_n476), .B2(new_n459), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT67), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G138), .B1(new_n484), .B2(KEYINPUT67), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n466), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G102), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2104), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n460), .A2(new_n496), .A3(new_n459), .A4(new_n485), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n488), .A2(new_n489), .A3(new_n493), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n507), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n504), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n502), .A2(KEYINPUT68), .A3(new_n503), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  INV_X1    g100(.A(new_n511), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT69), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(KEYINPUT69), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n502), .A2(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n530), .A2(G89), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n506), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n511), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n514), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(new_n523), .A2(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n506), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n511), .A2(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n514), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n530), .A2(G91), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n511), .A2(G53), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n556), .B1(new_n506), .B2(new_n557), .C1(new_n559), .C2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  OAI21_X1  g137(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n564));
  INV_X1    g139(.A(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n514), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n530), .A2(KEYINPUT70), .A3(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n511), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(new_n511), .A2(G48), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n514), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n506), .ZN(new_n576));
  AND2_X1   g151(.A1(KEYINPUT5), .A2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(KEYINPUT5), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G61), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(KEYINPUT71), .A3(G651), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n573), .B1(new_n576), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n506), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n530), .A2(G85), .B1(new_n511), .B2(G47), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G290));
  NAND3_X1  g163(.A1(G301), .A2(KEYINPUT72), .A3(G868), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n590));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(G171), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n511), .A2(G54), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n506), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT73), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n530), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n589), .B(new_n592), .C1(new_n600), .C2(G868), .ZN(G284));
  OAI211_X1 g176(.A(new_n589), .B(new_n592), .C1(new_n600), .C2(G868), .ZN(G321));
  NOR2_X1   g177(.A1(G299), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g179(.A(new_n603), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G860), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n599), .B1(G559), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT74), .ZN(G148));
  OR2_X1    g183(.A1(new_n599), .A2(G559), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(new_n591), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n549), .A2(new_n591), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(G282));
  INV_X1    g189(.A(new_n612), .ZN(G323));
  NAND2_X1  g190(.A1(new_n473), .A2(G2104), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT13), .Z(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2100), .ZN(new_n621));
  MUX2_X1   g196(.A(G99), .B(G111), .S(G2105), .Z(new_n622));
  AOI22_X1  g197(.A1(new_n473), .A2(G135), .B1(G2104), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G123), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n480), .B2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2096), .Z(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(G156));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT78), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT77), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n632), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT76), .B(KEYINPUT14), .Z(new_n635));
  NAND3_X1  g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT80), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n648), .B(KEYINPUT17), .Z(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n654), .C1(new_n651), .C2(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n651), .A3(new_n653), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n650), .A3(new_n648), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT81), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n668), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT20), .Z(new_n672));
  AOI211_X1 g247(.A(new_n670), .B(new_n672), .C1(new_n665), .C2(new_n669), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G229));
  XOR2_X1   g254(.A(KEYINPUT31), .B(G11), .Z(new_n680));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT30), .B(G28), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n625), .B2(new_n681), .ZN(new_n684));
  INV_X1    g259(.A(G103), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n469), .A2(KEYINPUT25), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(KEYINPUT25), .B1(new_n469), .B2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G139), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n686), .B(new_n687), .C1(new_n688), .C2(new_n466), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT90), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n460), .A2(G127), .ZN(new_n691));
  AND2_X1   g266(.A1(G115), .A2(G2104), .ZN(new_n692));
  OAI21_X1  g267(.A(G2105), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G29), .ZN(new_n695));
  NOR2_X1   g270(.A1(G29), .A2(G33), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT89), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(G2072), .Z(new_n699));
  INV_X1    g274(.A(G2084), .ZN(new_n700));
  INV_X1    g275(.A(G34), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(KEYINPUT24), .ZN(new_n702));
  AOI21_X1  g277(.A(G29), .B1(new_n701), .B2(KEYINPUT24), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(KEYINPUT91), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(KEYINPUT91), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G160), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n681), .ZN(new_n707));
  AOI211_X1 g282(.A(new_n684), .B(new_n699), .C1(new_n700), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n681), .A2(G32), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n473), .A2(G141), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT26), .Z(new_n712));
  INV_X1    g287(.A(G105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n710), .B(new_n712), .C1(new_n713), .C2(new_n469), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n479), .B2(G129), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n709), .B1(new_n715), .B2(new_n681), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT27), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n707), .A2(new_n700), .ZN(new_n720));
  NOR2_X1   g295(.A1(G27), .A2(G29), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G164), .B2(G29), .ZN(new_n722));
  INV_X1    g297(.A(G2078), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n708), .A2(new_n719), .A3(new_n720), .A4(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n726), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1961), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(G21), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G168), .B2(new_n726), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1966), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n725), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT93), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n479), .A2(G119), .ZN(new_n735));
  MUX2_X1   g310(.A(G95), .B(G107), .S(G2105), .Z(new_n736));
  AOI22_X1  g311(.A1(new_n473), .A2(G131), .B1(G2104), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G25), .B(new_n738), .S(G29), .Z(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n726), .A2(G24), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT82), .ZN(new_n743));
  INV_X1    g318(.A(G290), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n726), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n741), .B1(G1986), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G1986), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n726), .A2(G23), .ZN(new_n748));
  INV_X1    g323(.A(G288), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n726), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT33), .B(G1976), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G6), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n583), .B2(G16), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT32), .B(G1981), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G16), .A2(G22), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G166), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1971), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n752), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n747), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(KEYINPUT84), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT95), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n726), .A2(G20), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT23), .Z(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT96), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n774), .B2(new_n773), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n681), .A2(G26), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT28), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n473), .A2(G140), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G104), .B(G116), .S(G2105), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G2104), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT86), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n786), .B(new_n789), .C1(new_n479), .C2(G128), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT87), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n784), .B1(new_n791), .B2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2067), .ZN(new_n793));
  NOR2_X1   g368(.A1(G4), .A2(G16), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n600), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1348), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n726), .A2(G19), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT85), .Z(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n549), .B2(new_n726), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1341), .Z(new_n800));
  NAND3_X1  g375(.A1(new_n793), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n776), .B(new_n782), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n734), .A2(new_n769), .A3(new_n804), .ZN(G150));
  INV_X1    g380(.A(G150), .ZN(G311));
  AOI22_X1  g381(.A1(new_n530), .A2(G93), .B1(new_n511), .B2(G55), .ZN(new_n807));
  NAND2_X1  g382(.A1(G80), .A2(G543), .ZN(new_n808));
  INV_X1    g383(.A(G67), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n522), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n810), .A2(KEYINPUT97), .A3(G651), .ZN(new_n811));
  AOI21_X1  g386(.A(KEYINPUT97), .B1(new_n810), .B2(G651), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n807), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT37), .Z(new_n815));
  INV_X1    g390(.A(new_n549), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n813), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT38), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n600), .A2(G559), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT98), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n606), .B1(new_n824), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n815), .B1(new_n825), .B2(new_n826), .ZN(G145));
  AND2_X1   g402(.A1(new_n488), .A2(new_n497), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n493), .A2(new_n489), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n493), .A2(new_n489), .A3(KEYINPUT100), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n828), .A2(new_n829), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n833), .A2(new_n488), .A3(new_n497), .ZN(new_n835));
  AOI21_X1  g410(.A(KEYINPUT100), .B1(new_n493), .B2(new_n489), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT101), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n791), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n738), .B(new_n617), .ZN(new_n841));
  INV_X1    g416(.A(G118), .ZN(new_n842));
  AOI21_X1  g417(.A(KEYINPUT103), .B1(new_n842), .B2(G2105), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n842), .A2(KEYINPUT103), .A3(G2105), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n473), .A2(G142), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G130), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n480), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n841), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n840), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n852));
  INV_X1    g427(.A(new_n715), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n840), .A2(new_n850), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n851), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n854), .B1(new_n851), .B2(new_n855), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(G160), .B(new_n482), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n625), .B(KEYINPUT99), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n859), .B(new_n860), .Z(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n861), .B1(new_n856), .B2(new_n857), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(G395));
  XNOR2_X1  g443(.A(new_n819), .B(new_n609), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n599), .A2(G299), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n599), .A2(G299), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n873), .B1(new_n877), .B2(new_n869), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT42), .ZN(new_n879));
  XNOR2_X1  g454(.A(G290), .B(G288), .ZN(new_n880));
  XOR2_X1   g455(.A(G303), .B(new_n583), .Z(new_n881));
  XOR2_X1   g456(.A(new_n880), .B(new_n881), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n879), .B(new_n882), .ZN(new_n883));
  MUX2_X1   g458(.A(new_n813), .B(new_n883), .S(G868), .Z(G295));
  MUX2_X1   g459(.A(new_n813), .B(new_n883), .S(G868), .Z(G331));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  NAND2_X1  g461(.A1(G286), .A2(G301), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n528), .A2(G171), .A3(new_n529), .A4(new_n534), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n889), .B2(new_n819), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n819), .B2(new_n889), .ZN(new_n891));
  OR3_X1    g466(.A1(new_n889), .A2(new_n819), .A3(KEYINPUT106), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n872), .ZN(new_n894));
  INV_X1    g469(.A(new_n882), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n889), .B(new_n819), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n896), .A2(KEYINPUT105), .A3(new_n876), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT105), .B1(new_n896), .B2(new_n876), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n894), .B(new_n895), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n872), .ZN(new_n900));
  OAI22_X1  g475(.A1(new_n893), .A2(new_n877), .B1(new_n900), .B2(new_n896), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n882), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n902), .A3(new_n864), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT43), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n882), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n864), .A4(new_n899), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n904), .A2(new_n908), .A3(KEYINPUT44), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n903), .A2(new_n907), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n906), .A2(KEYINPUT43), .A3(new_n864), .A4(new_n899), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI22_X1  g490(.A1(new_n911), .A2(new_n912), .B1(KEYINPUT44), .B2(new_n915), .ZN(G397));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n838), .B2(G1384), .ZN(new_n918));
  INV_X1    g493(.A(G40), .ZN(new_n919));
  OR3_X1    g494(.A1(new_n463), .A2(new_n919), .A3(new_n470), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n791), .B(G2067), .ZN(new_n922));
  INV_X1    g497(.A(G1996), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n715), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n740), .B1(new_n735), .B2(new_n737), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n735), .A2(new_n737), .A3(new_n740), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n921), .A2(new_n923), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n715), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n921), .ZN(new_n933));
  NOR2_X1   g508(.A1(G290), .A2(G1986), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT108), .ZN(new_n935));
  NAND2_X1  g510(.A1(G290), .A2(G1986), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT124), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n835), .B2(new_n836), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n917), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n463), .A2(new_n919), .A3(new_n470), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT114), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n920), .B1(new_n943), .B2(new_n917), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT114), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT115), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n498), .A2(new_n953), .A3(KEYINPUT45), .A4(new_n942), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n947), .A2(new_n723), .A3(new_n950), .A4(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT121), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n941), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n958), .B2(new_n957), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n961));
  NAND4_X1  g536(.A1(new_n834), .A2(new_n837), .A3(KEYINPUT45), .A4(new_n942), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n498), .A2(new_n942), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n920), .B1(new_n917), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n961), .B1(new_n965), .B2(G2078), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n832), .A2(new_n488), .A3(new_n497), .A4(new_n833), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT50), .B1(new_n967), .B2(new_n942), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n498), .A2(KEYINPUT50), .A3(new_n942), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n945), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1961), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G301), .B1(new_n960), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(G8), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n967), .A2(KEYINPUT50), .A3(new_n942), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n963), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n920), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n965), .A2(new_n759), .B1(new_n981), .B2(new_n774), .ZN(new_n982));
  INV_X1    g557(.A(G8), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n977), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n967), .A2(new_n945), .A3(new_n942), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n985), .B(G8), .C1(G288), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT52), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n749), .B2(G1976), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n530), .A2(G86), .B1(new_n511), .B2(G48), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT111), .B(G1981), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT71), .B1(new_n581), .B2(G651), .ZN(new_n995));
  AOI211_X1 g570(.A(new_n574), .B(new_n506), .C1(new_n579), .C2(new_n580), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n993), .B(new_n994), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1981), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n583), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n985), .A2(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1001), .B1(new_n999), .B2(new_n1000), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n992), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n999), .A2(new_n1000), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT49), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1008), .A2(KEYINPUT113), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n991), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n965), .A2(new_n759), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n943), .A2(new_n979), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n920), .B1(new_n1012), .B2(new_n969), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n774), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n774), .B(new_n945), .C1(new_n968), .C2(new_n970), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1011), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n977), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(G8), .A3(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1010), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n975), .A2(new_n984), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G286), .A2(G8), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n955), .B1(new_n946), .B2(KEYINPUT114), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1966), .B1(new_n1024), .B2(new_n950), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n971), .A2(G2084), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT120), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1966), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n954), .B(new_n952), .C1(new_n948), .C2(new_n949), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n944), .A2(new_n949), .A3(new_n945), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1026), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1023), .B1(new_n1027), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1027), .A2(new_n1034), .ZN(new_n1036));
  OAI211_X1 g611(.A(KEYINPUT51), .B(G8), .C1(new_n1036), .C2(G286), .ZN(new_n1037));
  OAI21_X1  g612(.A(G8), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1023), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1035), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1022), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1035), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n947), .A2(new_n950), .A3(new_n956), .ZN(new_n1045));
  AOI211_X1 g620(.A(KEYINPUT120), .B(new_n1026), .C1(new_n1045), .C2(new_n1028), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1032), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1039), .B1(new_n1048), .B2(new_n1023), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1040), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1044), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT62), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n940), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1018), .A2(new_n1054), .A3(G8), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1054), .B1(new_n1018), .B2(G8), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n977), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(G8), .B(G168), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1057), .A2(new_n1021), .A3(KEYINPUT63), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1010), .A2(new_n1020), .A3(new_n984), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(new_n1058), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1062), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1060), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n749), .A2(new_n986), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n997), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1020), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1070), .A2(new_n1003), .B1(new_n1071), .B2(new_n1010), .ZN(new_n1072));
  XOR2_X1   g647(.A(G299), .B(KEYINPUT57), .Z(new_n1073));
  OR2_X1    g648(.A1(new_n981), .A2(G1956), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT56), .B(G2072), .Z(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n962), .A2(new_n964), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1073), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1077), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n981), .A2(G1956), .ZN(new_n1080));
  XNOR2_X1  g655(.A(G299), .B(KEYINPUT57), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT61), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1074), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT61), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n985), .A2(G2067), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1013), .B2(G1348), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1090), .A2(KEYINPUT60), .A3(new_n599), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1090), .B(new_n600), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(KEYINPUT60), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT59), .ZN(new_n1095));
  INV_X1    g670(.A(new_n985), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT58), .B(G1341), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n965), .A2(G1996), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1094), .A2(KEYINPUT59), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1098), .A2(new_n549), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1098), .B2(new_n549), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1095), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1088), .A2(new_n1093), .A3(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1090), .A2(new_n600), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1078), .B1(new_n1104), .B2(new_n1085), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n973), .B(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G171), .B(KEYINPUT54), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n920), .A2(new_n941), .A3(G2078), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n918), .A2(new_n962), .A3(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1108), .A2(new_n966), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(new_n984), .A3(new_n1020), .A4(new_n1010), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1109), .B1(new_n960), .B2(new_n974), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1106), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1067), .B(new_n1072), .C1(new_n1041), .C2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1053), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1043), .A2(new_n1052), .A3(new_n940), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n939), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n935), .A2(new_n933), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT48), .Z(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n930), .A2(KEYINPUT46), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n930), .A2(KEYINPUT46), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n921), .B1(new_n922), .B2(new_n853), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT47), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n925), .A2(new_n927), .A3(new_n931), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n791), .A2(G2067), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n921), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1125), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT126), .B1(new_n1120), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1117), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1022), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1051), .B2(KEYINPUT62), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1139));
  OAI21_X1  g714(.A(KEYINPUT124), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1140), .A3(new_n1119), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n938), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1134), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1135), .A2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g721(.A(G319), .ZN(new_n1148));
  NOR4_X1   g722(.A1(G229), .A2(G401), .A3(new_n1148), .A4(G227), .ZN(new_n1149));
  NAND4_X1  g723(.A1(new_n913), .A2(new_n866), .A3(new_n914), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n1151));
  XNOR2_X1  g725(.A(new_n1150), .B(new_n1151), .ZN(G308));
  XNOR2_X1  g726(.A(new_n1150), .B(KEYINPUT127), .ZN(G225));
endmodule


