

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U323 ( .A(n411), .B(KEYINPUT102), .ZN(n412) );
  XNOR2_X1 U324 ( .A(KEYINPUT41), .B(n573), .ZN(n555) );
  XNOR2_X1 U325 ( .A(n507), .B(KEYINPUT47), .ZN(n508) );
  XNOR2_X1 U326 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U327 ( .A(KEYINPUT91), .ZN(n387) );
  XNOR2_X1 U328 ( .A(n543), .B(KEYINPUT123), .ZN(n544) );
  NOR2_X1 U329 ( .A1(n408), .A2(n407), .ZN(n453) );
  XNOR2_X1 U330 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U331 ( .A(n545), .B(n544), .ZN(n546) );
  NOR2_X1 U332 ( .A1(n528), .A2(n491), .ZN(n513) );
  XNOR2_X1 U333 ( .A(n390), .B(n389), .ZN(n393) );
  XNOR2_X1 U334 ( .A(n446), .B(n445), .ZN(n499) );
  XNOR2_X1 U335 ( .A(KEYINPUT124), .B(n552), .ZN(n561) );
  XNOR2_X1 U336 ( .A(n413), .B(n412), .ZN(n484) );
  XNOR2_X1 U337 ( .A(n395), .B(n394), .ZN(n540) );
  XNOR2_X1 U338 ( .A(n449), .B(G43GAT), .ZN(n450) );
  XNOR2_X1 U339 ( .A(n451), .B(n450), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n291) );
  XNOR2_X1 U341 ( .A(G218GAT), .B(G92GAT), .ZN(n290) );
  XNOR2_X1 U342 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U343 ( .A(n292), .B(KEYINPUT11), .Z(n294) );
  XOR2_X1 U344 ( .A(G190GAT), .B(KEYINPUT78), .Z(n386) );
  XNOR2_X1 U345 ( .A(G36GAT), .B(n386), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n299) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n295), .B(KEYINPUT74), .ZN(n441) );
  XOR2_X1 U349 ( .A(KEYINPUT9), .B(n441), .Z(n297) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U352 ( .A(n299), .B(n298), .Z(n308) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n300), .B(G29GAT), .ZN(n301) );
  XOR2_X1 U355 ( .A(n301), .B(KEYINPUT70), .Z(n303) );
  XNOR2_X1 U356 ( .A(G50GAT), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n420) );
  XOR2_X1 U358 ( .A(KEYINPUT65), .B(G162GAT), .Z(n305) );
  XNOR2_X1 U359 ( .A(G134GAT), .B(G106GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n420), .B(n306), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n506) );
  XNOR2_X1 U363 ( .A(KEYINPUT36), .B(n506), .ZN(n579) );
  XNOR2_X1 U364 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n309), .B(KEYINPUT72), .ZN(n430) );
  XOR2_X1 U366 ( .A(n430), .B(KEYINPUT15), .Z(n311) );
  NAND2_X1 U367 ( .A1(G231GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U368 ( .A(n311), .B(n310), .ZN(n326) );
  XOR2_X1 U369 ( .A(KEYINPUT14), .B(G64GAT), .Z(n313) );
  XNOR2_X1 U370 ( .A(G8GAT), .B(G127GAT), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U372 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n315) );
  XNOR2_X1 U373 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n324) );
  XOR2_X1 U376 ( .A(G78GAT), .B(G211GAT), .Z(n319) );
  XNOR2_X1 U377 ( .A(G183GAT), .B(G71GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U379 ( .A(n320), .B(G155GAT), .Z(n322) );
  XOR2_X1 U380 ( .A(G15GAT), .B(G1GAT), .Z(n423) );
  XNOR2_X1 U381 ( .A(G22GAT), .B(n423), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n326), .B(n325), .ZN(n576) );
  INV_X1 U385 ( .A(n576), .ZN(n560) );
  XOR2_X1 U386 ( .A(G85GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U387 ( .A(G29GAT), .B(G141GAT), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U389 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n330) );
  XNOR2_X1 U390 ( .A(G120GAT), .B(G57GAT), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U392 ( .A(n332), .B(n331), .Z(n337) );
  XOR2_X1 U393 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n334) );
  NAND2_X1 U394 ( .A1(G225GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U396 ( .A(KEYINPUT88), .B(n335), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U398 ( .A(KEYINPUT6), .B(KEYINPUT87), .Z(n339) );
  XNOR2_X1 U399 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U401 ( .A(n341), .B(n340), .Z(n347) );
  XOR2_X1 U402 ( .A(G127GAT), .B(KEYINPUT0), .Z(n343) );
  XNOR2_X1 U403 ( .A(G113GAT), .B(G134GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n371) );
  XOR2_X1 U405 ( .A(G155GAT), .B(KEYINPUT3), .Z(n345) );
  XNOR2_X1 U406 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n371), .B(n348), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n547) );
  XOR2_X1 U410 ( .A(n348), .B(KEYINPUT24), .Z(n350) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .Z(n426) );
  XNOR2_X1 U412 ( .A(G50GAT), .B(n426), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n356) );
  XOR2_X1 U414 ( .A(G78GAT), .B(G148GAT), .Z(n352) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n442) );
  XOR2_X1 U417 ( .A(n442), .B(KEYINPUT84), .Z(n354) );
  NAND2_X1 U418 ( .A1(G228GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U420 ( .A(n356), .B(n355), .Z(n364) );
  XOR2_X1 U421 ( .A(KEYINPUT21), .B(G218GAT), .Z(n358) );
  XNOR2_X1 U422 ( .A(KEYINPUT85), .B(G211GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U424 ( .A(G197GAT), .B(n359), .Z(n384) );
  XOR2_X1 U425 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n361) );
  XNOR2_X1 U426 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n384), .B(n362), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n364), .B(n363), .ZN(n548) );
  XOR2_X1 U430 ( .A(G99GAT), .B(G190GAT), .Z(n366) );
  XNOR2_X1 U431 ( .A(G169GAT), .B(G43GAT), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U433 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n368) );
  XNOR2_X1 U434 ( .A(G15GAT), .B(KEYINPUT82), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n380) );
  XOR2_X1 U437 ( .A(G120GAT), .B(G71GAT), .Z(n429) );
  XOR2_X1 U438 ( .A(n429), .B(n371), .Z(n373) );
  NAND2_X1 U439 ( .A1(G227GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U441 ( .A(n374), .B(G176GAT), .Z(n378) );
  XOR2_X1 U442 ( .A(G183GAT), .B(KEYINPUT17), .Z(n376) );
  XNOR2_X1 U443 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n391), .B(KEYINPUT64), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n380), .B(n379), .ZN(n515) );
  INV_X1 U448 ( .A(n515), .ZN(n550) );
  XOR2_X1 U449 ( .A(G92GAT), .B(G64GAT), .Z(n382) );
  XNOR2_X1 U450 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U452 ( .A(G176GAT), .B(n383), .ZN(n443) );
  XNOR2_X1 U453 ( .A(n384), .B(n443), .ZN(n395) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(G36GAT), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n385), .B(G8GAT), .ZN(n425) );
  XOR2_X1 U456 ( .A(n386), .B(n425), .Z(n390) );
  NAND2_X1 U457 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U458 ( .A(n391), .B(KEYINPUT92), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n394) );
  NAND2_X1 U460 ( .A1(n550), .A2(n540), .ZN(n396) );
  NAND2_X1 U461 ( .A1(n548), .A2(n396), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n397), .B(KEYINPUT25), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n540), .B(KEYINPUT27), .ZN(n403) );
  NOR2_X1 U464 ( .A1(n548), .A2(n550), .ZN(n398) );
  XNOR2_X1 U465 ( .A(KEYINPUT26), .B(n398), .ZN(n567) );
  AND2_X1 U466 ( .A1(n403), .A2(n567), .ZN(n399) );
  NOR2_X1 U467 ( .A1(n400), .A2(n399), .ZN(n401) );
  XOR2_X1 U468 ( .A(KEYINPUT95), .B(n401), .Z(n402) );
  NOR2_X1 U469 ( .A1(n547), .A2(n402), .ZN(n408) );
  NAND2_X1 U470 ( .A1(n547), .A2(n403), .ZN(n528) );
  XOR2_X1 U471 ( .A(n548), .B(KEYINPUT28), .Z(n404) );
  XNOR2_X1 U472 ( .A(KEYINPUT66), .B(n404), .ZN(n491) );
  XOR2_X1 U473 ( .A(n513), .B(KEYINPUT93), .Z(n405) );
  NAND2_X1 U474 ( .A1(n515), .A2(n405), .ZN(n406) );
  XOR2_X1 U475 ( .A(KEYINPUT94), .B(n406), .Z(n407) );
  NOR2_X1 U476 ( .A1(n560), .A2(n453), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n409), .B(KEYINPUT101), .ZN(n410) );
  NOR2_X1 U478 ( .A1(n579), .A2(n410), .ZN(n413) );
  XOR2_X1 U479 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n411) );
  XOR2_X1 U480 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n415) );
  NAND2_X1 U481 ( .A1(G229GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U483 ( .A(n416), .B(KEYINPUT30), .Z(n422) );
  XOR2_X1 U484 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n418) );
  XNOR2_X1 U485 ( .A(G197GAT), .B(G113GAT), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U488 ( .A(n422), .B(n421), .Z(n424) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n529) );
  XOR2_X1 U492 ( .A(KEYINPUT71), .B(n529), .Z(n553) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n434) );
  INV_X1 U494 ( .A(n434), .ZN(n432) );
  AND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  INV_X1 U496 ( .A(n433), .ZN(n431) );
  NAND2_X1 U497 ( .A1(n432), .A2(n431), .ZN(n436) );
  NAND2_X1 U498 ( .A1(n434), .A2(n433), .ZN(n435) );
  NAND2_X1 U499 ( .A1(n436), .A2(n435), .ZN(n440) );
  XOR2_X1 U500 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n438) );
  XNOR2_X1 U501 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n437) );
  XOR2_X1 U502 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n444) );
  INV_X1 U505 ( .A(n499), .ZN(n573) );
  NAND2_X1 U506 ( .A1(n553), .A2(n573), .ZN(n456) );
  NOR2_X1 U507 ( .A1(n484), .A2(n456), .ZN(n448) );
  XNOR2_X1 U508 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n472) );
  NAND2_X1 U510 ( .A1(n472), .A2(n550), .ZN(n451) );
  XOR2_X1 U511 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n449) );
  XNOR2_X1 U512 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n461) );
  XOR2_X1 U513 ( .A(G1GAT), .B(KEYINPUT98), .Z(n459) );
  INV_X1 U514 ( .A(n506), .ZN(n564) );
  NOR2_X1 U515 ( .A1(n564), .A2(n576), .ZN(n452) );
  XNOR2_X1 U516 ( .A(n452), .B(KEYINPUT16), .ZN(n455) );
  INV_X1 U517 ( .A(n453), .ZN(n454) );
  NAND2_X1 U518 ( .A1(n455), .A2(n454), .ZN(n474) );
  NOR2_X1 U519 ( .A1(n456), .A2(n474), .ZN(n457) );
  XNOR2_X1 U520 ( .A(KEYINPUT96), .B(n457), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n547), .A2(n466), .ZN(n458) );
  XNOR2_X1 U522 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U523 ( .A(n461), .B(n460), .ZN(G1324GAT) );
  NAND2_X1 U524 ( .A1(n466), .A2(n540), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n462), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U526 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n464) );
  NAND2_X1 U527 ( .A1(n466), .A2(n550), .ZN(n463) );
  XNOR2_X1 U528 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U529 ( .A(G15GAT), .B(n465), .Z(G1326GAT) );
  NAND2_X1 U530 ( .A1(n466), .A2(n491), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n467), .B(KEYINPUT100), .ZN(n468) );
  XNOR2_X1 U532 ( .A(G22GAT), .B(n468), .ZN(G1327GAT) );
  NAND2_X1 U533 ( .A1(n547), .A2(n472), .ZN(n470) );
  XOR2_X1 U534 ( .A(G29GAT), .B(KEYINPUT39), .Z(n469) );
  XNOR2_X1 U535 ( .A(n470), .B(n469), .ZN(G1328GAT) );
  NAND2_X1 U536 ( .A1(n540), .A2(n472), .ZN(n471) );
  XNOR2_X1 U537 ( .A(n471), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U538 ( .A1(n491), .A2(n472), .ZN(n473) );
  XNOR2_X1 U539 ( .A(n473), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U540 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n476) );
  INV_X1 U541 ( .A(n529), .ZN(n569) );
  NAND2_X1 U542 ( .A1(n555), .A2(n569), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n483), .A2(n474), .ZN(n479) );
  NAND2_X1 U544 ( .A1(n547), .A2(n479), .ZN(n475) );
  XNOR2_X1 U545 ( .A(n476), .B(n475), .ZN(G1332GAT) );
  NAND2_X1 U546 ( .A1(n540), .A2(n479), .ZN(n477) );
  XNOR2_X1 U547 ( .A(n477), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U548 ( .A1(n550), .A2(n479), .ZN(n478) );
  XNOR2_X1 U549 ( .A(n478), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n481) );
  NAND2_X1 U551 ( .A1(n479), .A2(n491), .ZN(n480) );
  XNOR2_X1 U552 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U553 ( .A(G78GAT), .B(n482), .ZN(G1335GAT) );
  NOR2_X1 U554 ( .A1(n484), .A2(n483), .ZN(n492) );
  NAND2_X1 U555 ( .A1(n547), .A2(n492), .ZN(n485) );
  XNOR2_X1 U556 ( .A(G85GAT), .B(n485), .ZN(G1336GAT) );
  XOR2_X1 U557 ( .A(G92GAT), .B(KEYINPUT107), .Z(n487) );
  NAND2_X1 U558 ( .A1(n492), .A2(n540), .ZN(n486) );
  XNOR2_X1 U559 ( .A(n487), .B(n486), .ZN(G1337GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n489) );
  NAND2_X1 U561 ( .A1(n492), .A2(n550), .ZN(n488) );
  XNOR2_X1 U562 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U563 ( .A(G99GAT), .B(n490), .ZN(G1338GAT) );
  XNOR2_X1 U564 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n496) );
  XOR2_X1 U565 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n494) );
  NAND2_X1 U566 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U567 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U568 ( .A(n496), .B(n495), .ZN(G1339GAT) );
  INV_X1 U569 ( .A(n553), .ZN(n501) );
  NOR2_X1 U570 ( .A1(n579), .A2(n576), .ZN(n497) );
  XOR2_X1 U571 ( .A(KEYINPUT45), .B(n497), .Z(n498) );
  NOR2_X1 U572 ( .A1(n499), .A2(n498), .ZN(n500) );
  NAND2_X1 U573 ( .A1(n501), .A2(n500), .ZN(n511) );
  XNOR2_X1 U574 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n503) );
  AND2_X1 U575 ( .A1(n555), .A2(n529), .ZN(n502) );
  XNOR2_X1 U576 ( .A(n503), .B(n502), .ZN(n504) );
  NOR2_X1 U577 ( .A1(n560), .A2(n504), .ZN(n505) );
  NAND2_X1 U578 ( .A1(n506), .A2(n505), .ZN(n509) );
  XNOR2_X1 U579 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n507) );
  NAND2_X1 U580 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n512), .B(KEYINPUT48), .ZN(n541) );
  NAND2_X1 U582 ( .A1(n541), .A2(n513), .ZN(n514) );
  NOR2_X1 U583 ( .A1(n515), .A2(n514), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n524), .A2(n553), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n516), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n518) );
  NAND2_X1 U587 ( .A1(n524), .A2(n555), .ZN(n517) );
  XNOR2_X1 U588 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U589 ( .A(G120GAT), .B(n519), .Z(G1341GAT) );
  XNOR2_X1 U590 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n523) );
  XOR2_X1 U591 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n521) );
  NAND2_X1 U592 ( .A1(n524), .A2(n560), .ZN(n520) );
  XNOR2_X1 U593 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U594 ( .A(n523), .B(n522), .ZN(G1342GAT) );
  XOR2_X1 U595 ( .A(G134GAT), .B(KEYINPUT51), .Z(n526) );
  NAND2_X1 U596 ( .A1(n524), .A2(n564), .ZN(n525) );
  XNOR2_X1 U597 ( .A(n526), .B(n525), .ZN(G1343GAT) );
  NAND2_X1 U598 ( .A1(n541), .A2(n567), .ZN(n527) );
  NOR2_X1 U599 ( .A1(n528), .A2(n527), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n538), .A2(n529), .ZN(n530) );
  XNOR2_X1 U601 ( .A(n530), .B(KEYINPUT118), .ZN(n531) );
  XNOR2_X1 U602 ( .A(G141GAT), .B(n531), .ZN(G1344GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n533) );
  NAND2_X1 U604 ( .A1(n538), .A2(n555), .ZN(n532) );
  XNOR2_X1 U605 ( .A(n533), .B(n532), .ZN(n535) );
  XOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT52), .Z(n534) );
  XNOR2_X1 U607 ( .A(n535), .B(n534), .ZN(G1345GAT) );
  NAND2_X1 U608 ( .A1(n538), .A2(n560), .ZN(n536) );
  XNOR2_X1 U609 ( .A(n536), .B(KEYINPUT120), .ZN(n537) );
  XNOR2_X1 U610 ( .A(G155GAT), .B(n537), .ZN(G1346GAT) );
  NAND2_X1 U611 ( .A1(n564), .A2(n538), .ZN(n539) );
  XNOR2_X1 U612 ( .A(n539), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT121), .B(n540), .Z(n542) );
  NAND2_X1 U614 ( .A1(n542), .A2(n541), .ZN(n545) );
  XOR2_X1 U615 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n543) );
  NOR2_X1 U616 ( .A1(n547), .A2(n546), .ZN(n568) );
  NAND2_X1 U617 ( .A1(n548), .A2(n568), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n549), .B(KEYINPUT55), .ZN(n551) );
  AND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n561), .A2(n553), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n557) );
  NAND2_X1 U623 ( .A1(n555), .A2(n561), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT125), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT126), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(n563), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n564), .A2(n561), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n578) );
  NOR2_X1 U634 ( .A1(n569), .A2(n578), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n578), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n578), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

