

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579;

  NOR2_X1 U321 ( .A1(n533), .A2(n422), .ZN(n563) );
  XNOR2_X2 U322 ( .A(n442), .B(KEYINPUT117), .ZN(n556) );
  XNOR2_X1 U323 ( .A(KEYINPUT47), .B(KEYINPUT108), .ZN(n398) );
  XNOR2_X1 U324 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U325 ( .A(KEYINPUT45), .B(KEYINPUT109), .ZN(n400) );
  XNOR2_X1 U326 ( .A(n401), .B(n400), .ZN(n403) );
  XNOR2_X1 U327 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U328 ( .A(n399), .B(n398), .ZN(n405) );
  INV_X1 U329 ( .A(KEYINPUT77), .ZN(n374) );
  XNOR2_X1 U330 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U331 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U332 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U333 ( .A(n337), .B(n336), .ZN(n567) );
  XNOR2_X1 U334 ( .A(n445), .B(G183GAT), .ZN(n446) );
  XNOR2_X1 U335 ( .A(n447), .B(n446), .ZN(G1350GAT) );
  XOR2_X1 U336 ( .A(G141GAT), .B(G22GAT), .Z(n338) );
  XOR2_X1 U337 ( .A(G211GAT), .B(KEYINPUT21), .Z(n290) );
  XNOR2_X1 U338 ( .A(G197GAT), .B(G218GAT), .ZN(n289) );
  XNOR2_X1 U339 ( .A(n290), .B(n289), .ZN(n417) );
  XOR2_X1 U340 ( .A(n417), .B(G204GAT), .Z(n292) );
  NAND2_X1 U341 ( .A1(G228GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U343 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n294) );
  XNOR2_X1 U344 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U346 ( .A(n296), .B(n295), .Z(n300) );
  XNOR2_X1 U347 ( .A(G106GAT), .B(G78GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n297), .B(G148GAT), .ZN(n331) );
  XNOR2_X1 U349 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n298), .B(KEYINPUT2), .ZN(n313) );
  XNOR2_X1 U351 ( .A(n331), .B(n313), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n338), .B(n301), .ZN(n302) );
  XNOR2_X1 U354 ( .A(G50GAT), .B(G162GAT), .ZN(n381) );
  XNOR2_X1 U355 ( .A(n302), .B(n381), .ZN(n457) );
  XOR2_X1 U356 ( .A(G57GAT), .B(G148GAT), .Z(n304) );
  XNOR2_X1 U357 ( .A(G141GAT), .B(G1GAT), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n321) );
  XOR2_X1 U359 ( .A(G162GAT), .B(G127GAT), .Z(n306) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(G120GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U362 ( .A(G134GAT), .B(G85GAT), .Z(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n317) );
  XNOR2_X1 U364 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n309), .B(KEYINPUT1), .ZN(n310) );
  XOR2_X1 U366 ( .A(n310), .B(KEYINPUT5), .Z(n315) );
  XOR2_X1 U367 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n312) );
  XNOR2_X1 U368 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n435) );
  XNOR2_X1 U370 ( .A(n435), .B(n313), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n319) );
  NAND2_X1 U373 ( .A1(G225GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n533) );
  XOR2_X1 U376 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n358) );
  XNOR2_X1 U377 ( .A(G204GAT), .B(G92GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n322), .B(G64GAT), .ZN(n408) );
  XNOR2_X1 U379 ( .A(n408), .B(KEYINPUT72), .ZN(n324) );
  XOR2_X1 U380 ( .A(G85GAT), .B(KEYINPUT73), .Z(n380) );
  XNOR2_X1 U381 ( .A(G176GAT), .B(n380), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n329) );
  XNOR2_X1 U383 ( .A(G99GAT), .B(G71GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n325), .B(G120GAT), .ZN(n437) );
  XOR2_X1 U385 ( .A(n437), .B(KEYINPUT74), .Z(n327) );
  NAND2_X1 U386 ( .A1(G230GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n337) );
  XNOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n330), .B(KEYINPUT71), .ZN(n373) );
  XNOR2_X1 U391 ( .A(n331), .B(n373), .ZN(n335) );
  XOR2_X1 U392 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n333) );
  XNOR2_X1 U393 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n332) );
  XOR2_X1 U394 ( .A(n333), .B(n332), .Z(n334) );
  XOR2_X1 U395 ( .A(n567), .B(KEYINPUT41), .Z(n537) );
  XOR2_X1 U396 ( .A(G50GAT), .B(G43GAT), .Z(n340) );
  XOR2_X1 U397 ( .A(KEYINPUT69), .B(G1GAT), .Z(n368) );
  XNOR2_X1 U398 ( .A(n338), .B(n368), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U400 ( .A(n341), .B(G36GAT), .Z(n348) );
  XOR2_X1 U401 ( .A(G29GAT), .B(KEYINPUT7), .Z(n343) );
  XNOR2_X1 U402 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n393) );
  XOR2_X1 U404 ( .A(n393), .B(KEYINPUT67), .Z(n345) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(n346), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n356) );
  XOR2_X1 U409 ( .A(G8GAT), .B(G197GAT), .Z(n350) );
  XNOR2_X1 U410 ( .A(G113GAT), .B(G15GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U412 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n352) );
  XNOR2_X1 U413 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U415 ( .A(n354), .B(n353), .Z(n355) );
  XOR2_X1 U416 ( .A(n356), .B(n355), .Z(n564) );
  OR2_X1 U417 ( .A1(n537), .A2(n564), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n397) );
  XOR2_X1 U419 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n360) );
  XNOR2_X1 U420 ( .A(G64GAT), .B(KEYINPUT78), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n379) );
  XOR2_X1 U422 ( .A(G211GAT), .B(G78GAT), .Z(n362) );
  XNOR2_X1 U423 ( .A(G183GAT), .B(G71GAT), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U425 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n364) );
  XNOR2_X1 U426 ( .A(G22GAT), .B(G155GAT), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U428 ( .A(n366), .B(n365), .Z(n372) );
  XOR2_X1 U429 ( .A(G15GAT), .B(G127GAT), .Z(n427) );
  XOR2_X1 U430 ( .A(KEYINPUT76), .B(G8GAT), .Z(n411) );
  XOR2_X1 U431 ( .A(n427), .B(n411), .Z(n370) );
  NAND2_X1 U432 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n373), .B(KEYINPUT15), .ZN(n375) );
  XOR2_X1 U435 ( .A(n379), .B(n378), .Z(n572) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n383) );
  NAND2_X1 U437 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U439 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n385) );
  XNOR2_X1 U440 ( .A(KEYINPUT10), .B(G92GAT), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U442 ( .A(n387), .B(n386), .Z(n391) );
  XOR2_X1 U443 ( .A(G43GAT), .B(G134GAT), .Z(n428) );
  XNOR2_X1 U444 ( .A(G218GAT), .B(KEYINPUT64), .ZN(n388) );
  XOR2_X1 U445 ( .A(G36GAT), .B(G190GAT), .Z(n407) );
  XNOR2_X1 U446 ( .A(n388), .B(n407), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n428), .B(n389), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n392), .B(G106GAT), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n393), .B(G99GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n546) );
  AND2_X1 U452 ( .A1(n572), .A2(n546), .ZN(n396) );
  NAND2_X1 U453 ( .A1(n397), .A2(n396), .ZN(n399) );
  INV_X1 U454 ( .A(n572), .ZN(n526) );
  XOR2_X1 U455 ( .A(KEYINPUT36), .B(n546), .Z(n575) );
  NAND2_X1 U456 ( .A1(n526), .A2(n575), .ZN(n401) );
  INV_X1 U457 ( .A(n564), .ZN(n522) );
  AND2_X1 U458 ( .A1(n567), .A2(n564), .ZN(n402) );
  AND2_X1 U459 ( .A1(n403), .A2(n402), .ZN(n404) );
  NOR2_X1 U460 ( .A1(n405), .A2(n404), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n406), .B(KEYINPUT48), .ZN(n518) );
  XOR2_X1 U462 ( .A(n408), .B(n407), .Z(n410) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n412) );
  XOR2_X1 U465 ( .A(n412), .B(n411), .Z(n419) );
  XNOR2_X1 U466 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n413), .B(KEYINPUT17), .ZN(n414) );
  XOR2_X1 U468 ( .A(n414), .B(KEYINPUT18), .Z(n416) );
  XNOR2_X1 U469 ( .A(G169GAT), .B(G176GAT), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n438) );
  XNOR2_X1 U471 ( .A(n438), .B(n417), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n508) );
  XNOR2_X1 U473 ( .A(n508), .B(KEYINPUT115), .ZN(n420) );
  NOR2_X1 U474 ( .A1(n518), .A2(n420), .ZN(n421) );
  XOR2_X1 U475 ( .A(KEYINPUT54), .B(n421), .Z(n422) );
  NAND2_X1 U476 ( .A1(n457), .A2(n563), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n423), .B(KEYINPUT55), .ZN(n424) );
  XNOR2_X1 U478 ( .A(KEYINPUT116), .B(n424), .ZN(n441) );
  XOR2_X1 U479 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n426) );
  XNOR2_X1 U480 ( .A(KEYINPUT20), .B(KEYINPUT84), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U482 ( .A(KEYINPUT83), .B(G190GAT), .Z(n430) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U486 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U488 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n456) );
  BUF_X1 U491 ( .A(n456), .Z(n520) );
  NAND2_X1 U492 ( .A1(n441), .A2(n520), .ZN(n442) );
  NAND2_X1 U493 ( .A1(n556), .A2(n522), .ZN(n444) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(G1348GAT) );
  NAND2_X1 U496 ( .A1(n556), .A2(n526), .ZN(n447) );
  XOR2_X1 U497 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n445) );
  NAND2_X1 U498 ( .A1(n567), .A2(n522), .ZN(n479) );
  INV_X1 U499 ( .A(n546), .ZN(n555) );
  NOR2_X1 U500 ( .A1(n555), .A2(n572), .ZN(n448) );
  XNOR2_X1 U501 ( .A(KEYINPUT16), .B(n448), .ZN(n466) );
  XNOR2_X1 U502 ( .A(n520), .B(KEYINPUT87), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n508), .B(KEYINPUT27), .ZN(n459) );
  NAND2_X1 U504 ( .A1(n533), .A2(n459), .ZN(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n449), .B(n457), .ZN(n512) );
  NOR2_X1 U507 ( .A1(n450), .A2(n512), .ZN(n519) );
  NAND2_X1 U508 ( .A1(n451), .A2(n519), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n452), .B(KEYINPUT89), .ZN(n464) );
  NAND2_X1 U510 ( .A1(n456), .A2(n508), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n453), .B(KEYINPUT90), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n454), .A2(n457), .ZN(n455) );
  XOR2_X1 U513 ( .A(KEYINPUT25), .B(n455), .Z(n460) );
  NOR2_X1 U514 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(KEYINPUT26), .ZN(n562) );
  NAND2_X1 U516 ( .A1(n562), .A2(n459), .ZN(n532) );
  NAND2_X1 U517 ( .A1(n460), .A2(n532), .ZN(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT91), .B(n461), .ZN(n462) );
  NOR2_X1 U519 ( .A1(n533), .A2(n462), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT92), .B(n465), .Z(n476) );
  NAND2_X1 U522 ( .A1(n466), .A2(n476), .ZN(n492) );
  NOR2_X1 U523 ( .A1(n479), .A2(n492), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT93), .B(n467), .Z(n474) );
  NAND2_X1 U525 ( .A1(n533), .A2(n474), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(KEYINPUT34), .ZN(n469) );
  XNOR2_X1 U527 ( .A(G1GAT), .B(n469), .ZN(G1324GAT) );
  NAND2_X1 U528 ( .A1(n474), .A2(n508), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n472) );
  NAND2_X1 U531 ( .A1(n474), .A2(n520), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U533 ( .A(G15GAT), .B(n473), .ZN(G1326GAT) );
  NAND2_X1 U534 ( .A1(n512), .A2(n474), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n475), .B(G22GAT), .ZN(G1327GAT) );
  AND2_X1 U536 ( .A1(n572), .A2(n476), .ZN(n477) );
  NAND2_X1 U537 ( .A1(n575), .A2(n477), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT37), .B(n478), .Z(n503) );
  NOR2_X1 U539 ( .A1(n479), .A2(n503), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT38), .ZN(n490) );
  NAND2_X1 U541 ( .A1(n490), .A2(n533), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n482) );
  XNOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U546 ( .A(KEYINPUT95), .B(n485), .ZN(G1328GAT) );
  NAND2_X1 U547 ( .A1(n490), .A2(n508), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT98), .B(KEYINPUT40), .Z(n488) );
  NAND2_X1 U550 ( .A1(n490), .A2(n520), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U552 ( .A(G43GAT), .B(n489), .Z(G1330GAT) );
  NAND2_X1 U553 ( .A1(n490), .A2(n512), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n491), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT42), .B(KEYINPUT99), .Z(n494) );
  INV_X1 U556 ( .A(n537), .ZN(n552) );
  NAND2_X1 U557 ( .A1(n564), .A2(n552), .ZN(n504) );
  NOR2_X1 U558 ( .A1(n504), .A2(n492), .ZN(n498) );
  NAND2_X1 U559 ( .A1(n498), .A2(n533), .ZN(n493) );
  XNOR2_X1 U560 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n495), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n498), .A2(n508), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n496), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U564 ( .A1(n498), .A2(n520), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n497), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT100), .B(KEYINPUT43), .Z(n500) );
  NAND2_X1 U567 ( .A1(n498), .A2(n512), .ZN(n499) );
  XNOR2_X1 U568 ( .A(n500), .B(n499), .ZN(n502) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT101), .Z(n501) );
  XNOR2_X1 U570 ( .A(n502), .B(n501), .ZN(G1335GAT) );
  XOR2_X1 U571 ( .A(G85GAT), .B(KEYINPUT103), .Z(n507) );
  NOR2_X1 U572 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n505), .B(KEYINPUT102), .ZN(n513) );
  NAND2_X1 U574 ( .A1(n513), .A2(n533), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n508), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n509), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n520), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n510), .B(KEYINPUT104), .ZN(n511) );
  XNOR2_X1 U580 ( .A(G99GAT), .B(n511), .ZN(G1338GAT) );
  XNOR2_X1 U581 ( .A(G106GAT), .B(KEYINPUT105), .ZN(n517) );
  XOR2_X1 U582 ( .A(KEYINPUT106), .B(KEYINPUT44), .Z(n515) );
  NAND2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1339GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U587 ( .A1(n518), .A2(n521), .ZN(n529) );
  NAND2_X1 U588 ( .A1(n522), .A2(n529), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT49), .Z(n525) );
  NAND2_X1 U591 ( .A1(n529), .A2(n552), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  NAND2_X1 U593 ( .A1(n526), .A2(n529), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(KEYINPUT50), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(G134GAT), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U597 ( .A1(n529), .A2(n555), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1343GAT) );
  NOR2_X1 U599 ( .A1(n518), .A2(n532), .ZN(n534) );
  NAND2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n545) );
  NOR2_X1 U601 ( .A1(n564), .A2(n545), .ZN(n535) );
  XOR2_X1 U602 ( .A(KEYINPUT110), .B(n535), .Z(n536) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(n536), .ZN(G1344GAT) );
  NOR2_X1 U604 ( .A1(n545), .A2(n537), .ZN(n541) );
  XOR2_X1 U605 ( .A(KEYINPUT111), .B(KEYINPUT53), .Z(n539) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1345GAT) );
  NOR2_X1 U609 ( .A1(n572), .A2(n545), .ZN(n543) );
  XNOR2_X1 U610 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(n544), .ZN(G1346GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(G162GAT), .B(n547), .Z(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT114), .B(n548), .ZN(G1347GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n550) );
  XNOR2_X1 U617 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(KEYINPUT56), .B(n551), .Z(n554) );
  NAND2_X1 U620 ( .A1(n556), .A2(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1349GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n561) );
  XNOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n574) );
  NOR2_X1 U630 ( .A1(n564), .A2(n574), .ZN(n565) );
  XOR2_X1 U631 ( .A(n566), .B(n565), .Z(G1352GAT) );
  NOR2_X1 U632 ( .A1(n574), .A2(n567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n569) );
  XNOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n574), .ZN(n573) );
  XOR2_X1 U638 ( .A(G211GAT), .B(n573), .Z(G1354GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n578) );
  INV_X1 U640 ( .A(n574), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

