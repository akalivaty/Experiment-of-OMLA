//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT76), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G211gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT22), .B1(new_n211), .B2(G218gat), .ZN(new_n212));
  XOR2_X1   g011(.A(G197gat), .B(G204gat), .Z(new_n213));
  OAI21_X1  g012(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT22), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT76), .B(G211gat), .ZN(new_n216));
  INV_X1    g015(.A(G218gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n213), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT77), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G211gat), .B(G218gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n214), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n221), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT77), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(G141gat), .ZN(new_n228));
  INV_X1    g027(.A(G141gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT81), .A3(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(G141gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233));
  OR2_X1    g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(KEYINPUT2), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(G155gat), .A2(G162gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G141gat), .B(G148gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT2), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n225), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n222), .A2(new_n244), .A3(new_n224), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n242), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n236), .A2(new_n241), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n236), .A2(new_n241), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n253), .B1(new_n247), .B2(new_n242), .ZN(new_n254));
  OAI211_X1 g053(.A(G228gat), .B(G233gat), .C1(new_n254), .C2(KEYINPUT87), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n225), .A2(new_n245), .ZN(new_n256));
  OAI21_X1  g055(.A(G22gat), .B1(new_n256), .B2(new_n254), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n255), .B1(new_n252), .B2(new_n257), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n205), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n252), .A2(new_n257), .ZN(new_n261));
  INV_X1    g060(.A(new_n255), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n252), .A2(new_n255), .A3(new_n257), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n204), .A3(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G1gat), .B(G29gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT0), .ZN(new_n268));
  XNOR2_X1  g067(.A(G57gat), .B(G85gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G225gat), .A2(G233gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n273));
  INV_X1    g072(.A(G120gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G113gat), .ZN(new_n275));
  INV_X1    g074(.A(G113gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G120gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT1), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT71), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n279), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n276), .ZN(new_n288));
  NAND2_X1  g087(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(G120gat), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n275), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(KEYINPUT70), .A3(new_n275), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n280), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT4), .B1(new_n295), .B2(new_n253), .ZN(new_n296));
  AND2_X1   g095(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n297), .A2(new_n298), .A3(new_n274), .ZN(new_n299));
  INV_X1    g098(.A(new_n275), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n292), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n286), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n294), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n280), .ZN(new_n304));
  AND4_X1   g103(.A1(KEYINPUT4), .A2(new_n303), .A3(new_n253), .A4(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n273), .B1(new_n296), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n253), .A3(new_n304), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n295), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT85), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n290), .A2(KEYINPUT70), .A3(new_n275), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT70), .B1(new_n290), .B2(new_n275), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n314), .A2(new_n315), .A3(new_n286), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n316), .B2(new_n280), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n243), .A2(KEYINPUT82), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(new_n242), .B2(new_n253), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n303), .A2(KEYINPUT83), .A3(new_n304), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n249), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n317), .A2(new_n319), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n272), .B1(new_n312), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT39), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n271), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n317), .A2(new_n249), .A3(new_n320), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT84), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n317), .A2(new_n328), .A3(new_n249), .A4(new_n320), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n327), .A2(new_n272), .A3(new_n307), .A4(new_n329), .ZN(new_n330));
  AOI211_X1 g129(.A(new_n313), .B(new_n280), .C1(new_n293), .C2(new_n294), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT83), .B1(new_n303), .B2(new_n304), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n242), .B1(new_n236), .B2(new_n241), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(KEYINPUT82), .B2(new_n243), .ZN(new_n335));
  INV_X1    g134(.A(new_n321), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n306), .A2(new_n311), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n330), .B(KEYINPUT39), .C1(new_n338), .C2(new_n272), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n325), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT40), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n272), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT5), .B(new_n343), .C1(new_n333), .C2(new_n337), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n312), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n329), .A2(new_n307), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n272), .B1(new_n346), .B2(new_n327), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n296), .A2(new_n305), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n322), .A3(new_n272), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n345), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n271), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n354), .B(KEYINPUT78), .Z(new_n355));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT26), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(new_n356), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT68), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT27), .B(G183gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(G190gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G183gat), .ZN(new_n371));
  INV_X1    g170(.A(G183gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT27), .ZN(new_n373));
  AND4_X1   g172(.A1(new_n365), .A2(new_n368), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(KEYINPUT66), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT66), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G183gat), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT27), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT67), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n372), .B2(KEYINPUT27), .ZN(new_n381));
  INV_X1    g180(.A(G190gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n370), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n367), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n364), .B1(new_n375), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n358), .ZN(new_n388));
  NAND3_X1  g187(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n356), .A2(KEYINPUT23), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n390), .A2(new_n391), .A3(new_n360), .A4(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT25), .ZN(new_n395));
  AND4_X1   g194(.A1(KEYINPUT25), .A2(new_n391), .A3(new_n360), .A4(new_n393), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n358), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT24), .ZN(new_n399));
  NAND3_X1  g198(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n376), .A2(new_n378), .A3(new_n382), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n389), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n394), .A2(new_n395), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n355), .B1(new_n386), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n359), .A2(new_n363), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT66), .B(G183gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT27), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT28), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n368), .A2(new_n371), .A3(new_n373), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT68), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n366), .A2(new_n365), .A3(new_n368), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n406), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n388), .A2(new_n389), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n391), .A2(new_n360), .A3(new_n393), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n395), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n403), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n225), .B(new_n405), .C1(new_n421), .C2(new_n355), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n244), .B1(new_n386), .B2(new_n404), .ZN(new_n424));
  INV_X1    g223(.A(new_n355), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n225), .A4(new_n405), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n405), .B1(new_n421), .B2(new_n355), .ZN(new_n429));
  INV_X1    g228(.A(new_n225), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n423), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G8gat), .B(G36gat), .Z(new_n433));
  XOR2_X1   g232(.A(G64gat), .B(G92gat), .Z(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n353), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n353), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n423), .A2(new_n428), .A3(new_n431), .A4(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n435), .B(KEYINPUT80), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n325), .A2(KEYINPUT40), .A3(new_n339), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n342), .A2(new_n352), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n432), .A2(KEYINPUT37), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n423), .A2(new_n428), .A3(new_n431), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n436), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT38), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT88), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT88), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n451), .B(KEYINPUT38), .C1(new_n445), .C2(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n432), .A2(new_n436), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n422), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(KEYINPUT37), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n447), .B2(new_n458), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n351), .A2(new_n271), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n328), .B1(new_n333), .B2(new_n249), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n329), .A2(new_n307), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n343), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n343), .B1(new_n333), .B2(new_n337), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(new_n348), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n465), .A2(new_n468), .B1(new_n312), .B2(new_n344), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n460), .B1(new_n469), .B2(new_n270), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n468), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n471), .A2(new_n270), .A3(new_n345), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n459), .B(new_n462), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n266), .B(new_n444), .C1(new_n453), .C2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n295), .B1(new_n386), .B2(new_n404), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n303), .A2(new_n304), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n415), .A3(new_n420), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT34), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n479), .B(KEYINPUT64), .Z(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(KEYINPUT34), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G43gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT73), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT74), .ZN(new_n489));
  XNOR2_X1  g288(.A(G71gat), .B(G99gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT74), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n488), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n477), .A3(new_n482), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT72), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT32), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n498), .B2(KEYINPUT32), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT75), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT75), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n499), .B(new_n505), .C1(new_n501), .C2(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT32), .B(new_n498), .C1(new_n496), .C2(new_n497), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n486), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n508), .ZN(new_n510));
  AOI211_X1 g309(.A(new_n510), .B(new_n485), .C1(new_n504), .C2(new_n506), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT36), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n498), .A2(KEYINPUT32), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT72), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT32), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n505), .B1(new_n516), .B2(new_n499), .ZN(new_n517));
  INV_X1    g316(.A(new_n506), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n508), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n485), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT36), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n507), .A2(new_n508), .A3(new_n486), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n462), .B1(new_n470), .B2(new_n472), .ZN(new_n524));
  INV_X1    g323(.A(new_n442), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n260), .A2(new_n265), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n474), .A2(new_n512), .A3(new_n523), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n520), .A2(new_n522), .A3(new_n266), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT35), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n509), .A2(new_n511), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n469), .A2(new_n270), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n352), .A2(new_n533), .A3(new_n460), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n442), .B1(new_n534), .B2(new_n462), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT35), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n532), .A2(new_n535), .A3(new_n536), .A4(new_n266), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n529), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT13), .Z(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT16), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(G1gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(G1gat), .B2(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G8gat), .ZN(new_n546));
  INV_X1    g345(.A(G8gat), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n544), .B(new_n547), .C1(G1gat), .C2(new_n542), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G43gat), .B(G50gat), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  NOR2_X1   g350(.A1(G29gat), .A2(G36gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n555));
  NAND2_X1  g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT90), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n551), .A2(new_n554), .A3(new_n555), .A4(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n552), .B(KEYINPUT14), .ZN(new_n560));
  OAI211_X1 g359(.A(KEYINPUT15), .B(new_n550), .C1(new_n560), .C2(new_n557), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n561), .A3(KEYINPUT91), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n561), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n549), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n562), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n548), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT91), .B1(new_n559), .B2(new_n561), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n541), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n568), .B1(new_n567), .B2(new_n569), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(G229gat), .B2(G233gat), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT17), .B1(new_n565), .B2(new_n562), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n559), .A2(KEYINPUT17), .A3(new_n561), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n549), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n572), .B(new_n574), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT92), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n571), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n572), .B(new_n540), .C1(new_n575), .C2(new_n577), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n573), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT93), .ZN(new_n586));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT12), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n585), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n579), .A2(KEYINPUT92), .B1(new_n573), .B2(new_n583), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n592), .B1(new_n595), .B2(new_n582), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n593), .B1(new_n573), .B2(new_n583), .ZN(new_n597));
  INV_X1    g396(.A(new_n579), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT93), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n594), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n539), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n524), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G57gat), .B(G64gat), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(G71gat), .A2(G78gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n612), .B(new_n606), .C1(new_n607), .C2(new_n608), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G127gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n549), .B1(new_n617), .B2(new_n616), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT95), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n626));
  INV_X1    g425(.A(G155gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n625), .B(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n567), .A2(new_n569), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G99gat), .B(G106gat), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G85gat), .A2(G92gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT7), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  INV_X1    g438(.A(G85gat), .ZN(new_n640));
  INV_X1    g439(.A(G92gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(KEYINPUT8), .A2(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n636), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n636), .B1(new_n638), .B2(new_n642), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n634), .A2(new_n646), .B1(KEYINPUT41), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n646), .B(KEYINPUT96), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n649), .B(new_n576), .C1(new_n633), .C2(KEYINPUT17), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G190gat), .B(G218gat), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n647), .A2(KEYINPUT41), .ZN(new_n654));
  XNOR2_X1  g453(.A(G134gat), .B(G162gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n652), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n648), .A2(new_n650), .A3(new_n657), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n653), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n653), .B2(new_n658), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n614), .B(new_n615), .C1(new_n644), .C2(new_n645), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n614), .A2(new_n615), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n638), .A2(new_n642), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n635), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n643), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G230gat), .A2(G233gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT97), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(G176gat), .B(G204gat), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n667), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n646), .A2(KEYINPUT10), .A3(new_n664), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n669), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n675), .A2(KEYINPUT98), .A3(new_n678), .A4(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n683), .A2(new_n672), .A3(new_n678), .A4(new_n674), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n675), .A2(new_n683), .ZN(new_n689));
  INV_X1    g488(.A(new_n678), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n632), .A2(new_n662), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n604), .A2(new_n605), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g496(.A1(new_n603), .A2(new_n694), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n442), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT100), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n547), .B1(new_n698), .B2(new_n442), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT99), .Z(new_n706));
  NAND3_X1  g505(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(G1325gat));
  AND2_X1   g506(.A1(new_n512), .A2(new_n523), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n698), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G15gat), .ZN(new_n711));
  INV_X1    g510(.A(new_n532), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n694), .A2(G15gat), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n603), .B2(new_n713), .ZN(G1326gat));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n527), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  NOR3_X1   g516(.A1(new_n632), .A2(new_n662), .A3(new_n692), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n604), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n719), .A2(G29gat), .A3(new_n524), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT45), .Z(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n312), .A2(new_n322), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n324), .A3(new_n343), .ZN(new_n724));
  AND4_X1   g523(.A1(KEYINPUT40), .A2(new_n339), .A3(new_n724), .A4(new_n270), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT40), .B1(new_n325), .B2(new_n339), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n441), .A2(new_n439), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n728), .A2(new_n437), .B1(new_n271), .B2(new_n351), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n527), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n469), .A2(new_n270), .A3(new_n460), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n432), .A2(new_n436), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n457), .A2(KEYINPUT37), .ZN(new_n733));
  INV_X1    g532(.A(new_n456), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n447), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n450), .A3(new_n534), .A4(new_n452), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n730), .A2(new_n738), .B1(new_n526), .B2(new_n527), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n739), .A2(new_n708), .B1(new_n531), .B2(new_n537), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n722), .B1(new_n740), .B2(new_n662), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n539), .A2(KEYINPUT44), .A3(new_n661), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n632), .B(KEYINPUT101), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n743), .A2(new_n602), .A3(new_n693), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT102), .A4(new_n744), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n605), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G29gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n721), .A2(new_n750), .ZN(G1328gat));
  NOR3_X1   g550(.A1(new_n719), .A2(G36gat), .A3(new_n525), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n747), .A2(new_n442), .A3(new_n748), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G36gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1329gat));
  XOR2_X1   g556(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n758));
  NAND3_X1  g557(.A1(new_n747), .A2(new_n709), .A3(new_n748), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G43gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n712), .A2(G43gat), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n539), .A2(new_n602), .A3(new_n718), .A4(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n758), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(KEYINPUT47), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n741), .A2(new_n742), .A3(new_n709), .A4(new_n744), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(G43gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT105), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT106), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n766), .B(KEYINPUT105), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n771));
  INV_X1    g570(.A(new_n762), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n759), .B2(G43gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n770), .B(new_n771), .C1(new_n773), .C2(new_n758), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n769), .A2(new_n774), .ZN(G1330gat));
  NOR3_X1   g574(.A1(new_n719), .A2(G50gat), .A3(new_n266), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n747), .A2(new_n527), .A3(new_n748), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(G50gat), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(G50gat), .ZN(new_n782));
  INV_X1    g581(.A(new_n745), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n527), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n778), .A2(new_n779), .B1(new_n781), .B2(new_n784), .ZN(G1331gat));
  NAND3_X1  g584(.A1(new_n632), .A2(new_n662), .A3(new_n692), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n740), .A2(new_n602), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n605), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g588(.A(new_n525), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT108), .Z(new_n792));
  NOR2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1333gat));
  NAND3_X1  g593(.A1(new_n787), .A2(G71gat), .A3(new_n709), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n532), .B(KEYINPUT109), .ZN(new_n796));
  NOR4_X1   g595(.A1(new_n740), .A2(new_n602), .A3(new_n786), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n797), .B2(G71gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n798), .B(new_n799), .Z(G1334gat));
  NAND2_X1  g599(.A1(new_n787), .A2(new_n527), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  INV_X1    g601(.A(new_n632), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n601), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT111), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n539), .A3(new_n661), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT51), .Z(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n640), .A3(new_n605), .A4(new_n692), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n741), .A2(new_n742), .A3(new_n692), .A4(new_n805), .ZN(new_n809));
  OAI21_X1  g608(.A(G85gat), .B1(new_n809), .B2(new_n524), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT112), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n813), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1336gat));
  NAND4_X1  g614(.A1(new_n807), .A2(new_n641), .A3(new_n442), .A4(new_n692), .ZN(new_n816));
  OAI21_X1  g615(.A(G92gat), .B1(new_n809), .B2(new_n525), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1337gat));
  XOR2_X1   g621(.A(KEYINPUT113), .B(G99gat), .Z(new_n823));
  NOR3_X1   g622(.A1(new_n712), .A2(new_n693), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n809), .B2(new_n708), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1338gat));
  NOR3_X1   g626(.A1(new_n266), .A2(new_n693), .A3(G106gat), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT114), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n807), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G106gat), .B1(new_n809), .B2(new_n266), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g632(.A1(new_n680), .A2(new_n670), .A3(new_n681), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n670), .B1(new_n680), .B2(new_n681), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n678), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT115), .ZN(new_n842));
  INV_X1    g641(.A(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT55), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(new_n845), .A3(new_n840), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n842), .A2(new_n844), .A3(new_n688), .A4(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n585), .A2(new_n593), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT93), .A3(new_n599), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n843), .A2(KEYINPUT55), .B1(new_n684), .B2(new_n687), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n852), .A2(KEYINPUT116), .A3(new_n846), .A4(new_n842), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n849), .A2(new_n851), .A3(new_n594), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n575), .A2(new_n577), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n566), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n566), .A2(new_n570), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n856), .A2(new_n540), .B1(new_n857), .B2(new_n541), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n858), .A2(new_n591), .B1(new_n597), .B2(new_n598), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n692), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n661), .B1(new_n854), .B2(new_n860), .ZN(new_n861));
  AND4_X1   g660(.A1(new_n661), .A2(new_n849), .A3(new_n859), .A4(new_n853), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n743), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n694), .A2(new_n602), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n530), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n605), .A2(new_n525), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n602), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n288), .B2(new_n289), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n276), .B2(new_n869), .ZN(G1340gat));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n868), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n693), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(new_n274), .ZN(G1341gat));
  OAI21_X1  g673(.A(G127gat), .B1(new_n872), .B2(new_n743), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n803), .A2(G127gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n872), .B2(new_n876), .ZN(G1342gat));
  OAI21_X1  g676(.A(G134gat), .B1(new_n872), .B2(new_n662), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n661), .A2(new_n525), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT117), .Z(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(G134gat), .A3(new_n524), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT56), .B1(new_n866), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n866), .A2(KEYINPUT56), .A3(new_n881), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n882), .B2(new_n883), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n708), .A2(new_n527), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n605), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n886), .B2(new_n885), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n863), .A2(new_n865), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n442), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n602), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n229), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT55), .B1(new_n839), .B2(KEYINPUT118), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(KEYINPUT118), .B2(new_n839), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n852), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n894), .B(new_n860), .C1(new_n601), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n662), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n851), .A2(new_n594), .A3(new_n852), .A4(new_n896), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n894), .B1(new_n900), .B2(new_n860), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(new_n862), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n864), .B1(new_n903), .B2(new_n803), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT57), .B1(new_n904), .B2(new_n266), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n709), .A2(new_n867), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n266), .B1(new_n863), .B2(new_n865), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n602), .A2(G141gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n893), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n893), .B(KEYINPUT58), .C1(new_n910), .C2(new_n911), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1344gat));
  NAND3_X1  g715(.A1(new_n891), .A2(new_n227), .A3(new_n692), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n662), .B2(new_n847), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n859), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n662), .A2(new_n847), .A3(new_n919), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n899), .A2(new_n901), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n803), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n865), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n266), .B1(new_n925), .B2(KEYINPUT123), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n864), .B1(new_n923), .B2(new_n803), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT57), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n889), .A2(KEYINPUT57), .A3(new_n527), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n907), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n692), .B(new_n906), .C1(new_n930), .C2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n918), .B1(new_n936), .B2(G148gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n910), .A2(new_n693), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n918), .A2(G148gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n917), .B1(new_n937), .B2(new_n940), .ZN(G1345gat));
  OAI21_X1  g740(.A(G155gat), .B1(new_n910), .B2(new_n743), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n891), .A2(new_n627), .A3(new_n632), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1346gat));
  OAI21_X1  g743(.A(G162gat), .B1(new_n910), .B2(new_n662), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n880), .A2(G162gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n890), .B2(new_n946), .ZN(G1347gat));
  NAND3_X1  g746(.A1(new_n866), .A2(new_n442), .A3(new_n524), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n601), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n524), .A2(new_n442), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n796), .A2(new_n527), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n889), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n602), .A2(G169gat), .ZN(new_n953));
  OAI22_X1  g752(.A1(new_n949), .A2(G169gat), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT124), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n952), .B2(new_n693), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n693), .A2(G176gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n948), .B2(new_n957), .ZN(G1349gat));
  NOR2_X1   g757(.A1(new_n952), .A2(new_n743), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g759(.A(new_n408), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n961), .B1(new_n959), .B2(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n632), .A2(new_n366), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n960), .A2(new_n962), .B1(new_n948), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n952), .B2(new_n662), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT61), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n661), .A2(new_n382), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n948), .B2(new_n968), .ZN(G1351gat));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n930), .B2(new_n935), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n907), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT121), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n929), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n527), .B1(new_n927), .B2(new_n928), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n908), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n977), .A3(KEYINPUT126), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n709), .A2(new_n950), .ZN(new_n979));
  INV_X1    g778(.A(G197gat), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n601), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n971), .A2(new_n978), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n885), .A2(new_n950), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n889), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n984), .B2(new_n601), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n982), .A2(new_n985), .ZN(G1352gat));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n978), .A3(new_n692), .A4(new_n979), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(G204gat), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n984), .A2(G204gat), .A3(new_n693), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT62), .ZN(new_n991));
  XOR2_X1   g790(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n992));
  OAI21_X1  g791(.A(new_n991), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n988), .A2(new_n993), .ZN(G1353gat));
  OAI211_X1 g793(.A(new_n632), .B(new_n979), .C1(new_n930), .C2(new_n935), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n632), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n997), .B1(new_n974), .B2(new_n977), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT63), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n998), .A2(new_n999), .A3(new_n207), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n632), .A2(new_n216), .ZN(new_n1001));
  OAI22_X1  g800(.A1(new_n996), .A2(new_n1000), .B1(new_n984), .B2(new_n1001), .ZN(G1354gat));
  NOR2_X1   g801(.A1(new_n662), .A2(new_n217), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n971), .A2(new_n978), .A3(new_n979), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n217), .B1(new_n984), .B2(new_n662), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1355gat));
endmodule


