

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U325 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U326 ( .A(n448), .B(n447), .ZN(n503) );
  XOR2_X1 U327 ( .A(n364), .B(n363), .Z(n293) );
  XOR2_X1 U328 ( .A(n305), .B(n304), .Z(n294) );
  INV_X1 U329 ( .A(KEYINPUT6), .ZN(n368) );
  XNOR2_X1 U330 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U331 ( .A(n371), .B(n370), .ZN(n372) );
  INV_X1 U332 ( .A(KEYINPUT48), .ZN(n465) );
  XNOR2_X1 U333 ( .A(n365), .B(n293), .ZN(n374) );
  XNOR2_X1 U334 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n468) );
  XNOR2_X1 U335 ( .A(n466), .B(n465), .ZN(n534) );
  XNOR2_X1 U336 ( .A(n374), .B(n373), .ZN(n378) );
  XNOR2_X1 U337 ( .A(n469), .B(n468), .ZN(n571) );
  XNOR2_X1 U338 ( .A(n306), .B(n294), .ZN(n307) );
  XNOR2_X1 U339 ( .A(n381), .B(n404), .ZN(n382) );
  XNOR2_X1 U340 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U341 ( .A(n308), .B(n307), .ZN(n578) );
  XNOR2_X1 U342 ( .A(n383), .B(n382), .ZN(n440) );
  INV_X1 U343 ( .A(G43GAT), .ZN(n449) );
  XNOR2_X1 U344 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n478) );
  XNOR2_X1 U345 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U346 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n452), .B(n451), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT99), .B(KEYINPUT38), .Z(n448) );
  XNOR2_X1 U349 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n296) );
  AND2_X1 U350 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(n297), .B(KEYINPUT68), .Z(n303) );
  XOR2_X1 U353 ( .A(G64GAT), .B(G92GAT), .Z(n299) );
  XNOR2_X1 U354 ( .A(G176GAT), .B(G204GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n386) );
  XOR2_X1 U356 ( .A(KEYINPUT67), .B(KEYINPUT13), .Z(n301) );
  XNOR2_X1 U357 ( .A(G71GAT), .B(G78GAT), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n355) );
  XNOR2_X1 U359 ( .A(n386), .B(n355), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n308) );
  XOR2_X1 U361 ( .A(G120GAT), .B(G148GAT), .Z(n375) );
  XOR2_X1 U362 ( .A(G99GAT), .B(G85GAT), .Z(n328) );
  XNOR2_X1 U363 ( .A(n375), .B(n328), .ZN(n306) );
  XOR2_X1 U364 ( .A(KEYINPUT69), .B(KEYINPUT32), .Z(n305) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(G57GAT), .ZN(n304) );
  XOR2_X1 U366 ( .A(G1GAT), .B(G141GAT), .Z(n310) );
  XNOR2_X1 U367 ( .A(G169GAT), .B(G197GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U369 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n312) );
  XNOR2_X1 U370 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n325) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n315), .B(KEYINPUT7), .ZN(n327) );
  XOR2_X1 U375 ( .A(n327), .B(KEYINPUT65), .Z(n317) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n318), .B(G29GAT), .ZN(n323) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G36GAT), .Z(n321) );
  XNOR2_X1 U380 ( .A(G15GAT), .B(G22GAT), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n319), .B(KEYINPUT64), .ZN(n347) );
  XNOR2_X1 U382 ( .A(G113GAT), .B(n347), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n574) );
  INV_X1 U386 ( .A(n574), .ZN(n506) );
  NOR2_X1 U387 ( .A1(n578), .A2(n506), .ZN(n487) );
  XNOR2_X1 U388 ( .A(G36GAT), .B(G190GAT), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n326), .B(G218GAT), .ZN(n388) );
  XNOR2_X1 U390 ( .A(n327), .B(n388), .ZN(n341) );
  XOR2_X1 U391 ( .A(G29GAT), .B(G134GAT), .Z(n376) );
  XOR2_X1 U392 ( .A(n376), .B(n328), .Z(n330) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U395 ( .A(G92GAT), .B(KEYINPUT72), .Z(n332) );
  XNOR2_X1 U396 ( .A(G162GAT), .B(KEYINPUT70), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U398 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U399 ( .A(G50GAT), .B(G106GAT), .Z(n416) );
  XOR2_X1 U400 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n336) );
  XNOR2_X1 U401 ( .A(KEYINPUT10), .B(KEYINPUT71), .ZN(n335) );
  XNOR2_X1 U402 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n416), .B(n337), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n561) );
  XNOR2_X1 U406 ( .A(n561), .B(KEYINPUT36), .ZN(n584) );
  XOR2_X1 U407 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n343) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U409 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U410 ( .A(n344), .B(KEYINPUT75), .Z(n349) );
  XOR2_X1 U411 ( .A(KEYINPUT73), .B(G211GAT), .Z(n346) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(G183GAT), .ZN(n345) );
  XNOR2_X1 U413 ( .A(n346), .B(n345), .ZN(n387) );
  XNOR2_X1 U414 ( .A(n347), .B(n387), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U416 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n351) );
  XNOR2_X1 U417 ( .A(G155GAT), .B(G64GAT), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U419 ( .A(n353), .B(n352), .Z(n358) );
  XOR2_X1 U420 ( .A(G1GAT), .B(G127GAT), .Z(n354) );
  XNOR2_X1 U421 ( .A(G57GAT), .B(n354), .ZN(n381) );
  INV_X1 U422 ( .A(n381), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n582) );
  XNOR2_X1 U425 ( .A(G155GAT), .B(KEYINPUT81), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n359), .B(KEYINPUT2), .ZN(n360) );
  XOR2_X1 U427 ( .A(n360), .B(KEYINPUT3), .Z(n362) );
  XNOR2_X1 U428 ( .A(G141GAT), .B(G162GAT), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n362), .B(n361), .ZN(n429) );
  XNOR2_X1 U430 ( .A(n429), .B(KEYINPUT4), .ZN(n365) );
  XOR2_X1 U431 ( .A(KEYINPUT85), .B(KEYINPUT89), .Z(n364) );
  XNOR2_X1 U432 ( .A(G85GAT), .B(KEYINPUT88), .ZN(n363) );
  XOR2_X1 U433 ( .A(KEYINPUT1), .B(KEYINPUT86), .Z(n367) );
  XNOR2_X1 U434 ( .A(KEYINPUT84), .B(KEYINPUT87), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n371) );
  NAND2_X1 U436 ( .A1(G225GAT), .A2(G233GAT), .ZN(n369) );
  XOR2_X1 U437 ( .A(n372), .B(KEYINPUT5), .Z(n373) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U440 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n380) );
  XNOR2_X1 U441 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n380), .B(n379), .ZN(n404) );
  XNOR2_X1 U443 ( .A(KEYINPUT90), .B(n440), .ZN(n570) );
  XOR2_X1 U444 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n385) );
  XNOR2_X1 U445 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n403) );
  XNOR2_X1 U447 ( .A(n403), .B(n386), .ZN(n395) );
  XOR2_X1 U448 ( .A(G197GAT), .B(KEYINPUT21), .Z(n415) );
  XOR2_X1 U449 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n390) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U452 ( .A(n415), .B(n391), .Z(n393) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U455 ( .A(n395), .B(n394), .Z(n522) );
  XNOR2_X1 U456 ( .A(n522), .B(KEYINPUT27), .ZN(n437) );
  NOR2_X1 U457 ( .A1(n570), .A2(n437), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n396), .B(KEYINPUT93), .ZN(n533) );
  XOR2_X1 U459 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n398) );
  XNOR2_X1 U460 ( .A(KEYINPUT20), .B(KEYINPUT78), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n414) );
  XOR2_X1 U462 ( .A(G183GAT), .B(G134GAT), .Z(n400) );
  XNOR2_X1 U463 ( .A(G43GAT), .B(G15GAT), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U465 ( .A(G190GAT), .B(G99GAT), .Z(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U468 ( .A(G120GAT), .B(G127GAT), .Z(n406) );
  XNOR2_X1 U469 ( .A(G71GAT), .B(G176GAT), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n412) );
  NAND2_X1 U473 ( .A1(G227GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n524) );
  INV_X1 U476 ( .A(n524), .ZN(n535) );
  NOR2_X1 U477 ( .A1(n533), .A2(n535), .ZN(n432) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n418) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n419), .B(G211GAT), .Z(n424) );
  XOR2_X1 U482 ( .A(G78GAT), .B(G148GAT), .Z(n421) );
  XNOR2_X1 U483 ( .A(KEYINPUT82), .B(G204GAT), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n422), .B(G218GAT), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U487 ( .A(KEYINPUT22), .B(KEYINPUT83), .Z(n426) );
  NAND2_X1 U488 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n431) );
  XNOR2_X1 U491 ( .A(G22GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n470) );
  XNOR2_X1 U493 ( .A(n470), .B(KEYINPUT28), .ZN(n538) );
  INV_X1 U494 ( .A(n538), .ZN(n529) );
  NAND2_X1 U495 ( .A1(n432), .A2(n529), .ZN(n443) );
  NOR2_X1 U496 ( .A1(n524), .A2(n522), .ZN(n433) );
  NOR2_X1 U497 ( .A1(n470), .A2(n433), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n434), .B(KEYINPUT25), .ZN(n439) );
  XOR2_X1 U499 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n436) );
  NAND2_X1 U500 ( .A1(n470), .A2(n524), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n550) );
  INV_X1 U502 ( .A(n550), .ZN(n572) );
  OR2_X1 U503 ( .A1(n572), .A2(n437), .ZN(n438) );
  NAND2_X1 U504 ( .A1(n439), .A2(n438), .ZN(n441) );
  NAND2_X1 U505 ( .A1(n441), .A2(n440), .ZN(n442) );
  NAND2_X1 U506 ( .A1(n443), .A2(n442), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n444), .B(KEYINPUT95), .ZN(n486) );
  NOR2_X1 U508 ( .A1(n582), .A2(n486), .ZN(n445) );
  NAND2_X1 U509 ( .A1(n584), .A2(n445), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n446), .B(KEYINPUT37), .ZN(n518) );
  NAND2_X1 U511 ( .A1(n487), .A2(n518), .ZN(n447) );
  NOR2_X1 U512 ( .A1(n503), .A2(n524), .ZN(n452) );
  XNOR2_X1 U513 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n450) );
  XOR2_X1 U514 ( .A(KEYINPUT41), .B(n578), .Z(n556) );
  NAND2_X1 U515 ( .A1(n556), .A2(n574), .ZN(n454) );
  XOR2_X1 U516 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n453) );
  XNOR2_X1 U517 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X1 U518 ( .A1(n561), .A2(n455), .ZN(n456) );
  XNOR2_X1 U519 ( .A(KEYINPUT111), .B(n582), .ZN(n568) );
  NAND2_X1 U520 ( .A1(n456), .A2(n568), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n457), .B(KEYINPUT113), .ZN(n458) );
  XNOR2_X1 U522 ( .A(n458), .B(KEYINPUT47), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n584), .A2(n582), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n459), .B(KEYINPUT114), .ZN(n460) );
  XNOR2_X1 U525 ( .A(n460), .B(KEYINPUT45), .ZN(n461) );
  NOR2_X1 U526 ( .A1(n578), .A2(n461), .ZN(n462) );
  NAND2_X1 U527 ( .A1(n462), .A2(n506), .ZN(n463) );
  NAND2_X1 U528 ( .A1(n464), .A2(n463), .ZN(n466) );
  XOR2_X1 U529 ( .A(n522), .B(KEYINPUT121), .Z(n467) );
  NOR2_X1 U530 ( .A1(n534), .A2(n467), .ZN(n469) );
  INV_X1 U531 ( .A(n470), .ZN(n471) );
  AND2_X1 U532 ( .A1(n570), .A2(n471), .ZN(n472) );
  AND2_X1 U533 ( .A1(n571), .A2(n472), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT124), .B(KEYINPUT55), .ZN(n474) );
  INV_X1 U535 ( .A(KEYINPUT123), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n524), .A2(n477), .ZN(n566) );
  NAND2_X1 U537 ( .A1(n566), .A2(n561), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n566), .A2(n556), .ZN(n482) );
  XOR2_X1 U539 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(G176GAT), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(G1349GAT) );
  INV_X1 U542 ( .A(n582), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n561), .A2(n483), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n507) );
  NAND2_X1 U546 ( .A1(n487), .A2(n507), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT96), .B(n488), .ZN(n496) );
  NOR2_X1 U548 ( .A1(n570), .A2(n496), .ZN(n489) );
  XOR2_X1 U549 ( .A(G1GAT), .B(n489), .Z(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT34), .B(n490), .ZN(G1324GAT) );
  NOR2_X1 U551 ( .A1(n496), .A2(n522), .ZN(n491) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n491), .Z(G1325GAT) );
  NOR2_X1 U553 ( .A1(n524), .A2(n496), .ZN(n495) );
  XOR2_X1 U554 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n493) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n529), .A2(n496), .ZN(n497) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n497), .Z(G1327GAT) );
  NOR2_X1 U560 ( .A1(n503), .A2(n570), .ZN(n501) );
  XOR2_X1 U561 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n499) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n503), .A2(n522), .ZN(n502) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n505) );
  NOR2_X1 U568 ( .A1(n529), .A2(n503), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  AND2_X1 U570 ( .A1(n506), .A2(n556), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n507), .A2(n517), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n570), .A2(n514), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n510), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n522), .A2(n514), .ZN(n511) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n524), .A2(n514), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n529), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n528) );
  NOR2_X1 U585 ( .A1(n570), .A2(n528), .ZN(n520) );
  XNOR2_X1 U586 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n522), .A2(n528), .ZN(n523) );
  XOR2_X1 U590 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U591 ( .A1(n524), .A2(n528), .ZN(n526) );
  XNOR2_X1 U592 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U596 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U598 ( .A(G106GAT), .B(n532), .Z(G1339GAT) );
  NOR2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n549) );
  NAND2_X1 U600 ( .A1(n535), .A2(n549), .ZN(n536) );
  XOR2_X1 U601 ( .A(KEYINPUT115), .B(n536), .Z(n537) );
  NOR2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n545), .A2(n574), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U606 ( .A1(n545), .A2(n556), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  INV_X1 U608 ( .A(n545), .ZN(n542) );
  NOR2_X1 U609 ( .A1(n568), .A2(n542), .ZN(n543) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n547) );
  NAND2_X1 U613 ( .A1(n545), .A2(n561), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT117), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n574), .A2(n562), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(n555), .Z(n558) );
  NAND2_X1 U624 ( .A1(n562), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n562), .A2(n582), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(KEYINPUT120), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U631 ( .A(G169GAT), .B(KEYINPUT125), .Z(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n574), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  INV_X1 U634 ( .A(n566), .ZN(n567) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n585) );
  NAND2_X1 U640 ( .A1(n585), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

