//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT74), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n204), .B1(G155gat), .B2(G162gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT75), .B(G141gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(new_n208), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT76), .B(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n214), .A3(new_n202), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n207), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n207), .A2(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT3), .ZN(new_n220));
  INV_X1    g019(.A(G113gat), .ZN(new_n221));
  INV_X1    g020(.A(G120gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT1), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n221), .B2(new_n222), .ZN(new_n224));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT77), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n218), .A2(new_n220), .A3(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n207), .A2(new_n215), .A3(new_n226), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT79), .B1(new_n230), .B2(KEYINPUT4), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n230), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n235));
  OAI211_X1 g034(.A(KEYINPUT5), .B(new_n228), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G225gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT5), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n218), .A2(new_n220), .A3(new_n227), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n229), .A2(new_n232), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(KEYINPUT4), .B2(new_n229), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n238), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n219), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT80), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n246), .A3(new_n219), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n230), .A3(new_n247), .ZN(new_n248));
  OR3_X1    g047(.A1(new_n248), .A2(new_n238), .A3(new_n237), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G1gat), .B(G29gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT0), .ZN(new_n252));
  XNOR2_X1  g051(.A(G57gat), .B(G85gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n243), .A2(new_n249), .A3(new_n254), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n250), .A2(KEYINPUT6), .A3(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262));
  INV_X1    g061(.A(G22gat), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  INV_X1    g063(.A(G218gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G197gat), .ZN(new_n267));
  INV_X1    g066(.A(G204gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(G197gat), .A2(G204gat), .ZN(new_n270));
  OAI22_X1  g069(.A1(KEYINPUT22), .A2(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n265), .ZN(new_n272));
  NAND2_X1  g071(.A1(G211gat), .A2(G218gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(KEYINPUT69), .A3(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n271), .B(new_n274), .Z(new_n275));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n218), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT3), .B1(new_n275), .B2(new_n276), .ZN(new_n279));
  OAI211_X1 g078(.A(G228gat), .B(G233gat), .C1(new_n279), .C2(new_n216), .ZN(new_n280));
  OR3_X1    g079(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n277), .B2(new_n280), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT81), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n285), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n286), .A2(new_n273), .A3(new_n272), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n276), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n216), .B1(new_n291), .B2(new_n217), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n284), .B1(new_n277), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n263), .B1(new_n283), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n282), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n277), .A2(new_n280), .A3(new_n278), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n263), .B(new_n293), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n262), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G78gat), .B(G106gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT31), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(G50gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G22gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT83), .A3(new_n297), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n297), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n262), .A3(new_n302), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n314), .A2(new_n315), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n316), .A2(new_n318), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  XOR2_X1   g118(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n320));
  INV_X1    g119(.A(KEYINPUT65), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT27), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT64), .B1(new_n322), .B2(G183gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT27), .B(G183gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n321), .B(new_n323), .C1(new_n324), .C2(KEYINPUT64), .ZN(new_n325));
  INV_X1    g124(.A(G183gat), .ZN(new_n326));
  OR4_X1    g125(.A1(KEYINPUT64), .A2(new_n321), .A3(new_n326), .A4(KEYINPUT27), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n320), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n324), .A2(KEYINPUT28), .A3(new_n329), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n319), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(KEYINPUT24), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(KEYINPUT23), .B2(new_n317), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(new_n329), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(KEYINPUT24), .A3(new_n333), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n317), .A2(KEYINPUT23), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .A4(new_n311), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(new_n226), .ZN(new_n343));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT34), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n346), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G15gat), .B(G43gat), .Z(new_n352));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n343), .A2(new_n344), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(KEYINPUT33), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n355), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n349), .A2(new_n356), .A3(new_n350), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n358), .B2(new_n362), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n342), .A2(G226gat), .A3(G233gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT70), .ZN(new_n367));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n342), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(KEYINPUT29), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n275), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n366), .A2(KEYINPUT71), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n366), .A2(KEYINPUT71), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n275), .B(new_n370), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT72), .ZN(new_n378));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n373), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT73), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT73), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n373), .A2(new_n385), .A3(new_n376), .A4(new_n381), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n373), .B2(new_n376), .ZN(new_n388));
  INV_X1    g187(.A(new_n382), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(KEYINPUT30), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n310), .A2(new_n365), .A3(new_n387), .A4(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n261), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT35), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n358), .A2(new_n362), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n360), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n307), .A3(new_n309), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n390), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT35), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n261), .ZN(new_n401));
  AND4_X1   g200(.A1(new_n260), .A2(new_n259), .A3(new_n383), .A4(new_n386), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT37), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n373), .A2(new_n403), .A3(new_n376), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n380), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n373), .B2(new_n376), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT38), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT86), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n409), .B(KEYINPUT38), .C1(new_n405), .C2(new_n406), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n403), .B1(new_n371), .B2(new_n275), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n275), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT38), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n380), .A4(new_n404), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n402), .A2(new_n408), .A3(new_n410), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n307), .A2(new_n309), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n254), .B1(new_n243), .B2(new_n249), .ZN(new_n418));
  XOR2_X1   g217(.A(KEYINPUT84), .B(KEYINPUT40), .Z(new_n419));
  INV_X1    g218(.A(new_n237), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n239), .B2(new_n241), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT39), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n255), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n421), .B(KEYINPUT39), .C1(new_n248), .C2(new_n420), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n419), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(KEYINPUT40), .A3(new_n425), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT85), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT40), .A4(new_n425), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n418), .B(new_n426), .C1(new_n428), .C2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n417), .B1(new_n398), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n261), .A2(new_n387), .A3(new_n390), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT36), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n363), .B2(new_n364), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n395), .A2(KEYINPUT36), .A3(new_n396), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n417), .A2(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n393), .A2(new_n401), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G113gat), .B(G141gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT88), .ZN(new_n441));
  XOR2_X1   g240(.A(G169gat), .B(G197gat), .Z(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT12), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G15gat), .B(G22gat), .ZN(new_n448));
  INV_X1    g247(.A(G1gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT16), .A3(new_n449), .ZN(new_n450));
  OR2_X1    g249(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n450), .B(new_n451), .C1(new_n449), .C2(new_n448), .ZN(new_n452));
  NAND2_X1  g251(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(G43gat), .B(G50gat), .Z(new_n456));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G29gat), .A2(G36gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n457), .ZN(new_n460));
  OR3_X1    g259(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n465), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n461), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n468), .A2(new_n459), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n464), .B1(new_n469), .B2(new_n458), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n464), .B(KEYINPUT17), .C1(new_n469), .C2(new_n458), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n470), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT18), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n474), .A2(KEYINPUT18), .A3(new_n475), .A4(new_n476), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n454), .B(new_n470), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n475), .B(KEYINPUT13), .Z(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n447), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n447), .A2(new_n484), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n439), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT101), .ZN(new_n490));
  XNOR2_X1  g289(.A(G120gat), .B(G148gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n495));
  XNOR2_X1  g294(.A(G99gat), .B(G106gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT7), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(G85gat), .A3(G92gat), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT8), .ZN(new_n503));
  INV_X1    g302(.A(G85gat), .ZN(new_n504));
  INV_X1    g303(.A(G92gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n495), .B(new_n496), .C1(new_n501), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n496), .A2(new_n495), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n498), .A2(new_n500), .ZN(new_n510));
  OR2_X1    g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(KEYINPUT95), .A3(new_n502), .ZN(new_n512));
  AOI22_X1  g311(.A1(KEYINPUT8), .A2(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n509), .A2(new_n510), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G57gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G64gat), .ZN(new_n517));
  INV_X1    g316(.A(G64gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G57gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G71gat), .B(G78gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT9), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G71gat), .ZN(new_n526));
  INV_X1    g325(.A(G78gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT92), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G71gat), .B2(G78gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(G71gat), .A3(G78gat), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(new_n529), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n517), .A2(new_n519), .B1(new_n523), .B2(new_n522), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n525), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n515), .A2(new_n537), .A3(KEYINPUT10), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n515), .A2(new_n537), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT10), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(new_n508), .A3(new_n514), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n515), .A2(new_n537), .A3(KEYINPUT97), .A4(KEYINPUT10), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT100), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT100), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n541), .A2(new_n543), .ZN(new_n553));
  INV_X1    g352(.A(new_n547), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n494), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT98), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n558), .A3(new_n554), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n559), .A2(new_n493), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(KEYINPUT98), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n548), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT99), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT99), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n560), .A2(new_n548), .A3(new_n564), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n557), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n472), .A2(new_n473), .A3(new_n508), .A4(new_n514), .ZN(new_n569));
  AND2_X1   g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n470), .A2(new_n515), .B1(KEYINPUT41), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n575));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT96), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n577), .A2(KEYINPUT96), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n455), .B1(new_n583), .B2(new_n536), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n536), .A2(new_n583), .ZN(new_n585));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT93), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT94), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n588), .B(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n568), .A2(new_n582), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n489), .A2(new_n490), .A3(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n416), .A2(new_n432), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n434), .A2(new_n417), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n436), .A2(new_n437), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n400), .B1(new_n399), .B2(new_n261), .ZN(new_n604));
  NOR4_X1   g403(.A1(new_n397), .A2(new_n398), .A3(new_n392), .A4(KEYINPUT35), .ZN(new_n605));
  OAI22_X1  g404(.A1(new_n600), .A2(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n487), .A3(new_n598), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT101), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n261), .B1(new_n599), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n449), .ZN(G1324gat));
  INV_X1    g409(.A(KEYINPUT42), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT102), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT16), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n490), .B1(new_n489), .B2(new_n598), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n607), .A2(KEYINPUT101), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n398), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(G8gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n608), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n398), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n611), .ZN(new_n620));
  INV_X1    g419(.A(G8gat), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n618), .A2(new_n621), .A3(new_n398), .A4(new_n613), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n620), .A3(new_n622), .ZN(G1325gat));
  INV_X1    g422(.A(G15gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n624), .A3(new_n365), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n602), .B1(new_n599), .B2(new_n608), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(new_n624), .B2(new_n626), .ZN(G1326gat));
  AOI21_X1  g426(.A(new_n310), .B1(new_n599), .B2(new_n608), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT43), .B(G22gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(G1327gat));
  INV_X1    g430(.A(new_n582), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n567), .A2(new_n596), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT103), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n606), .A2(new_n487), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G29gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(new_n392), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT45), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n439), .B2(new_n582), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n604), .A2(new_n605), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n603), .B1(new_n416), .B2(new_n432), .ZN(new_n643));
  OAI211_X1 g442(.A(KEYINPUT44), .B(new_n632), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645));
  INV_X1    g444(.A(new_n486), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n447), .A2(new_n484), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n485), .A2(KEYINPUT104), .A3(new_n486), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n633), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT105), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n641), .A2(new_n644), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G29gat), .B1(new_n653), .B2(new_n261), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n654), .ZN(G1328gat));
  INV_X1    g454(.A(new_n398), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(G36gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n641), .A2(new_n644), .A3(new_n398), .A4(new_n652), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(G36gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(G1329gat));
  INV_X1    g465(.A(new_n602), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n641), .A2(new_n644), .A3(new_n667), .A4(new_n652), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(G43gat), .ZN(new_n669));
  INV_X1    g468(.A(G43gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n636), .A2(new_n670), .A3(new_n365), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT47), .B1(new_n671), .B2(KEYINPUT107), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n669), .B(new_n671), .C1(KEYINPUT107), .C2(KEYINPUT47), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(G1330gat));
  NOR2_X1   g475(.A1(new_n310), .A2(G50gat), .ZN(new_n677));
  AND4_X1   g476(.A1(new_n487), .A2(new_n606), .A3(new_n635), .A4(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n641), .A2(new_n644), .A3(new_n417), .A4(new_n652), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(G50gat), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT48), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI211_X1 g481(.A(KEYINPUT48), .B(new_n678), .C1(new_n679), .C2(G50gat), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(G1331gat));
  INV_X1    g483(.A(new_n596), .ZN(new_n685));
  NOR4_X1   g484(.A1(new_n650), .A2(new_n632), .A3(new_n685), .A4(new_n568), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n606), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n261), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(new_n516), .ZN(G1332gat));
  AOI211_X1 g488(.A(new_n656), .B(new_n687), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1333gat));
  OAI21_X1  g491(.A(G71gat), .B1(new_n687), .B2(new_n602), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n365), .A2(new_n526), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n687), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1334gat));
  NOR2_X1   g496(.A1(new_n687), .A2(new_n310), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(new_n527), .ZN(G1335gat));
  NOR2_X1   g498(.A1(new_n439), .A2(new_n582), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT51), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n650), .A2(new_n596), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n700), .A2(KEYINPUT110), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n606), .A2(new_n632), .A3(new_n702), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n701), .A2(KEYINPUT110), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(KEYINPUT110), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n261), .A2(G85gat), .A3(new_n568), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n650), .A2(new_n596), .A3(new_n568), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n641), .A2(new_n644), .A3(new_n392), .A4(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G85gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n711), .A2(new_n712), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n709), .B1(new_n714), .B2(new_n715), .ZN(G1336gat));
  NOR3_X1   g515(.A1(new_n656), .A2(G92gat), .A3(new_n568), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n703), .A2(new_n707), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n641), .A2(new_n644), .A3(new_n398), .A4(new_n710), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G92gat), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n704), .A2(new_n723), .A3(new_n701), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n701), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n700), .A2(new_n702), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n727), .A2(new_n717), .B1(G92gat), .B2(new_n719), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n722), .B1(new_n728), .B2(new_n721), .ZN(G1337gat));
  NOR2_X1   g528(.A1(new_n568), .A2(G99gat), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n703), .A2(new_n707), .A3(new_n365), .A4(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n641), .A2(new_n644), .A3(new_n710), .ZN(new_n732));
  OAI21_X1  g531(.A(G99gat), .B1(new_n732), .B2(new_n602), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1338gat));
  NOR3_X1   g533(.A1(new_n310), .A2(G106gat), .A3(new_n568), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n703), .A2(new_n707), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n641), .A2(new_n644), .A3(new_n417), .A4(new_n710), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G106gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT53), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n727), .A2(new_n735), .B1(G106gat), .B2(new_n737), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n739), .ZN(G1339gat));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n549), .A2(new_n743), .A3(new_n551), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n546), .B2(new_n547), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n540), .A2(new_n544), .A3(new_n545), .A4(new_n554), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n493), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n744), .A2(KEYINPUT55), .A3(new_n747), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(new_n566), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n747), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI211_X1 g552(.A(KEYINPUT113), .B(KEYINPUT55), .C1(new_n744), .C2(new_n747), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n749), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT114), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n749), .B(new_n757), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n650), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n481), .A2(new_n482), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT115), .Z(new_n761));
  AOI21_X1  g560(.A(new_n475), .B1(new_n474), .B2(new_n476), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n445), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n567), .A3(new_n485), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n632), .B1(new_n759), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n632), .A2(new_n485), .A3(new_n763), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n766), .A2(new_n756), .A3(new_n758), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n685), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n650), .A2(new_n597), .A3(KEYINPUT112), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT112), .B1(new_n650), .B2(new_n597), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n261), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n399), .ZN(new_n774));
  AOI21_X1  g573(.A(G113gat), .B1(new_n774), .B2(new_n650), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n488), .A2(new_n221), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(G1340gat));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n567), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g578(.A1(new_n774), .A2(new_n596), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G127gat), .ZN(G1342gat));
  INV_X1    g580(.A(G134gat), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n773), .A2(new_n782), .A3(new_n399), .A4(new_n632), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT116), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n784), .A2(KEYINPUT56), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(KEYINPUT56), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n774), .A2(new_n632), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n785), .B(new_n786), .C1(new_n782), .C2(new_n787), .ZN(G1343gat));
  NOR2_X1   g587(.A1(new_n398), .A2(new_n261), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n602), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n602), .A2(new_n789), .A3(KEYINPUT117), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n766), .A2(new_n756), .A3(new_n758), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n751), .A2(new_n752), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n487), .A2(new_n749), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n764), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n582), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n596), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n417), .B1(new_n800), .B2(new_n771), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n794), .B1(KEYINPUT57), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n310), .B1(new_n768), .B2(new_n772), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n210), .B1(new_n806), .B2(new_n488), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n667), .A2(new_n310), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n773), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n773), .A2(KEYINPUT118), .A3(new_n810), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n656), .A3(new_n814), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n488), .A2(G141gat), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n811), .A2(new_n398), .A3(new_n816), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n805), .A3(new_n650), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n210), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n809), .A2(new_n817), .B1(new_n808), .B2(new_n820), .ZN(G1344gat));
  INV_X1    g620(.A(new_n815), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n208), .A3(new_n567), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n806), .A2(new_n568), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(KEYINPUT59), .A3(new_n208), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n803), .A2(new_n804), .ZN(new_n827));
  INV_X1    g626(.A(new_n794), .ZN(new_n828));
  INV_X1    g627(.A(new_n755), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n766), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n596), .B1(new_n830), .B2(new_n799), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n597), .A2(new_n487), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n804), .B(new_n417), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n827), .A2(new_n567), .A3(new_n828), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n826), .B1(new_n834), .B2(G148gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n823), .B1(new_n825), .B2(new_n835), .ZN(G1345gat));
  OAI21_X1  g635(.A(G155gat), .B1(new_n806), .B2(new_n685), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n596), .A2(new_n213), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n815), .B2(new_n838), .ZN(G1346gat));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n212), .A3(new_n632), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n806), .B2(new_n582), .ZN(new_n842));
  INV_X1    g641(.A(new_n212), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n806), .A2(new_n841), .A3(new_n582), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(G1347gat));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n656), .A2(new_n397), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n759), .A2(new_n764), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n582), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n596), .B1(new_n850), .B2(new_n795), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n261), .B(new_n848), .C1(new_n851), .C2(new_n771), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n392), .B1(new_n768), .B2(new_n772), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n855), .A3(new_n848), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n487), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G169gat), .ZN(new_n859));
  INV_X1    g658(.A(new_n650), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n852), .A2(G169gat), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n847), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g662(.A(KEYINPUT121), .B(new_n861), .C1(new_n858), .C2(G169gat), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(G1348gat));
  INV_X1    g664(.A(new_n852), .ZN(new_n866));
  INV_X1    g665(.A(G176gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n567), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n568), .B1(new_n853), .B2(new_n856), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n867), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT122), .ZN(G1349gat));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT60), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(KEYINPUT60), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n326), .B1(new_n857), .B2(new_n596), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n596), .A2(new_n324), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n854), .A2(new_n848), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n877), .B(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n879), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n854), .A2(new_n855), .A3(new_n848), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n855), .B1(new_n854), .B2(new_n848), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n596), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G183gat), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n877), .B(KEYINPUT123), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n884), .A2(new_n872), .A3(KEYINPUT60), .A4(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n880), .A2(new_n886), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n866), .A2(new_n329), .A3(new_n632), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n329), .B1(new_n857), .B2(new_n632), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(G1351gat));
  AND3_X1   g692(.A1(new_n854), .A2(new_n398), .A3(new_n810), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(new_n650), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n667), .A2(new_n392), .A3(new_n656), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n833), .B(new_n896), .C1(new_n803), .C2(new_n804), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n487), .A2(G197gat), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n895), .A2(G197gat), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(G1352gat));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n268), .A3(new_n567), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT62), .Z(new_n902));
  NAND3_X1  g701(.A1(new_n827), .A2(new_n567), .A3(new_n833), .ZN(new_n903));
  INV_X1    g702(.A(new_n896), .ZN(new_n904));
  OAI21_X1  g703(.A(G204gat), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(G1353gat));
  NAND3_X1  g705(.A1(new_n894), .A2(new_n264), .A3(new_n596), .ZN(new_n907));
  INV_X1    g706(.A(new_n897), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n596), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT63), .B1(new_n909), .B2(G211gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(G1354gat));
  AOI21_X1  g712(.A(G218gat), .B1(new_n894), .B2(new_n632), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n632), .A2(G218gat), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT126), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n915), .A2(new_n916), .B1(new_n908), .B2(new_n918), .ZN(G1355gat));
endmodule


