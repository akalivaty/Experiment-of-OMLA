//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G140), .Z(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT83), .ZN(new_n190));
  INV_X1    g004(.A(G227), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  XOR2_X1   g006(.A(new_n190), .B(new_n192), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT0), .B(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n197), .B2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n195), .A2(KEYINPUT64), .A3(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT65), .B1(new_n195), .B2(G143), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n197), .A3(G146), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n205), .A2(new_n207), .A3(new_n208), .A4(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n208), .A2(new_n210), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n214), .A2(KEYINPUT66), .A3(new_n207), .A4(new_n205), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n201), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT3), .B1(new_n217), .B2(G107), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G101), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(G101), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n218), .A2(new_n221), .A3(new_n227), .A4(new_n222), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n216), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n214), .A2(new_n231), .A3(G128), .A4(new_n205), .ZN(new_n232));
  OAI21_X1  g046(.A(G128), .B1(new_n198), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n196), .B2(new_n198), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n222), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n217), .A2(G107), .ZN(new_n237));
  OAI21_X1  g051(.A(G101), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n238), .A2(new_n228), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(KEYINPUT10), .A3(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n195), .A2(KEYINPUT64), .A3(G143), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT64), .B1(new_n195), .B2(G143), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n208), .B(new_n210), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n233), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT84), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(KEYINPUT84), .A3(new_n233), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n232), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n239), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT85), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT85), .ZN(new_n252));
  AOI211_X1 g066(.A(new_n252), .B(KEYINPUT10), .C1(new_n248), .C2(new_n239), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n230), .B(new_n240), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT87), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n239), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n243), .A2(KEYINPUT84), .A3(new_n233), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT84), .B1(new_n243), .B2(new_n233), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n257), .B1(new_n260), .B2(new_n232), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n252), .B1(new_n261), .B2(KEYINPUT10), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n249), .A2(KEYINPUT85), .A3(new_n250), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n264), .A2(KEYINPUT87), .A3(new_n230), .A4(new_n240), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT11), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n266), .A2(new_n267), .A3(G137), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n266), .B1(new_n267), .B2(G137), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G131), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n267), .A2(G137), .ZN(new_n273));
  OAI211_X1 g087(.A(KEYINPUT67), .B(new_n266), .C1(new_n267), .C2(G137), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n271), .A2(new_n272), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n269), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n267), .A2(G137), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT11), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n276), .A2(new_n278), .A3(new_n273), .A4(new_n274), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G131), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n256), .A2(new_n265), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n254), .A2(new_n281), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n194), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n257), .A2(new_n234), .A3(new_n232), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n249), .A2(new_n286), .B1(new_n280), .B2(new_n275), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n287), .A2(KEYINPUT86), .A3(KEYINPUT12), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT86), .B1(new_n287), .B2(KEYINPUT12), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n287), .A2(KEYINPUT12), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n194), .B1(new_n254), .B2(new_n281), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n187), .B(new_n188), .C1(new_n285), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(G469), .A2(G902), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n284), .A3(new_n194), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n193), .B1(new_n291), .B2(new_n283), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(G469), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(G125), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n232), .A2(new_n301), .A3(new_n234), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n213), .A2(new_n215), .ZN(new_n303));
  INV_X1    g117(.A(new_n201), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT89), .B1(new_n305), .B2(G125), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT89), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n216), .A2(new_n307), .A3(new_n301), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n302), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT90), .B(G224), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G953), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n311), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n302), .B(new_n313), .C1(new_n306), .C2(new_n308), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(G110), .B(G122), .Z(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT2), .B(G113), .ZN(new_n318));
  INV_X1    g132(.A(G119), .ZN(new_n319));
  OR2_X1    g133(.A1(KEYINPUT69), .A2(G116), .ZN(new_n320));
  NAND2_X1  g134(.A1(KEYINPUT69), .A2(G116), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(G116), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n318), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n318), .ZN(new_n326));
  AND2_X1   g140(.A1(KEYINPUT69), .A2(G116), .ZN(new_n327));
  NOR2_X1   g141(.A1(KEYINPUT69), .A2(G116), .ZN(new_n328));
  OAI21_X1  g142(.A(G119), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n329), .A3(new_n323), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n229), .A3(new_n225), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(KEYINPUT5), .A3(new_n323), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(G113), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n239), .A3(new_n330), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n317), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n337), .A2(KEYINPUT6), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n332), .A2(new_n336), .A3(new_n317), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT88), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT88), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n332), .A2(new_n336), .A3(new_n341), .A4(new_n317), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n337), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n315), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G210), .B1(G237), .B2(G902), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n302), .B1(new_n216), .B2(new_n301), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n313), .A2(KEYINPUT7), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n335), .A2(new_n330), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n257), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n336), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n316), .B(KEYINPUT8), .Z(new_n353));
  AOI22_X1  g167(.A1(new_n348), .A2(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n340), .A2(new_n342), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n313), .A2(KEYINPUT91), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n302), .B(new_n356), .C1(new_n306), .C2(new_n308), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT7), .B1(new_n313), .B2(KEYINPUT91), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n354), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  AND4_X1   g173(.A1(new_n188), .A2(new_n346), .A3(new_n347), .A4(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n315), .B2(new_n345), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n347), .B1(new_n361), .B2(new_n359), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n300), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G113), .B(G122), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(new_n217), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n301), .A2(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT16), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT75), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G125), .B(G140), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT16), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n367), .B2(KEYINPUT16), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n370), .A2(new_n366), .A3(KEYINPUT76), .A4(G125), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n195), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n371), .A2(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G146), .ZN(new_n383));
  NOR2_X1   g197(.A1(G237), .A2(G953), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n197), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(G143), .A3(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT17), .A3(G131), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(G131), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT17), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n272), .A3(new_n387), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n381), .A2(new_n383), .A3(new_n389), .A4(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n372), .B(new_n195), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n272), .ZN(new_n397));
  OAI221_X1 g211(.A(new_n395), .B1(new_n388), .B2(new_n397), .C1(new_n390), .C2(new_n396), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n365), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT92), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n394), .A2(new_n365), .A3(new_n398), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n400), .B(new_n188), .C1(new_n403), .C2(new_n399), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G475), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n390), .A2(new_n392), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n369), .A2(KEYINPUT19), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n369), .A2(KEYINPUT19), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n195), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n383), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n398), .ZN(new_n411));
  INV_X1    g225(.A(new_n365), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(G475), .B1(new_n413), .B2(new_n401), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n188), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(KEYINPUT20), .A3(new_n188), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n405), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G953), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G952), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(G234), .B2(G237), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT21), .B(G898), .Z(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(G234), .A2(G237), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(G902), .A3(G953), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G122), .B1(new_n327), .B2(new_n328), .ZN(new_n431));
  INV_X1    g245(.A(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G116), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n431), .A2(new_n435), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(G107), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n220), .ZN(new_n439));
  XNOR2_X1  g253(.A(G128), .B(G143), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(new_n267), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(KEYINPUT13), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n197), .A2(G128), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n443), .B(G134), .C1(KEYINPUT13), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n267), .ZN(new_n446));
  INV_X1    g260(.A(new_n439), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n434), .A2(new_n220), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n445), .B(new_n446), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n442), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT9), .B(G234), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G217), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n452), .A2(new_n453), .A3(G953), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n442), .A2(new_n449), .A3(new_n454), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G478), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n459), .A2(KEYINPUT15), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n188), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n458), .B2(new_n188), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n420), .A2(new_n430), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n363), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G221), .B1(new_n452), .B2(G902), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n299), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n421), .A2(G221), .A3(G234), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(G137), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n381), .A2(new_n383), .ZN(new_n474));
  INV_X1    g288(.A(G128), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G119), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT74), .ZN(new_n477));
  AND2_X1   g291(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n478));
  NOR2_X1   g292(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n319), .A2(G128), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g296(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n484));
  AND4_X1   g298(.A1(new_n477), .A2(new_n483), .A3(new_n481), .A4(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n476), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n476), .A2(KEYINPUT23), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(G110), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n476), .A2(new_n481), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT24), .B(G110), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n474), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n369), .A2(G146), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n382), .B2(G146), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT77), .B(G110), .Z(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n486), .B2(new_n488), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(new_n491), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT78), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n494), .B(KEYINPUT79), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n495), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n483), .A2(new_n481), .A3(new_n484), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT74), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n480), .A2(new_n477), .A3(new_n481), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n503), .A2(new_n504), .B1(G119), .B2(new_n475), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n501), .B1(new_n505), .B2(new_n487), .ZN(new_n506));
  INV_X1    g320(.A(new_n498), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT79), .B1(new_n508), .B2(new_n494), .ZN(new_n509));
  OAI211_X1 g323(.A(KEYINPUT80), .B(new_n492), .C1(new_n500), .C2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT79), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n499), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT80), .B1(new_n515), .B2(new_n492), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n473), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n473), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n492), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n188), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT25), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n453), .B1(G234), .B2(new_n188), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n517), .A2(new_n523), .A3(new_n188), .A4(new_n519), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n517), .A2(new_n519), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n522), .A2(G902), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT68), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n216), .A2(new_n281), .ZN(new_n534));
  INV_X1    g348(.A(new_n273), .ZN(new_n535));
  OAI21_X1  g349(.A(G131), .B1(new_n535), .B2(new_n277), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n235), .A2(new_n275), .A3(new_n536), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(new_n537), .ZN(new_n538));
  AND4_X1   g352(.A1(new_n530), .A2(new_n534), .A3(new_n531), .A4(new_n537), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n331), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n331), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n543), .A3(new_n537), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n534), .A2(new_n537), .ZN(new_n545));
  INV_X1    g359(.A(new_n532), .ZN(new_n546));
  INV_X1    g360(.A(new_n533), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n534), .A2(new_n537), .A3(new_n530), .A4(new_n531), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT70), .A3(new_n331), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n544), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n384), .A2(G210), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n227), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n554), .B(new_n555), .Z(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n559));
  INV_X1    g373(.A(new_n544), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n543), .B1(new_n534), .B2(new_n537), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT28), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT71), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n544), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(KEYINPUT71), .A3(KEYINPUT28), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n544), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n556), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n558), .A2(new_n559), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n562), .A2(KEYINPUT29), .A3(new_n556), .A4(new_n570), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n558), .A2(KEYINPUT72), .A3(new_n571), .A4(new_n559), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n574), .A2(new_n188), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G472), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n556), .B1(new_n568), .B2(new_n570), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n542), .A2(new_n556), .A3(new_n544), .A4(new_n551), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT31), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT32), .ZN(new_n586));
  NOR2_X1   g400(.A1(G472), .A2(G902), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT70), .B1(new_n550), .B2(new_n331), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n541), .B(new_n543), .C1(new_n548), .C2(new_n549), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n591), .A2(KEYINPUT31), .A3(new_n556), .A4(new_n544), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n581), .A2(new_n582), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n579), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n587), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT32), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n529), .B1(new_n578), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT82), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(G472), .A2(new_n577), .B1(new_n588), .B2(new_n596), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n601), .A2(KEYINPUT82), .A3(new_n529), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n469), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  OAI21_X1  g418(.A(G472), .B1(new_n594), .B2(G902), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n585), .A2(new_n587), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n525), .A4(new_n528), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n299), .A2(new_n467), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n363), .A2(KEYINPUT93), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n346), .A2(new_n188), .A3(new_n359), .ZN(new_n611));
  INV_X1    g425(.A(new_n347), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n361), .A2(new_n347), .A3(new_n359), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n300), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n457), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n454), .B1(new_n442), .B2(new_n449), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT33), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n456), .B2(new_n457), .ZN(new_n623));
  OAI211_X1 g437(.A(G478), .B(new_n188), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT94), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n458), .A2(KEYINPUT33), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n456), .A2(new_n622), .A3(new_n457), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n628), .A2(new_n629), .A3(G478), .A4(new_n188), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n619), .A2(new_n620), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n459), .B1(new_n631), .B2(G902), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n625), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n419), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n618), .A2(new_n429), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n609), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT34), .B(G104), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  INV_X1    g453(.A(new_n464), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n420), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n618), .A2(new_n429), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n609), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n644), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n605), .A2(new_n606), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n511), .A2(new_n516), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n473), .A2(KEYINPUT36), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n527), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n525), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n468), .A2(new_n649), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT37), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  AOI21_X1  g473(.A(new_n656), .B1(new_n578), .B2(new_n597), .ZN(new_n660));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n423), .B1(new_n428), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n641), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n608), .A2(new_n618), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  XOR2_X1   g480(.A(new_n615), .B(KEYINPUT38), .Z(new_n667));
  INV_X1    g481(.A(new_n300), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n640), .A2(new_n419), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n655), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT97), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(KEYINPUT97), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n662), .B(KEYINPUT39), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n608), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n552), .A2(new_n556), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n188), .B1(new_n566), .B2(new_n556), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n597), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n673), .A2(new_n676), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  INV_X1    g497(.A(new_n634), .ZN(new_n684));
  INV_X1    g498(.A(new_n662), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n660), .A2(new_n684), .A3(new_n685), .A4(new_n664), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NAND2_X1  g501(.A1(new_n282), .A2(new_n284), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n293), .B1(new_n688), .B2(new_n193), .ZN(new_n689));
  OAI21_X1  g503(.A(G469), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n467), .A3(new_n294), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT98), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n690), .A2(KEYINPUT98), .A3(new_n467), .A4(new_n294), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n598), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n635), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND3_X1  g513(.A1(new_n598), .A2(new_n695), .A3(new_n642), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  INV_X1    g515(.A(new_n465), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n690), .A2(new_n467), .A3(new_n294), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n610), .A2(new_n617), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT99), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT99), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n691), .A2(new_n618), .A3(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n702), .B(new_n660), .C1(new_n705), .C2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NAND2_X1  g523(.A1(new_n562), .A2(new_n570), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n557), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n583), .B2(new_n584), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n587), .B(KEYINPUT100), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(G472), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n585), .B2(new_n188), .ZN(new_n717));
  NOR4_X1   g531(.A1(new_n715), .A2(new_n717), .A3(new_n529), .A4(new_n669), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n430), .A3(new_n704), .A4(new_n695), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NAND3_X1  g534(.A1(new_n633), .A2(new_n419), .A3(new_n685), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT102), .Z(new_n722));
  NAND3_X1  g536(.A1(new_n605), .A2(new_n714), .A3(new_n655), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT101), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n605), .A2(new_n714), .A3(new_n655), .A4(KEYINPUT101), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n722), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT99), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n706), .B1(new_n691), .B2(new_n618), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  INV_X1    g546(.A(new_n722), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n615), .A2(new_n668), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n608), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n598), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n598), .A2(new_n733), .A3(new_n736), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT104), .B(G131), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G33));
  AND3_X1   g558(.A1(new_n598), .A2(new_n663), .A3(new_n736), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n267), .ZN(G36));
  NAND2_X1  g560(.A1(new_n633), .A2(new_n420), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n649), .A2(new_n749), .A3(new_n655), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n735), .B1(new_n751), .B2(KEYINPUT44), .ZN(new_n752));
  INV_X1    g566(.A(new_n674), .ZN(new_n753));
  INV_X1    g567(.A(new_n467), .ZN(new_n754));
  INV_X1    g568(.A(new_n294), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n296), .A2(new_n297), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n296), .A2(KEYINPUT45), .A3(new_n297), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(G469), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n295), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n755), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(KEYINPUT46), .A3(new_n295), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n754), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n750), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n752), .A2(new_n753), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT105), .B(G137), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G39));
  NAND2_X1  g584(.A1(new_n763), .A2(new_n764), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n467), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n765), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n578), .A2(new_n597), .ZN(new_n778));
  AOI211_X1 g592(.A(new_n721), .B(new_n778), .C1(new_n525), .C2(new_n528), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n734), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  NOR2_X1   g595(.A1(G952), .A2(G953), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT115), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n715), .A2(new_n717), .A3(new_n529), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n423), .A3(new_n749), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n668), .A3(new_n667), .A4(new_n703), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT109), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(KEYINPUT109), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n703), .A2(KEYINPUT110), .A3(new_n734), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n691), .B2(new_n735), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n793), .A2(new_n423), .A3(new_n795), .A4(new_n749), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n725), .B2(new_n726), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n793), .A2(new_n795), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n681), .A2(new_n529), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n423), .A2(new_n798), .A3(new_n420), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n633), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n690), .A2(new_n754), .A3(new_n294), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n774), .B2(new_n776), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n734), .A3(new_n785), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n792), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT51), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n805), .B2(KEYINPUT111), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n805), .A3(new_n792), .A4(new_n802), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n422), .B(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n785), .A2(new_n730), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT113), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n798), .A2(new_n423), .A3(new_n684), .A4(new_n799), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n796), .A2(new_n601), .A3(new_n529), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT48), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n809), .A2(new_n812), .A3(new_n813), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n817), .A2(new_n819), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n808), .B2(new_n806), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n813), .A4(new_n812), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n745), .B1(new_n739), .B2(new_n741), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n634), .A2(new_n641), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n300), .A3(new_n615), .A4(new_n430), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n607), .A2(new_n608), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n657), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n700), .A2(new_n708), .A3(new_n719), .A4(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n464), .A2(new_n660), .A3(new_n420), .A4(new_n685), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n736), .B1(new_n834), .B2(new_n727), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n598), .A2(new_n599), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT82), .B1(new_n601), .B2(new_n529), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n838), .A2(new_n469), .B1(new_n696), .B2(new_n635), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n828), .A2(new_n833), .A3(new_n835), .A4(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n731), .A2(new_n665), .A3(new_n686), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n608), .A2(new_n618), .A3(new_n669), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n656), .A3(new_n685), .A4(new_n681), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(KEYINPUT108), .A3(KEYINPUT52), .A4(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n778), .A2(new_n655), .A3(new_n664), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n845), .A2(new_n663), .B1(new_n727), .B2(new_n730), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT52), .A3(new_n686), .A4(new_n843), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n731), .A2(new_n665), .A3(new_n686), .A4(new_n843), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT108), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n844), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n848), .B(KEYINPUT52), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n833), .A2(new_n828), .A3(new_n835), .A4(new_n839), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n855), .A2(new_n854), .A3(new_n856), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n856), .A2(KEYINPUT107), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n603), .A2(new_n697), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n708), .A2(new_n719), .A3(new_n832), .A4(new_n700), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT107), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n828), .A4(new_n835), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n861), .A2(new_n866), .A3(new_n844), .A4(new_n852), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n860), .B1(new_n867), .B2(new_n854), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n859), .B1(new_n868), .B2(new_n858), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n783), .B1(new_n827), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n690), .A2(new_n294), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT49), .Z(new_n872));
  AND4_X1   g686(.A1(new_n420), .A2(new_n872), .A3(new_n633), .A4(new_n667), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n300), .A3(new_n467), .A4(new_n799), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n874), .ZN(G75));
  AOI21_X1  g689(.A(new_n188), .B1(new_n853), .B2(new_n857), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT56), .B1(new_n876), .B2(G210), .ZN(new_n877));
  INV_X1    g691(.A(new_n345), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n315), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT55), .Z(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n877), .A2(new_n881), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n421), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  XNOR2_X1  g699(.A(new_n295), .B(KEYINPUT116), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT57), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n853), .A2(new_n858), .A3(new_n857), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n858), .B1(new_n853), .B2(new_n857), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT117), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n892), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n689), .B(KEYINPUT118), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n876), .A2(G469), .A3(new_n759), .A4(new_n758), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n884), .B1(new_n895), .B2(new_n896), .ZN(G54));
  NAND2_X1  g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n876), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n413), .A2(new_n401), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n884), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n876), .A2(new_n902), .A3(new_n899), .A4(new_n900), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n904), .A2(KEYINPUT120), .A3(new_n905), .A4(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(G60));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT59), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n628), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n888), .B2(new_n889), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n917), .A2(KEYINPUT121), .A3(new_n905), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n628), .B1(new_n869), .B2(new_n914), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT121), .B1(new_n917), .B2(new_n905), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(G63));
  AND2_X1   g735(.A1(new_n853), .A2(new_n857), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n652), .A2(new_n653), .ZN(new_n923));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT60), .ZN(new_n925));
  OR3_X1    g739(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n526), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n922), .B2(new_n925), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n905), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n926), .A2(KEYINPUT61), .A3(new_n905), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(G66));
  OAI21_X1  g747(.A(G953), .B1(new_n425), .B2(new_n310), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(KEYINPUT122), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n864), .B2(G953), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(KEYINPUT122), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n878), .B1(G898), .B2(new_n421), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n937), .B(new_n938), .Z(G69));
  XOR2_X1   g753(.A(new_n550), .B(KEYINPUT123), .Z(new_n940));
  AND2_X1   g754(.A1(new_n407), .A2(new_n408), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n940), .B(new_n941), .Z(new_n942));
  AND2_X1   g756(.A1(new_n829), .A2(new_n734), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n838), .A2(new_n675), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n768), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n768), .A2(new_n944), .A3(KEYINPUT125), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n780), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n682), .ZN(new_n953));
  NAND2_X1  g767(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n731), .A2(new_n665), .A3(new_n686), .A4(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n841), .A2(new_n950), .A3(new_n951), .A4(new_n682), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n949), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n942), .B1(new_n959), .B2(new_n421), .ZN(new_n960));
  NAND2_X1  g774(.A1(G900), .A2(G953), .ZN(new_n961));
  INV_X1    g775(.A(new_n942), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n618), .A2(new_n669), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n765), .A2(new_n598), .A3(new_n753), .A4(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n828), .A2(new_n964), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n768), .A2(new_n965), .A3(new_n780), .A4(new_n841), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n962), .B1(new_n966), .B2(new_n421), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n960), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n191), .B2(new_n661), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n591), .A2(new_n557), .A3(new_n544), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n677), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n868), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n966), .B2(new_n864), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n905), .B1(new_n977), .B2(new_n974), .ZN(new_n978));
  INV_X1    g792(.A(new_n864), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n949), .A2(new_n958), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT126), .B1(new_n980), .B2(new_n973), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n947), .A2(new_n780), .A3(new_n948), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(new_n864), .A3(new_n956), .A4(new_n957), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(new_n984), .A3(new_n972), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n981), .A2(new_n985), .A3(new_n678), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n981), .A2(new_n985), .A3(new_n988), .A4(new_n678), .ZN(new_n989));
  AOI211_X1 g803(.A(new_n976), .B(new_n978), .C1(new_n987), .C2(new_n989), .ZN(G57));
endmodule


