

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  INV_X2 U325 ( .A(n557), .ZN(n562) );
  XOR2_X1 U326 ( .A(n309), .B(n308), .Z(n549) );
  XOR2_X1 U327 ( .A(n545), .B(KEYINPUT28), .Z(n516) );
  XOR2_X1 U328 ( .A(KEYINPUT101), .B(KEYINPUT34), .Z(n455) );
  XOR2_X1 U329 ( .A(G15GAT), .B(G127GAT), .Z(n399) );
  XNOR2_X1 U330 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n293) );
  XNOR2_X1 U331 ( .A(n293), .B(G120GAT), .ZN(n342) );
  XOR2_X1 U332 ( .A(n399), .B(n342), .Z(n295) );
  XNOR2_X1 U333 ( .A(G43GAT), .B(G134GAT), .ZN(n294) );
  XNOR2_X1 U334 ( .A(n295), .B(n294), .ZN(n301) );
  XOR2_X1 U335 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n297) );
  XNOR2_X1 U336 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n361) );
  XOR2_X1 U338 ( .A(n361), .B(G176GAT), .Z(n299) );
  NAND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U341 ( .A(n301), .B(n300), .Z(n309) );
  XOR2_X1 U342 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n303) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G190GAT), .ZN(n302) );
  XNOR2_X1 U344 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U345 ( .A(KEYINPUT87), .B(G71GAT), .Z(n305) );
  XNOR2_X1 U346 ( .A(KEYINPUT86), .B(G183GAT), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U348 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U349 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n311) );
  NAND2_X1 U350 ( .A1(G228GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U351 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U352 ( .A(n312), .B(KEYINPUT90), .Z(n317) );
  XOR2_X1 U353 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n314) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(G218GAT), .ZN(n313) );
  XNOR2_X1 U355 ( .A(n314), .B(n313), .ZN(n354) );
  XNOR2_X1 U356 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n315) );
  XNOR2_X1 U357 ( .A(n315), .B(KEYINPUT2), .ZN(n341) );
  XNOR2_X1 U358 ( .A(n354), .B(n341), .ZN(n316) );
  XNOR2_X1 U359 ( .A(n317), .B(n316), .ZN(n324) );
  XOR2_X1 U360 ( .A(G204GAT), .B(G211GAT), .Z(n319) );
  XNOR2_X1 U361 ( .A(KEYINPUT92), .B(KEYINPUT23), .ZN(n318) );
  XNOR2_X1 U362 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U363 ( .A(n320), .B(KEYINPUT89), .Z(n322) );
  XOR2_X1 U364 ( .A(G22GAT), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U365 ( .A(n398), .B(KEYINPUT93), .ZN(n321) );
  XNOR2_X1 U366 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U367 ( .A(n324), .B(n323), .Z(n328) );
  XNOR2_X1 U368 ( .A(G50GAT), .B(KEYINPUT81), .ZN(n325) );
  XNOR2_X1 U369 ( .A(n325), .B(G162GAT), .ZN(n393) );
  XNOR2_X1 U370 ( .A(G106GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U371 ( .A(n326), .B(G148GAT), .ZN(n423) );
  XNOR2_X1 U372 ( .A(n393), .B(n423), .ZN(n327) );
  XNOR2_X1 U373 ( .A(n328), .B(n327), .ZN(n545) );
  XOR2_X1 U374 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n330) );
  XNOR2_X1 U375 ( .A(G1GAT), .B(G57GAT), .ZN(n329) );
  XNOR2_X1 U376 ( .A(n330), .B(n329), .ZN(n337) );
  XOR2_X1 U377 ( .A(G155GAT), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U378 ( .A(G127GAT), .B(G162GAT), .ZN(n331) );
  XNOR2_X1 U379 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U380 ( .A(G134GAT), .B(KEYINPUT82), .Z(n377) );
  XOR2_X1 U381 ( .A(n333), .B(n377), .Z(n335) );
  XNOR2_X1 U382 ( .A(G29GAT), .B(G85GAT), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U384 ( .A(n337), .B(n336), .ZN(n346) );
  XOR2_X1 U385 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n339) );
  NAND2_X1 U386 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U387 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U388 ( .A(n340), .B(KEYINPUT5), .Z(n344) );
  XNOR2_X1 U389 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U390 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U391 ( .A(n346), .B(n345), .ZN(n543) );
  XOR2_X1 U392 ( .A(G36GAT), .B(G190GAT), .Z(n384) );
  INV_X1 U393 ( .A(G64GAT), .ZN(n347) );
  NAND2_X1 U394 ( .A1(G92GAT), .A2(n347), .ZN(n350) );
  INV_X1 U395 ( .A(G92GAT), .ZN(n348) );
  NAND2_X1 U396 ( .A1(n348), .A2(G64GAT), .ZN(n349) );
  NAND2_X1 U397 ( .A1(n350), .A2(n349), .ZN(n352) );
  XNOR2_X1 U398 ( .A(G204GAT), .B(KEYINPUT77), .ZN(n351) );
  XNOR2_X1 U399 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U400 ( .A(G176GAT), .B(n353), .ZN(n431) );
  XOR2_X1 U401 ( .A(n354), .B(n431), .Z(n356) );
  XOR2_X1 U402 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n355) );
  XNOR2_X1 U403 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U404 ( .A(n384), .B(n357), .Z(n359) );
  NAND2_X1 U405 ( .A1(G226GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U406 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U407 ( .A(n361), .B(n360), .ZN(n363) );
  XOR2_X1 U408 ( .A(G8GAT), .B(G183GAT), .Z(n362) );
  XOR2_X1 U409 ( .A(G211GAT), .B(n362), .Z(n402) );
  XNOR2_X1 U410 ( .A(n363), .B(n402), .ZN(n496) );
  INV_X1 U411 ( .A(n496), .ZN(n540) );
  XOR2_X1 U412 ( .A(KEYINPUT27), .B(n540), .Z(n370) );
  NAND2_X1 U413 ( .A1(n543), .A2(n370), .ZN(n514) );
  NOR2_X1 U414 ( .A1(n516), .A2(n514), .ZN(n364) );
  XNOR2_X1 U415 ( .A(n364), .B(KEYINPUT97), .ZN(n365) );
  NOR2_X1 U416 ( .A1(n549), .A2(n365), .ZN(n376) );
  NAND2_X1 U417 ( .A1(n496), .A2(n549), .ZN(n366) );
  NAND2_X1 U418 ( .A1(n545), .A2(n366), .ZN(n367) );
  XOR2_X1 U419 ( .A(KEYINPUT25), .B(n367), .Z(n372) );
  NOR2_X1 U420 ( .A1(n545), .A2(n549), .ZN(n369) );
  XNOR2_X1 U421 ( .A(KEYINPUT26), .B(KEYINPUT98), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n566) );
  NAND2_X1 U423 ( .A1(n566), .A2(n370), .ZN(n371) );
  NAND2_X1 U424 ( .A1(n372), .A2(n371), .ZN(n373) );
  XNOR2_X1 U425 ( .A(KEYINPUT99), .B(n373), .ZN(n374) );
  NOR2_X1 U426 ( .A1(n543), .A2(n374), .ZN(n375) );
  NOR2_X1 U427 ( .A1(n376), .A2(n375), .ZN(n463) );
  XOR2_X1 U428 ( .A(KEYINPUT10), .B(n377), .Z(n379) );
  XOR2_X1 U429 ( .A(G99GAT), .B(G85GAT), .Z(n424) );
  XNOR2_X1 U430 ( .A(G218GAT), .B(n424), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U432 ( .A(KEYINPUT65), .B(G92GAT), .Z(n381) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U435 ( .A(n383), .B(n382), .Z(n386) );
  XNOR2_X1 U436 ( .A(G106GAT), .B(n384), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U438 ( .A(KEYINPUT66), .B(KEYINPUT83), .Z(n388) );
  XNOR2_X1 U439 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U441 ( .A(n390), .B(n389), .Z(n395) );
  XOR2_X1 U442 ( .A(G29GAT), .B(G43GAT), .Z(n392) );
  XNOR2_X1 U443 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n447) );
  XNOR2_X1 U445 ( .A(n447), .B(n393), .ZN(n394) );
  XNOR2_X1 U446 ( .A(n395), .B(n394), .ZN(n561) );
  XOR2_X1 U447 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n397) );
  XNOR2_X1 U448 ( .A(KEYINPUT84), .B(KEYINPUT14), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n413) );
  XOR2_X1 U450 ( .A(G64GAT), .B(n398), .Z(n401) );
  XNOR2_X1 U451 ( .A(n399), .B(G78GAT), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n406) );
  XOR2_X1 U453 ( .A(n402), .B(KEYINPUT85), .Z(n404) );
  NAND2_X1 U454 ( .A1(G231GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U455 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U456 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U457 ( .A(KEYINPUT72), .B(G1GAT), .Z(n446) );
  XOR2_X1 U458 ( .A(KEYINPUT75), .B(G57GAT), .Z(n408) );
  XNOR2_X1 U459 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n407) );
  XNOR2_X1 U460 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U461 ( .A(KEYINPUT74), .B(n409), .Z(n428) );
  XNOR2_X1 U462 ( .A(n446), .B(n428), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U464 ( .A(n413), .B(n412), .ZN(n577) );
  INV_X1 U465 ( .A(n577), .ZN(n507) );
  NOR2_X1 U466 ( .A1(n561), .A2(n507), .ZN(n414) );
  XOR2_X1 U467 ( .A(KEYINPUT16), .B(n414), .Z(n415) );
  NOR2_X1 U468 ( .A1(n463), .A2(n415), .ZN(n416) );
  XOR2_X1 U469 ( .A(KEYINPUT100), .B(n416), .Z(n481) );
  XOR2_X1 U470 ( .A(KEYINPUT79), .B(KEYINPUT32), .Z(n418) );
  XNOR2_X1 U471 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U473 ( .A(KEYINPUT78), .B(KEYINPUT33), .Z(n420) );
  XNOR2_X1 U474 ( .A(KEYINPUT80), .B(KEYINPUT76), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U476 ( .A(n422), .B(n421), .Z(n430) );
  XOR2_X1 U477 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U478 ( .A1(G230GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U482 ( .A(n432), .B(n431), .ZN(n572) );
  XOR2_X1 U483 ( .A(G141GAT), .B(G197GAT), .Z(n434) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(G22GAT), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U486 ( .A(KEYINPUT73), .B(G8GAT), .Z(n436) );
  XNOR2_X1 U487 ( .A(G113GAT), .B(G15GAT), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U489 ( .A(n438), .B(n437), .Z(n443) );
  XOR2_X1 U490 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n440) );
  NAND2_X1 U491 ( .A1(G229GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U493 ( .A(KEYINPUT67), .B(n441), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n453) );
  XOR2_X1 U495 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n445) );
  XNOR2_X1 U496 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n451) );
  XOR2_X1 U498 ( .A(n446), .B(G50GAT), .Z(n449) );
  XNOR2_X1 U499 ( .A(n447), .B(G36GAT), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U501 ( .A(n451), .B(n450), .Z(n452) );
  XNOR2_X1 U502 ( .A(n453), .B(n452), .ZN(n568) );
  NAND2_X1 U503 ( .A1(n572), .A2(n568), .ZN(n466) );
  NOR2_X1 U504 ( .A1(n481), .A2(n466), .ZN(n460) );
  NAND2_X1 U505 ( .A1(n460), .A2(n543), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U507 ( .A(G1GAT), .B(n456), .ZN(G1324GAT) );
  NAND2_X1 U508 ( .A1(n460), .A2(n496), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U510 ( .A(G15GAT), .B(KEYINPUT35), .Z(n459) );
  NAND2_X1 U511 ( .A1(n460), .A2(n549), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(G1326GAT) );
  NAND2_X1 U513 ( .A1(n460), .A2(n516), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n461), .B(KEYINPUT102), .ZN(n462) );
  XNOR2_X1 U515 ( .A(G22GAT), .B(n462), .ZN(G1327GAT) );
  XOR2_X1 U516 ( .A(KEYINPUT36), .B(n561), .Z(n581) );
  NOR2_X1 U517 ( .A1(n581), .A2(n463), .ZN(n464) );
  NAND2_X1 U518 ( .A1(n507), .A2(n464), .ZN(n465) );
  XOR2_X1 U519 ( .A(KEYINPUT37), .B(n465), .Z(n494) );
  NOR2_X1 U520 ( .A1(n466), .A2(n494), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n467), .B(KEYINPUT38), .ZN(n477) );
  NAND2_X1 U522 ( .A1(n477), .A2(n543), .ZN(n470) );
  XNOR2_X1 U523 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n468) );
  XNOR2_X1 U524 ( .A(n468), .B(KEYINPUT103), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n470), .B(n469), .ZN(G1328GAT) );
  XOR2_X1 U526 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n472) );
  NAND2_X1 U527 ( .A1(n496), .A2(n477), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U529 ( .A(G36GAT), .B(n473), .ZN(G1329GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n475) );
  NAND2_X1 U531 ( .A1(n477), .A2(n549), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U533 ( .A(G43GAT), .B(n476), .Z(G1330GAT) );
  XOR2_X1 U534 ( .A(G50GAT), .B(KEYINPUT107), .Z(n479) );
  NAND2_X1 U535 ( .A1(n516), .A2(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1331GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n483) );
  INV_X1 U538 ( .A(n568), .ZN(n527) );
  XNOR2_X1 U539 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n572), .B(n480), .ZN(n531) );
  XNOR2_X1 U541 ( .A(n531), .B(KEYINPUT108), .ZN(n554) );
  NAND2_X1 U542 ( .A1(n527), .A2(n554), .ZN(n493) );
  NOR2_X1 U543 ( .A1(n481), .A2(n493), .ZN(n490) );
  NAND2_X1 U544 ( .A1(n490), .A2(n543), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U546 ( .A(G57GAT), .B(n484), .ZN(G1332GAT) );
  NAND2_X1 U547 ( .A1(n490), .A2(n496), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n485), .B(KEYINPUT110), .ZN(n486) );
  XNOR2_X1 U549 ( .A(G64GAT), .B(n486), .ZN(G1333GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n488) );
  NAND2_X1 U551 ( .A1(n490), .A2(n549), .ZN(n487) );
  XNOR2_X1 U552 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U553 ( .A(G71GAT), .B(n489), .ZN(G1334GAT) );
  XOR2_X1 U554 ( .A(G78GAT), .B(KEYINPUT43), .Z(n492) );
  NAND2_X1 U555 ( .A1(n490), .A2(n516), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(G1335GAT) );
  NOR2_X1 U557 ( .A1(n494), .A2(n493), .ZN(n499) );
  NAND2_X1 U558 ( .A1(n543), .A2(n499), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G85GAT), .B(n495), .ZN(G1336GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n496), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U562 ( .A1(n549), .A2(n499), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U564 ( .A1(n499), .A2(n516), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(KEYINPUT44), .ZN(n501) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(n501), .ZN(G1339GAT) );
  NAND2_X1 U567 ( .A1(n531), .A2(n568), .ZN(n502) );
  XNOR2_X1 U568 ( .A(KEYINPUT46), .B(n502), .ZN(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT113), .B(n577), .ZN(n558) );
  NAND2_X1 U570 ( .A1(n503), .A2(n558), .ZN(n504) );
  NOR2_X1 U571 ( .A1(n561), .A2(n504), .ZN(n505) );
  XOR2_X1 U572 ( .A(KEYINPUT114), .B(n505), .Z(n506) );
  XNOR2_X1 U573 ( .A(n506), .B(KEYINPUT47), .ZN(n512) );
  NOR2_X1 U574 ( .A1(n581), .A2(n507), .ZN(n508) );
  XNOR2_X1 U575 ( .A(KEYINPUT45), .B(n508), .ZN(n509) );
  NAND2_X1 U576 ( .A1(n509), .A2(n572), .ZN(n510) );
  NOR2_X1 U577 ( .A1(n568), .A2(n510), .ZN(n511) );
  NOR2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(KEYINPUT48), .B(n513), .ZN(n539) );
  NOR2_X1 U580 ( .A1(n539), .A2(n514), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n526), .A2(n549), .ZN(n515) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n523), .A2(n568), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(n517), .ZN(G1340GAT) );
  XOR2_X1 U585 ( .A(G120GAT), .B(KEYINPUT49), .Z(n519) );
  NAND2_X1 U586 ( .A1(n523), .A2(n554), .ZN(n518) );
  XNOR2_X1 U587 ( .A(n519), .B(n518), .ZN(G1341GAT) );
  INV_X1 U588 ( .A(n523), .ZN(n520) );
  NOR2_X1 U589 ( .A1(n558), .A2(n520), .ZN(n521) );
  XOR2_X1 U590 ( .A(KEYINPUT50), .B(n521), .Z(n522) );
  XNOR2_X1 U591 ( .A(G127GAT), .B(n522), .ZN(G1342GAT) );
  XOR2_X1 U592 ( .A(G134GAT), .B(KEYINPUT51), .Z(n525) );
  NAND2_X1 U593 ( .A1(n523), .A2(n561), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n525), .B(n524), .ZN(G1343GAT) );
  NAND2_X1 U595 ( .A1(n566), .A2(n526), .ZN(n530) );
  NOR2_X1 U596 ( .A1(n527), .A2(n530), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(G1344GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n533) );
  INV_X1 U600 ( .A(n530), .ZN(n537) );
  NAND2_X1 U601 ( .A1(n537), .A2(n531), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U603 ( .A(G148GAT), .B(n534), .ZN(G1345GAT) );
  NAND2_X1 U604 ( .A1(n577), .A2(n537), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n535), .B(KEYINPUT116), .ZN(n536) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(n536), .ZN(G1346GAT) );
  NAND2_X1 U607 ( .A1(n537), .A2(n561), .ZN(n538) );
  XNOR2_X1 U608 ( .A(n538), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U609 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n547) );
  NOR2_X1 U610 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U611 ( .A(KEYINPUT54), .B(KEYINPUT117), .ZN(n541) );
  XNOR2_X1 U612 ( .A(n542), .B(n541), .ZN(n544) );
  NOR2_X1 U613 ( .A1(n544), .A2(n543), .ZN(n567) );
  NAND2_X1 U614 ( .A1(n567), .A2(n545), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n568), .A2(n562), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n552) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(n553), .Z(n556) );
  NAND2_X1 U623 ( .A1(n562), .A2(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(G190GAT), .B(n565), .Z(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n580) );
  INV_X1 U634 ( .A(n580), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n576), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n574) );
  OR2_X1 U639 ( .A1(n580), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT124), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(n584), .B(KEYINPUT126), .Z(n586) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1355GAT) );
endmodule

