//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT64), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT64), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(KEYINPUT65), .B(G125), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT64), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n478), .B(new_n479), .C1(new_n466), .C2(new_n467), .ZN(new_n480));
  INV_X1    g055(.A(G137), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n472), .A2(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n466), .A2(new_n467), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n463), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n484), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n477), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n484), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n480), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n473), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n500), .A2(new_n463), .A3(new_n501), .A4(G138), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n494), .B1(new_n496), .B2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT66), .B(G651), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT68), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n504), .B2(new_n511), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(G88), .A3(new_n506), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(G50), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n514), .A2(KEYINPUT67), .A3(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n506), .B(KEYINPUT69), .ZN(new_n527));
  INV_X1    g102(.A(G63), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n531), .B1(new_n514), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g108(.A(KEYINPUT70), .B(new_n513), .C1(new_n504), .C2(new_n511), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT71), .B(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n514), .A2(new_n506), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n530), .A2(new_n536), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n542), .B1(new_n529), .B2(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(KEYINPUT72), .A3(new_n536), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(G168));
  NAND2_X1  g124(.A1(new_n514), .A2(new_n532), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n550), .A2(G543), .A3(new_n534), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G64), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n527), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(new_n505), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n514), .A2(new_n506), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G90), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n552), .A2(new_n556), .A3(new_n558), .ZN(G171));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n527), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT73), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n564), .B(new_n560), .C1(new_n527), .C2(new_n561), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n505), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n551), .A2(G43), .B1(G81), .B2(new_n557), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(G860), .A3(new_n567), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  NAND3_X1  g148(.A1(new_n550), .A2(G543), .A3(new_n534), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n533), .A2(new_n577), .A3(G53), .A4(new_n534), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  OR3_X1    g156(.A1(new_n580), .A2(new_n581), .A3(new_n512), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n580), .B2(new_n512), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n582), .A2(new_n583), .B1(G91), .B2(new_n557), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n579), .A2(new_n584), .ZN(G299));
  NAND3_X1  g160(.A1(new_n552), .A2(new_n556), .A3(new_n558), .ZN(G301));
  NOR2_X1   g161(.A1(new_n544), .A2(new_n545), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT72), .B1(new_n547), .B2(new_n536), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(G286));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n506), .B(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n591), .B2(G74), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n557), .A2(G87), .ZN(new_n593));
  INV_X1    g168(.A(G49), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n574), .ZN(G288));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n506), .A2(G61), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n504), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n596), .A2(new_n540), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AND2_X1   g177(.A1(G48), .A2(G543), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n599), .A2(new_n600), .B1(new_n514), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(new_n551), .A2(G47), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n527), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n505), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n557), .A2(G85), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT77), .Z(new_n614));
  INV_X1    g189(.A(G54), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n574), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n616), .B2(new_n574), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n557), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n540), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n506), .A2(G66), .ZN(new_n623));
  INV_X1    g198(.A(G79), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(new_n531), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n619), .A2(new_n622), .B1(G651), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n614), .B1(G868), .B2(new_n627), .ZN(G284));
  OAI21_X1  g203(.A(new_n614), .B1(G868), .B2(new_n627), .ZN(G321));
  NOR2_X1   g204(.A1(G299), .A2(G868), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g206(.A(new_n630), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n627), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n566), .A2(new_n567), .ZN(new_n635));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n618), .A2(new_n626), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n638), .A2(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n637), .B1(new_n639), .B2(new_n636), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g216(.A1(G123), .A2(new_n485), .B1(new_n488), .B2(G135), .ZN(new_n642));
  OAI221_X1 g217(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(G2096), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n500), .A2(new_n474), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT12), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n646), .A2(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2451), .B(G2454), .Z(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n665), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(G401));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2100), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2096), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(KEYINPUT24), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G34), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT82), .B(G29), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n698), .B2(G34), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n699), .B1(new_n701), .B2(KEYINPUT93), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(KEYINPUT93), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT94), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  INV_X1    g280(.A(G160), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G2084), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT31), .B(G11), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n711), .B2(G28), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(G28), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n712), .B2(KEYINPUT96), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n710), .B1(new_n713), .B2(new_n715), .C1(new_n645), .C2(new_n700), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n705), .A2(G32), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT26), .Z(new_n719));
  INV_X1    g294(.A(new_n485), .ZN(new_n720));
  INV_X1    g295(.A(G129), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n474), .A2(G105), .ZN(new_n723));
  INV_X1    g298(.A(new_n488), .ZN(new_n724));
  INV_X1    g299(.A(G141), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n717), .B1(new_n727), .B2(new_n705), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT27), .B(G1996), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n709), .A2(new_n716), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n700), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G27), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G164), .B2(new_n732), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT97), .B(G2078), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n707), .B2(new_n708), .ZN(new_n738));
  INV_X1    g313(.A(G16), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G5), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G171), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n731), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n705), .A2(G33), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT25), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n500), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n463), .B1(new_n750), .B2(KEYINPUT91), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(KEYINPUT91), .B2(new_n750), .ZN(new_n752));
  INV_X1    g327(.A(G139), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n724), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n745), .B1(new_n757), .B2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G2072), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n744), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n762));
  NAND2_X1  g337(.A1(G286), .A2(G16), .ZN(new_n763));
  INV_X1    g338(.A(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(G16), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT95), .B(G1966), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n763), .B(new_n766), .C1(G16), .C2(new_n764), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n758), .A2(new_n759), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n761), .A2(new_n762), .A3(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(G16), .A2(G19), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n635), .B2(new_n739), .ZN(new_n775));
  INV_X1    g350(.A(G1341), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n700), .A2(G26), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  OAI221_X1 g355(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT88), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n488), .A2(G140), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT87), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n485), .A2(G128), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(G29), .ZN(new_n787));
  INV_X1    g362(.A(G2067), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n775), .A2(new_n776), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n732), .A2(G35), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n732), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT29), .B(G2090), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n777), .A2(new_n789), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n739), .A2(G20), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT23), .Z(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G299), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT100), .B(G1956), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n739), .A2(G4), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n627), .B2(new_n739), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1348), .Z(new_n803));
  AND3_X1   g378(.A1(new_n795), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n773), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n762), .B1(new_n761), .B2(new_n772), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n739), .A2(G23), .ZN(new_n808));
  INV_X1    g383(.A(G288), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n739), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT84), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT84), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT33), .B(G1976), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G6), .B(G305), .S(G16), .Z(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n811), .A2(new_n814), .A3(new_n812), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n739), .A2(G22), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G166), .B2(new_n739), .ZN(new_n822));
  INV_X1    g397(.A(G1971), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n816), .A2(new_n819), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(KEYINPUT34), .ZN(new_n826));
  MUX2_X1   g401(.A(G24), .B(G290), .S(G16), .Z(new_n827));
  INV_X1    g402(.A(G1986), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT86), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n732), .A2(G25), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n485), .A2(G119), .ZN(new_n832));
  OAI221_X1 g407(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n488), .A2(G131), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n831), .B1(new_n836), .B2(new_n732), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT83), .Z(new_n838));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G1991), .Z(new_n839));
  AOI21_X1  g414(.A(new_n830), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n829), .B(new_n840), .C1(new_n839), .C2(new_n838), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n826), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n825), .A2(KEYINPUT85), .A3(KEYINPUT34), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT85), .B1(new_n825), .B2(KEYINPUT34), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n842), .B(KEYINPUT36), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n807), .A2(new_n847), .A3(new_n848), .ZN(G311));
  NAND3_X1  g424(.A1(new_n807), .A2(new_n847), .A3(new_n848), .ZN(G150));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n527), .B2(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n853), .A2(new_n505), .B1(G93), .B2(new_n557), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n551), .A2(G55), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT102), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n627), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n856), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n566), .A2(new_n567), .A3(new_n855), .A4(new_n854), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n861), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT101), .Z(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n865), .B2(new_n866), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n859), .B1(new_n868), .B2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n786), .B(G164), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(new_n726), .B2(new_n722), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n496), .A2(new_n502), .ZN(new_n874));
  INV_X1    g449(.A(new_n494), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n786), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n727), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n757), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n835), .B(KEYINPUT103), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(new_n648), .Z(new_n883));
  AOI22_X1  g458(.A1(G130), .A2(new_n485), .B1(new_n488), .B2(G142), .ZN(new_n884));
  OAI221_X1 g459(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n883), .B(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n873), .B(new_n878), .C1(new_n749), .C2(new_n754), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n881), .B2(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n881), .A2(new_n887), .A3(KEYINPUT104), .A4(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n645), .B(G160), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(G162), .Z(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n881), .A2(new_n888), .ZN(new_n899));
  INV_X1    g474(.A(new_n887), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(new_n896), .A3(new_n889), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT40), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n896), .B1(new_n892), .B2(new_n893), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n907), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n906), .A2(new_n909), .ZN(G395));
  OR2_X1    g485(.A1(new_n864), .A2(new_n639), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n864), .A2(new_n639), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n638), .A2(G299), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n618), .A2(new_n579), .A3(new_n584), .A4(new_n626), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n914), .A2(KEYINPUT105), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT105), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n915), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n914), .A2(KEYINPUT41), .A3(new_n915), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n913), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n927), .A2(KEYINPUT107), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n930));
  AND2_X1   g505(.A1(G290), .A2(G288), .ZN(new_n931));
  NOR2_X1   g506(.A1(G290), .A2(G288), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(G305), .B(G303), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n809), .A2(new_n606), .A3(new_n610), .A4(new_n611), .ZN(new_n936));
  NAND2_X1  g511(.A1(G290), .A2(G288), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(KEYINPUT106), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n934), .A2(KEYINPUT106), .A3(new_n937), .A4(new_n936), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(KEYINPUT107), .B2(new_n927), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n919), .B(new_n925), .C1(KEYINPUT107), .C2(new_n927), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n929), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n929), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n856), .A2(new_n636), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(G295));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n948), .ZN(G331));
  NAND3_X1  g525(.A1(new_n546), .A2(new_n548), .A3(G301), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G301), .B1(new_n546), .B2(new_n548), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n864), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(G168), .A2(G171), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(new_n862), .A3(new_n951), .A4(new_n863), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n954), .B(new_n956), .C1(new_n917), .C2(new_n916), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n956), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n957), .A2(KEYINPUT108), .B1(new_n924), .B2(new_n958), .ZN(new_n959));
  OR3_X1    g534(.A1(new_n958), .A2(new_n918), .A3(KEYINPUT108), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n941), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n954), .A2(new_n956), .A3(new_n914), .A4(new_n915), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n954), .A2(new_n956), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n922), .A2(new_n923), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n941), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n903), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n961), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n966), .A2(new_n903), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n942), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT43), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n961), .A2(KEYINPUT43), .A3(new_n967), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n962), .B1(new_n969), .B2(new_n971), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(G397));
  XNOR2_X1  g553(.A(new_n786), .B(new_n788), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n979), .A2(new_n727), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT109), .B(G1384), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(G164), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n478), .A2(new_n479), .ZN(new_n984));
  INV_X1    g559(.A(G125), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n498), .B2(new_n499), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n464), .B1(new_n986), .B2(KEYINPUT65), .ZN(new_n987));
  INV_X1    g562(.A(new_n471), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n482), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(G40), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n983), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n994));
  INV_X1    g569(.A(G1996), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n993), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n980), .A2(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT47), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n993), .A2(G1986), .A3(G290), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT48), .Z(new_n1001));
  XNOR2_X1  g576(.A(new_n727), .B(G1996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n979), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n835), .B(new_n839), .Z(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1001), .B1(new_n1005), .B2(new_n993), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n836), .A2(new_n839), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n1003), .A2(new_n1007), .B1(G2067), .B2(new_n786), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n992), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n999), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n876), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n991), .B1(new_n1012), .B2(KEYINPUT50), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n876), .A2(new_n1015), .A3(new_n1011), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1013), .A2(new_n1014), .A3(new_n708), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1018));
  INV_X1    g593(.A(G40), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n472), .A2(new_n1019), .A3(new_n482), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1016), .A2(new_n1018), .A3(new_n708), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT119), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(G164), .B2(G1384), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1020), .B(new_n1024), .C1(new_n1012), .C2(new_n981), .ZN(new_n1025));
  INV_X1    g600(.A(G1966), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1017), .A2(new_n1022), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT113), .B(G8), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(G286), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT126), .B(KEYINPUT51), .Z(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(G8), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n546), .A2(new_n548), .A3(new_n1029), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1030), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1018), .A2(new_n1020), .A3(KEYINPUT118), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1016), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT118), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1040), .A2(G2090), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G164), .A2(new_n982), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n991), .B1(new_n1043), .B2(KEYINPUT45), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n981), .B1(G164), .B2(G1384), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1971), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1029), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n521), .A2(new_n522), .ZN(new_n1050));
  OAI211_X1 g625(.A(G8), .B(new_n1049), .C1(new_n1050), .C2(new_n516), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n517), .B2(new_n523), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1047), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1961), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n1059));
  INV_X1    g634(.A(new_n982), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1020), .A3(new_n1045), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1062), .A2(G2078), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1058), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1059), .A2(G2078), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1025), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(G301), .B(KEYINPUT54), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT127), .B(G2078), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n991), .A2(new_n1059), .A3(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1061), .A2(new_n983), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1066), .A2(new_n1067), .B1(new_n1071), .B2(new_n1064), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n602), .B2(new_n604), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n514), .A2(new_n603), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n597), .A2(new_n598), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n505), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1079), .B2(KEYINPUT76), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1080), .A2(new_n601), .A3(G1981), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1074), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n602), .A2(new_n1075), .A3(new_n604), .ZN(new_n1083));
  OAI21_X1  g658(.A(G1981), .B1(new_n1080), .B2(new_n601), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1083), .B(new_n1084), .C1(new_n1073), .C2(KEYINPUT49), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G164), .A2(G1384), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1020), .A2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1087), .A2(new_n1029), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(G288), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1088), .B(new_n1091), .C1(new_n1090), .C2(G288), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1087), .B(new_n1029), .C1(G288), .C2(new_n1090), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT52), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G2090), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1016), .A2(new_n1018), .A3(new_n1096), .A4(new_n1020), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1055), .B(G8), .C1(new_n1046), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT112), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1062), .A2(new_n823), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1052), .B1(new_n1101), .B2(new_n1097), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n1055), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1095), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1038), .A2(new_n1057), .A3(new_n1072), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1087), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1020), .A2(new_n1086), .A3(KEYINPUT122), .ZN(new_n1109));
  AOI21_X1  g684(.A(G2067), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1348), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n627), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND3_X1  g690(.A1(new_n1108), .A2(new_n1109), .A3(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1061), .A2(new_n1020), .A3(new_n1045), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n995), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n635), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g696(.A(KEYINPUT59), .B(new_n635), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1114), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1112), .A2(new_n638), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n627), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1113), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(G299), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n579), .A2(new_n584), .A3(new_n1130), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1956), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT56), .B(G2072), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1117), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1134), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1129), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT124), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1141), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(KEYINPUT125), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1134), .A2(new_n1136), .A3(new_n1146), .A4(new_n1138), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT61), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1149), .B(new_n1129), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1127), .A2(new_n1143), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1125), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1141), .B1(new_n1152), .B2(new_n1139), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1106), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1089), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1028), .A2(G168), .A3(new_n1029), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1155), .A2(new_n1057), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1099), .A2(KEYINPUT112), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1103), .B1(new_n1102), .B2(new_n1055), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1156), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(G8), .B1(new_n1046), .B2(new_n1098), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1159), .B1(new_n1165), .B2(new_n1056), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1157), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1161), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1105), .A2(KEYINPUT120), .A3(new_n1157), .A4(new_n1166), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1160), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1155), .A2(new_n1095), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1089), .A2(new_n1090), .A3(new_n809), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1081), .B(KEYINPUT116), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1174), .A2(KEYINPUT117), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1088), .B(KEYINPUT115), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1174), .B2(KEYINPUT117), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1171), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1170), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1155), .A2(new_n1057), .A3(new_n1156), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1066), .A2(G171), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1184), .B(new_n1030), .C1(new_n1034), .C2(new_n1037), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1180), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1154), .A2(new_n1179), .A3(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(G290), .B(new_n828), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n993), .B1(new_n1005), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1010), .B1(new_n1187), .B2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g765(.A1(new_n975), .A2(new_n976), .ZN(new_n1192));
  OR3_X1    g766(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1193));
  NOR2_X1   g767(.A1(G229), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n1194), .B1(new_n907), .B2(new_n904), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1192), .A2(new_n1195), .ZN(G308));
  OAI221_X1 g770(.A(new_n1194), .B1(new_n907), .B2(new_n904), .C1(new_n975), .C2(new_n976), .ZN(G225));
endmodule


