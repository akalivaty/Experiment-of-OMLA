//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT97), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n203), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n211), .A2(KEYINPUT17), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT17), .B1(new_n211), .B2(new_n212), .ZN(new_n214));
  INV_X1    g013(.A(G8gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(G1gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n217), .B2(KEYINPUT98), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n218), .B(new_n221), .ZN(new_n222));
  OR3_X1    g021(.A1(new_n213), .A2(new_n214), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n211), .A2(new_n212), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n222), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT18), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n225), .B(new_n222), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n224), .B(KEYINPUT13), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G113gat), .B(G141gat), .Z(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT96), .B(KEYINPUT11), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G169gat), .B(G197gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n229), .A2(new_n232), .A3(new_n233), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  INV_X1    g046(.A(G113gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(G120gat), .ZN(new_n249));
  INV_X1    g048(.A(G120gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(G113gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n246), .B(new_n247), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  INV_X1    g052(.A(G127gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(G134gat), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G127gat), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n253), .A2(KEYINPUT1), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT2), .ZN(new_n261));
  INV_X1    g060(.A(G148gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(G141gat), .ZN(new_n263));
  INV_X1    g062(.A(G141gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G148gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G155gat), .ZN(new_n267));
  INV_X1    g066(.A(G162gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n260), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n269), .B2(new_n260), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT80), .ZN(new_n275));
  XNOR2_X1  g074(.A(G155gat), .B(G162gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT79), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n271), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT80), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n266), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n263), .A2(KEYINPUT81), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n262), .B2(G141gat), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n281), .B(new_n283), .C1(new_n264), .C2(G148gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n260), .B1(new_n269), .B2(KEYINPUT2), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n275), .A2(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n259), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n285), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT80), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n279), .B1(new_n278), .B2(new_n266), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n289), .B(new_n259), .C1(new_n290), .C2(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT4), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n286), .A2(new_n297), .A3(new_n259), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n302));
  INV_X1    g101(.A(new_n259), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n295), .ZN(new_n305));
  INV_X1    g104(.A(new_n300), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n288), .B2(new_n293), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n286), .A2(new_n310), .A3(new_n297), .A4(new_n259), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT84), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .A4(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G1gat), .B(G29gat), .Z(new_n315));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT85), .B(KEYINPUT6), .ZN(new_n321));
  INV_X1    g120(.A(new_n319), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n308), .A2(new_n322), .A3(new_n313), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n308), .B2(new_n313), .ZN(new_n325));
  INV_X1    g124(.A(new_n321), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n325), .A2(KEYINPUT86), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT86), .B1(new_n325), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n331));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT24), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G183gat), .B(G190gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(G169gat), .ZN(new_n339));
  INV_X1    g138(.A(G176gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT65), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G176gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT23), .ZN(new_n346));
  INV_X1    g145(.A(G169gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n340), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n331), .B1(new_n337), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n331), .B1(new_n352), .B2(KEYINPUT23), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G183gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G183gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n333), .B1(new_n359), .B2(KEYINPUT24), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT66), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n357), .C1(new_n355), .C2(KEYINPUT27), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT27), .ZN(new_n367));
  AOI21_X1  g166(.A(G190gat), .B1(new_n367), .B2(G183gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n355), .A2(KEYINPUT27), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n368), .A2(KEYINPUT66), .A3(new_n365), .A4(new_n369), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT26), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n348), .A2(new_n373), .A3(new_n345), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n352), .A2(KEYINPUT26), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n375), .A2(new_n332), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n371), .A2(new_n372), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n362), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G226gat), .ZN(new_n379));
  INV_X1    g178(.A(G233gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT72), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT72), .ZN(new_n383));
  INV_X1    g182(.A(new_n381), .ZN(new_n384));
  INV_X1    g183(.A(new_n372), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n364), .A2(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n373), .B1(G169gat), .B2(G176gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n345), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n375), .B(new_n332), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n351), .B2(new_n361), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n383), .B(new_n384), .C1(new_n391), .C2(KEYINPUT29), .ZN(new_n392));
  NAND2_X1  g191(.A1(G211gat), .A2(G218gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT22), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G197gat), .B(G204gat), .ZN(new_n396));
  INV_X1    g195(.A(G211gat), .ZN(new_n397));
  INV_X1    g196(.A(G218gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT71), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n393), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n399), .B2(new_n393), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n395), .B(new_n396), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n396), .A2(new_n395), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n362), .A2(new_n377), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n381), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n382), .A2(new_n392), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n382), .A2(new_n392), .A3(new_n411), .A4(KEYINPUT73), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n384), .B1(new_n391), .B2(KEYINPUT29), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n410), .A2(new_n381), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n408), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n330), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n419), .B1(new_n414), .B2(new_n415), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT78), .A3(new_n424), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n329), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n420), .A4(new_n424), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT76), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n428), .A2(KEYINPUT76), .A3(KEYINPUT30), .A4(new_n424), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT74), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT74), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n439), .A3(new_n425), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT75), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n416), .B2(new_n420), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT74), .B(new_n419), .C1(new_n414), .C2(new_n415), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(KEYINPUT75), .A3(new_n425), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n436), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n431), .B1(new_n447), .B2(KEYINPUT77), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n434), .A2(new_n435), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT75), .B1(new_n445), .B2(new_n425), .ZN(new_n450));
  NOR4_X1   g249(.A1(new_n443), .A2(new_n444), .A3(new_n441), .A4(new_n424), .ZN(new_n451));
  OAI211_X1 g250(.A(KEYINPUT77), .B(new_n449), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT65), .B(G176gat), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n455), .A2(new_n339), .B1(new_n348), .B2(new_n346), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT25), .B1(new_n456), .B2(new_n360), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n349), .A2(new_n353), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n337), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n377), .B(new_n259), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n362), .A2(new_n462), .A3(new_n377), .A4(new_n259), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n359), .A2(KEYINPUT24), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(new_n334), .A3(new_n344), .A4(new_n349), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n465), .A2(new_n331), .B1(new_n354), .B2(new_n360), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n303), .B1(new_n466), .B2(new_n390), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n461), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G227gat), .A2(G233gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT64), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n454), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G43gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT68), .ZN(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n471), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT33), .B1(new_n468), .B2(new_n470), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n479));
  NOR4_X1   g278(.A1(new_n471), .A2(new_n478), .A3(new_n479), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n468), .A2(new_n470), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n481), .B2(KEYINPUT32), .ZN(new_n482));
  INV_X1    g281(.A(new_n478), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT69), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n477), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT34), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n487), .B(new_n477), .C1(new_n480), .C2(new_n484), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n468), .A2(new_n470), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT29), .B1(new_n404), .B2(new_n407), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n292), .B1(KEYINPUT3), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n287), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n409), .ZN(new_n500));
  INV_X1    g299(.A(G228gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(new_n380), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n292), .B(KEYINPUT88), .C1(KEYINPUT3), .C2(new_n493), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n496), .A2(new_n500), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G22gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n404), .A2(new_n407), .A3(KEYINPUT87), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n506), .B(new_n498), .C1(KEYINPUT87), .C2(new_n407), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n286), .B1(new_n507), .B2(new_n287), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n408), .B1(new_n497), .B2(new_n498), .ZN(new_n509));
  OAI22_X1  g308(.A1(new_n508), .A2(new_n509), .B1(new_n501), .B2(new_n380), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n505), .B1(new_n504), .B2(new_n510), .ZN(new_n512));
  OAI21_X1  g311(.A(G78gat), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n504), .A2(new_n510), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(G78gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT31), .B(G50gat), .ZN(new_n519));
  INV_X1    g318(.A(G106gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n513), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n513), .B2(new_n518), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n486), .A2(new_n490), .A3(new_n488), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n492), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n448), .A2(new_n453), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT35), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT95), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n486), .A2(new_n490), .A3(new_n488), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n490), .B1(new_n486), .B2(new_n488), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n492), .A2(KEYINPUT95), .A3(new_n525), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n449), .B(new_n430), .C1(new_n450), .C2(new_n451), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT89), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n442), .A2(new_n446), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n449), .A4(new_n430), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n513), .A2(new_n518), .A3(new_n521), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n513), .A2(new_n518), .ZN(new_n541));
  INV_X1    g340(.A(new_n521), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND4_X1   g342(.A1(new_n528), .A2(new_n329), .A3(new_n540), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  OAI22_X1  g344(.A1(new_n527), .A2(new_n528), .B1(new_n534), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n540), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n448), .B2(new_n453), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n551), .B(new_n552), .C1(new_n530), .C2(new_n531), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n492), .A2(new_n549), .A3(new_n550), .A4(new_n525), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT39), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n312), .A2(new_n294), .A3(new_n311), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT90), .A3(new_n306), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT90), .B1(new_n557), .B2(new_n306), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n305), .A2(new_n306), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(new_n556), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n565), .A3(new_n322), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT40), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(KEYINPUT91), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(KEYINPUT91), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n566), .A2(KEYINPUT91), .A3(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n320), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n536), .B2(new_n539), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n417), .A2(new_n408), .A3(new_n418), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT92), .Z(new_n576));
  NAND3_X1  g375(.A1(new_n382), .A2(new_n392), .A3(new_n418), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n409), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT93), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n578), .A2(KEYINPUT93), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT37), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n583));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n424), .B1(new_n428), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n328), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n325), .A2(KEYINPUT86), .A3(new_n326), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n426), .A2(new_n429), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n586), .A2(new_n589), .A3(new_n590), .A4(new_n324), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n583), .B1(new_n592), .B2(new_n585), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n524), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n548), .B(new_n555), .C1(new_n574), .C2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n245), .B1(new_n546), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G57gat), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT99), .B1(new_n597), .B2(G64gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n599));
  INV_X1    g398(.A(G64gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(G57gat), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n598), .B(new_n601), .C1(G57gat), .C2(new_n600), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT100), .ZN(new_n603));
  NAND2_X1  g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(G71gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n516), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT9), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G57gat), .B(G64gat), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n604), .B(new_n606), .C1(new_n610), .C2(new_n607), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(new_n254), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n222), .B1(new_n612), .B2(KEYINPUT21), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT101), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G155gat), .ZN(new_n621));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n618), .A2(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(G230gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n380), .ZN(new_n629));
  XNOR2_X1  g428(.A(G99gat), .B(G106gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n612), .B1(KEYINPUT103), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G85gat), .A2(G92gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT7), .ZN(new_n633));
  NAND2_X1  g432(.A1(G99gat), .A2(G106gat), .ZN(new_n634));
  INV_X1    g433(.A(G85gat), .ZN(new_n635));
  INV_X1    g434(.A(G92gat), .ZN(new_n636));
  AOI22_X1  g435(.A1(KEYINPUT8), .A2(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n630), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n631), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n631), .A2(new_n640), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n639), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n629), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n629), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n641), .B2(new_n643), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G120gat), .B(G148gat), .Z(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n225), .A2(new_n639), .B1(KEYINPUT41), .B2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n213), .A2(new_n214), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n639), .B(KEYINPUT102), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G190gat), .B(G218gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n656), .A2(KEYINPUT41), .ZN(new_n663));
  XNOR2_X1  g462(.A(G134gat), .B(G162gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n662), .B(new_n665), .Z(new_n666));
  NOR3_X1   g465(.A1(new_n627), .A2(new_n655), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n596), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n596), .A2(KEYINPUT104), .A3(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n329), .B(KEYINPUT105), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g474(.A1(new_n536), .A2(new_n539), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT16), .B(G8gat), .Z(new_n677));
  AND3_X1   g476(.A1(new_n672), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n215), .B1(new_n672), .B2(new_n676), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT42), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(KEYINPUT42), .B2(new_n678), .ZN(G1325gat));
  INV_X1    g480(.A(new_n672), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n682), .A2(G15gat), .A3(new_n534), .ZN(new_n683));
  OAI21_X1  g482(.A(G15gat), .B1(new_n682), .B2(new_n555), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n672), .A2(new_n547), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(new_n666), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n626), .A2(new_n655), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n596), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n673), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n691), .A2(G29gat), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT45), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n655), .B(KEYINPUT106), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(new_n245), .A3(new_n626), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n546), .A2(new_n595), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n666), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n666), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n546), .B2(new_n595), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n699), .A2(KEYINPUT44), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n697), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n707), .A2(new_n673), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n694), .B1(new_n708), .B2(new_n206), .ZN(G1328gat));
  INV_X1    g508(.A(new_n676), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n691), .A2(G36gat), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n707), .A2(new_n676), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(new_n207), .ZN(G1329gat));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n555), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n707), .B2(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n691), .A2(G43gat), .A3(new_n534), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT109), .B(KEYINPUT47), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  INV_X1    g519(.A(new_n701), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n548), .A2(new_n555), .ZN(new_n722));
  INV_X1    g521(.A(new_n573), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n594), .B1(new_n676), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n545), .ZN(new_n726));
  INV_X1    g525(.A(new_n534), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n530), .A2(new_n547), .A3(new_n531), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT77), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n728), .A2(new_n452), .A3(new_n731), .A4(new_n431), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n726), .A2(new_n727), .B1(new_n732), .B2(KEYINPUT35), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n703), .B(new_n721), .C1(new_n725), .C2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n689), .B1(new_n546), .B2(new_n595), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n716), .B(new_n696), .C1(new_n737), .C2(new_n705), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n718), .B1(new_n738), .B2(G43gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n720), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n719), .A2(new_n741), .ZN(G1330gat));
  INV_X1    g541(.A(G50gat), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n707), .B2(new_n547), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n691), .A2(G50gat), .A3(new_n524), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n746));
  OR3_X1    g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n744), .B2(new_n745), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  INV_X1    g548(.A(new_n695), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n626), .A2(new_n245), .A3(new_n689), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n750), .B(new_n751), .C1(new_n546), .C2(new_n595), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n673), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n676), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT49), .B(G64gat), .Z(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(G1333gat));
  AOI21_X1  g557(.A(new_n605), .B1(new_n752), .B2(new_n716), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n534), .A2(G71gat), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n752), .A2(new_n547), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n626), .A2(new_n244), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n699), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n698), .A2(new_n666), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n673), .A2(new_n635), .A3(new_n655), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT112), .Z(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n655), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n768), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n704), .B2(new_n706), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n673), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n780), .B2(new_n635), .ZN(G1336gat));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n750), .A2(new_n710), .A3(G92gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n772), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n779), .A2(new_n676), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n782), .B(new_n784), .C1(new_n785), .C2(new_n636), .ZN(new_n786));
  INV_X1    g585(.A(new_n784), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n636), .B1(new_n779), .B2(new_n676), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT52), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(G1337gat));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n716), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G99gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n534), .A2(G99gat), .A3(new_n776), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT113), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n772), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1338gat));
  OAI211_X1 g595(.A(new_n547), .B(new_n777), .C1(new_n737), .C2(new_n705), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G106gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n695), .A2(new_n520), .A3(new_n547), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT114), .Z(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT115), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n772), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805));
  AOI211_X1 g604(.A(new_n689), .B(new_n768), .C1(new_n546), .C2(new_n595), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n771), .B(new_n800), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n769), .A2(new_n810), .A3(new_n771), .A4(new_n800), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n805), .A2(new_n798), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT53), .B1(new_n797), .B2(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n805), .B1(new_n815), .B2(new_n812), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n804), .B1(new_n814), .B2(new_n816), .ZN(G1339gat));
  NAND2_X1  g616(.A1(new_n644), .A2(new_n645), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n647), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n644), .A2(new_n629), .A3(new_n645), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n652), .B1(new_n646), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(new_n823), .A3(KEYINPUT55), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n654), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n224), .B1(new_n223), .B2(new_n226), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n230), .A2(new_n231), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n239), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n831), .A2(KEYINPUT118), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(KEYINPUT118), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n243), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n828), .A2(new_n689), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n826), .A2(new_n244), .A3(new_n654), .A4(new_n827), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n655), .A2(new_n243), .A3(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n666), .B1(new_n839), .B2(KEYINPUT119), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n837), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n836), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI22_X1  g642(.A1(new_n843), .A2(new_n626), .B1(new_n655), .B2(new_n751), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n692), .A2(new_n676), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n728), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n248), .A3(new_n244), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n844), .A2(new_n524), .A3(new_n727), .A4(new_n845), .ZN(new_n849));
  OAI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n245), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT120), .ZN(G1340gat));
  NOR3_X1   g651(.A1(new_n849), .A2(new_n250), .A3(new_n750), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n847), .A2(new_n655), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n250), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n847), .A2(new_n254), .A3(new_n626), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n849), .B2(new_n627), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT121), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n847), .A2(new_n256), .A3(new_n666), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n849), .B2(new_n689), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n839), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT122), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n689), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n836), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n626), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n751), .A2(new_n655), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n547), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n844), .A2(new_n875), .A3(new_n547), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n716), .A2(new_n676), .A3(new_n692), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n874), .A2(new_n244), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n865), .B1(new_n878), .B2(G141gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n716), .A2(new_n524), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n244), .A2(new_n264), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT123), .Z(new_n882));
  AND4_X1   g681(.A1(new_n844), .A2(new_n845), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n878), .B2(G141gat), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n879), .A2(new_n884), .A3(KEYINPUT58), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886));
  AOI221_X4 g685(.A(new_n883), .B1(new_n865), .B2(new_n886), .C1(new_n878), .C2(G141gat), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n885), .A2(new_n887), .ZN(G1344gat));
  AND2_X1   g687(.A1(new_n846), .A2(new_n880), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n262), .A3(new_n655), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n776), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(KEYINPUT59), .A3(new_n262), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n873), .A2(new_n875), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n844), .A2(KEYINPUT57), .A3(new_n547), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n655), .B(new_n877), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n894), .B1(new_n898), .B2(G148gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n890), .B1(new_n893), .B2(new_n899), .ZN(G1345gat));
  OAI21_X1  g699(.A(G155gat), .B1(new_n891), .B2(new_n627), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n889), .A2(new_n267), .A3(new_n626), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n889), .B2(new_n666), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n891), .A2(new_n268), .A3(new_n689), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n692), .A2(new_n676), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n526), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n844), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n244), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n844), .A2(new_n524), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n534), .A3(new_n907), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n245), .A2(new_n347), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n909), .B2(new_n655), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n750), .A2(new_n455), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n912), .B2(new_n916), .ZN(G1349gat));
  AOI21_X1  g716(.A(new_n355), .B1(new_n912), .B2(new_n626), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n367), .A2(G183gat), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n909), .A2(new_n919), .A3(new_n369), .A4(new_n626), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n918), .A2(new_n921), .A3(KEYINPUT60), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT60), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1350gat));
  AOI21_X1  g723(.A(new_n357), .B1(new_n912), .B2(new_n666), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n909), .A2(new_n357), .A3(new_n666), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1351gat));
  NOR2_X1   g728(.A1(new_n716), .A2(new_n907), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n895), .B2(new_n897), .ZN(new_n931));
  INV_X1    g730(.A(G197gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n931), .A2(new_n932), .A3(new_n245), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n844), .A2(new_n547), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n244), .A3(new_n930), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n932), .B2(new_n935), .ZN(G1352gat));
  INV_X1    g735(.A(G204gat), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n695), .B(new_n930), .C1(new_n895), .C2(new_n897), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(KEYINPUT126), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(KEYINPUT126), .B2(new_n938), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n934), .A2(new_n930), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n941), .A2(G204gat), .A3(new_n776), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(G1353gat));
  AND4_X1   g743(.A1(new_n397), .A2(new_n934), .A3(new_n626), .A4(new_n930), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n626), .B(new_n930), .C1(new_n895), .C2(new_n897), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G211gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT63), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n948), .A2(new_n951), .A3(G211gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(new_n950), .A3(new_n952), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n931), .B2(new_n689), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n666), .A2(new_n398), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n941), .B2(new_n955), .ZN(G1355gat));
endmodule


