//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n583, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n607, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n642, new_n643, new_n644,
    new_n645, new_n648, new_n650, new_n651, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n468), .A2(G137), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT67), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(new_n471), .A3(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n481), .A2(new_n483), .A3(new_n470), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n479), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  OR2_X1    g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n486), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n477), .B1(new_n487), .B2(new_n488), .ZN(G160));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n465), .A2(new_n467), .ZN(new_n491));
  INV_X1    g066(.A(G112), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n484), .A2(new_n468), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n495), .A2(new_n496), .B1(G124), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n481), .A2(new_n483), .A3(new_n464), .A4(new_n470), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G136), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G162));
  AND2_X1   g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n481), .A2(new_n483), .A3(new_n470), .A4(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n506), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n465), .A2(new_n467), .A3(G138), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT4), .B1(new_n484), .B2(new_n511), .ZN(new_n512));
  OR3_X1    g087(.A1(new_n511), .A2(new_n473), .A3(KEYINPUT4), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n509), .A2(new_n510), .B1(new_n512), .B2(new_n513), .ZN(G164));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI21_X1  g101(.A(G543), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n520), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  AND3_X1   g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(G76), .A2(G543), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n534), .A2(new_n536), .B1(new_n538), .B2(G651), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n537), .A2(new_n539), .B1(new_n525), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g116(.A1(G63), .A2(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n517), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(new_n527), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT72), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G543), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT6), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(new_n519), .ZN(new_n549));
  NAND2_X1  g124(.A1(KEYINPUT6), .A2(G651), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G51), .B1(new_n517), .B2(new_n542), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n515), .A2(new_n516), .B1(new_n549), .B2(new_n550), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G89), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n534), .A2(new_n536), .ZN(new_n555));
  INV_X1    g130(.A(new_n532), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n552), .A2(new_n554), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n546), .A2(new_n561), .ZN(G168));
  INV_X1    g137(.A(G90), .ZN(new_n563));
  INV_X1    g138(.A(G52), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n525), .A2(new_n563), .B1(new_n527), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(G64), .B1(new_n522), .B2(new_n521), .ZN(new_n566));
  NAND2_X1  g141(.A1(G77), .A2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n519), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(G171));
  NAND2_X1  g144(.A1(G68), .A2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n522), .A2(new_n521), .ZN(new_n571));
  INV_X1    g146(.A(G56), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT73), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n576), .A3(G651), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n553), .A2(G81), .B1(new_n551), .B2(G43), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G860), .ZN(G153));
  NAND4_X1  g156(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g157(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n583));
  NAND2_X1  g158(.A1(G1), .A2(G3), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(G319), .A2(G483), .A3(G661), .A4(new_n585), .ZN(G188));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(G65), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(G65), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n517), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G78), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(KEYINPUT77), .A3(new_n591), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n594), .A2(G651), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G53), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT9), .B1(new_n527), .B2(new_n597), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n527), .A2(KEYINPUT9), .A3(new_n597), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n553), .A2(KEYINPUT75), .A3(G91), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n601));
  INV_X1    g176(.A(G91), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n525), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n598), .A2(new_n599), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n596), .A2(new_n604), .ZN(G299));
  INV_X1    g180(.A(G171), .ZN(G301));
  AND3_X1   g181(.A1(new_n546), .A2(KEYINPUT78), .A3(new_n561), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT78), .B1(new_n546), .B2(new_n561), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G286));
  INV_X1    g185(.A(G74), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n519), .B1(new_n571), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G49), .B2(new_n551), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n553), .A2(G87), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(G288));
  AOI22_X1  g190(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(new_n519), .ZN(new_n617));
  INV_X1    g192(.A(G86), .ZN(new_n618));
  INV_X1    g193(.A(G48), .ZN(new_n619));
  OAI22_X1  g194(.A1(new_n525), .A2(new_n618), .B1(new_n527), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(G305));
  AOI22_X1  g197(.A1(new_n553), .A2(G85), .B1(new_n551), .B2(G47), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT79), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n519), .B2(new_n625), .ZN(G290));
  NAND2_X1  g201(.A1(G301), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G79), .A2(G543), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT80), .ZN(new_n629));
  INV_X1    g204(.A(G66), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n571), .ZN(new_n631));
  AOI22_X1  g206(.A1(new_n631), .A2(G651), .B1(G54), .B2(new_n551), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n553), .A2(KEYINPUT10), .A3(G92), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT10), .ZN(new_n634));
  INV_X1    g209(.A(G92), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n525), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n627), .B1(new_n639), .B2(G868), .ZN(G284));
  OAI21_X1  g215(.A(new_n627), .B1(new_n639), .B2(G868), .ZN(G321));
  NAND2_X1  g216(.A1(G286), .A2(G868), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(KEYINPUT81), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(KEYINPUT81), .ZN(new_n644));
  INV_X1    g219(.A(G299), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n643), .B(new_n644), .C1(G868), .C2(new_n645), .ZN(G297));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(G868), .C2(new_n645), .ZN(G280));
  INV_X1    g222(.A(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n639), .B1(new_n648), .B2(G860), .ZN(G148));
  NAND2_X1  g224(.A1(new_n639), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G868), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(G868), .B2(new_n580), .ZN(G323));
  XNOR2_X1  g227(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g228(.A1(new_n474), .A2(new_n478), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  INV_X1    g232(.A(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n500), .A2(G135), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT83), .ZN(new_n661));
  OAI21_X1  g236(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n662));
  INV_X1    g237(.A(G111), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n491), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n497), .B2(G123), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G2096), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(G2096), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n659), .A2(new_n669), .A3(new_n670), .ZN(G156));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT84), .B(G2438), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2427), .B(G2430), .Z(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(KEYINPUT14), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2451), .B(G2454), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT16), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1341), .B(G1348), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n678), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2443), .B(G2446), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  AND3_X1   g261(.A1(new_n685), .A2(G14), .A3(new_n686), .ZN(G401));
  INV_X1    g262(.A(KEYINPUT18), .ZN(new_n688));
  XOR2_X1   g263(.A(G2084), .B(G2090), .Z(new_n689));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(KEYINPUT17), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(new_n658), .ZN(new_n695));
  XOR2_X1   g270(.A(G2072), .B(G2078), .Z(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n691), .B2(KEYINPUT18), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(new_n668), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(G227));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT19), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1956), .B(G2474), .Z(new_n703));
  XOR2_X1   g278(.A(G1961), .B(G1966), .Z(new_n704));
  AND2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n703), .A2(new_n704), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(new_n710), .B(new_n709), .S(new_n702), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1991), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1981), .B(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n719), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT87), .Z(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(G1971), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(G1971), .ZN(new_n724));
  NOR2_X1   g299(.A1(G6), .A2(G16), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n621), .B2(G16), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT32), .B(G1981), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n719), .A2(G23), .ZN(new_n729));
  INV_X1    g304(.A(G288), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n719), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT33), .B(G1976), .Z(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT86), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n731), .B(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n723), .A2(new_n724), .A3(new_n728), .A4(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT34), .ZN(new_n737));
  MUX2_X1   g312(.A(G24), .B(G290), .S(G16), .Z(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G1986), .Z(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G25), .ZN(new_n741));
  OAI221_X1 g316(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n742));
  INV_X1    g317(.A(new_n497), .ZN(new_n743));
  INV_X1    g318(.A(G119), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n500), .A2(G131), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(new_n740), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT35), .B(G1991), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT85), .Z(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n748), .B(new_n751), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n736), .A2(new_n737), .A3(new_n739), .A4(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n740), .A2(G35), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G162), .B2(new_n740), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT29), .Z(new_n758));
  INV_X1    g333(.A(G2090), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n740), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(KEYINPUT89), .B(new_n766), .C1(new_n468), .C2(G116), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n768));
  AOI21_X1  g343(.A(G116), .B1(new_n465), .B2(new_n467), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n765), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n767), .A2(new_n770), .B1(new_n497), .B2(G128), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n500), .A2(KEYINPUT88), .A3(G140), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT88), .ZN(new_n773));
  INV_X1    g348(.A(G140), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n499), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n764), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2067), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n760), .A2(new_n761), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n740), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n740), .ZN(new_n782));
  INV_X1    g357(.A(G2078), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n719), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G168), .B2(new_n719), .ZN(new_n786));
  INV_X1    g361(.A(G1966), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n740), .B1(new_n789), .B2(G34), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n789), .B2(G34), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G160), .B2(G29), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n784), .B(new_n788), .C1(G2084), .C2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(G28), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n740), .B1(new_n794), .B2(G28), .ZN(new_n796));
  AND2_X1   g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  NOR2_X1   g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  OAI22_X1  g373(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n719), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n719), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n799), .B1(new_n801), .B2(G1961), .ZN(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT26), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n805), .A2(new_n806), .B1(G105), .B2(new_n478), .ZN(new_n807));
  INV_X1    g382(.A(G129), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n743), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n500), .A2(G141), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n740), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n740), .B2(G32), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT27), .B(G1996), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n802), .B1(G1961), .B2(new_n801), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n639), .A2(new_n719), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G4), .B2(new_n719), .ZN(new_n818));
  INV_X1    g393(.A(G1348), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n818), .A2(new_n819), .B1(G29), .B2(new_n667), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n819), .B2(new_n818), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n719), .A2(G20), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT23), .Z(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G299), .B2(G16), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT93), .B(G1956), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G2084), .B2(new_n792), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n830));
  NAND2_X1  g405(.A1(G103), .A2(G2104), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n491), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n500), .A2(G139), .ZN(new_n834));
  NAND2_X1  g409(.A1(G115), .A2(G2104), .ZN(new_n835));
  INV_X1    g410(.A(G127), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n473), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n491), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n833), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(KEYINPUT91), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(KEYINPUT91), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n740), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n740), .B2(G33), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT92), .B(G2072), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(G16), .A2(G19), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n580), .B2(G16), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G1341), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n814), .B2(new_n815), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n822), .A2(new_n828), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  NOR4_X1   g427(.A1(new_n755), .A2(new_n780), .A3(new_n793), .A4(new_n852), .ZN(G311));
  OR4_X1    g428(.A1(new_n755), .A2(new_n780), .A3(new_n793), .A4(new_n852), .ZN(G150));
  AOI22_X1  g429(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n519), .ZN(new_n856));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  INV_X1    g432(.A(G55), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n525), .A2(new_n857), .B1(new_n527), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT95), .B(KEYINPUT37), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n639), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT38), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n856), .A2(new_n859), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n579), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n866), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT94), .Z(new_n872));
  OAI21_X1  g447(.A(new_n861), .B1(new_n869), .B2(new_n870), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n864), .B1(new_n872), .B2(new_n873), .ZN(G145));
  INV_X1    g449(.A(new_n656), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n839), .A2(KEYINPUT98), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n508), .B1(new_n513), .B2(new_n512), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n777), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n513), .A2(new_n512), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n771), .B(new_n776), .C1(new_n880), .C2(new_n508), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n879), .A2(new_n811), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n811), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n812), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT91), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n839), .A2(new_n887), .A3(KEYINPUT98), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n843), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n879), .A2(new_n811), .A3(new_n881), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n500), .A2(G142), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n468), .A2(G118), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n497), .A2(KEYINPUT99), .A3(G130), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT99), .B1(new_n497), .B2(G130), .ZN(new_n897));
  OAI221_X1 g472(.A(new_n893), .B1(new_n894), .B2(new_n895), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n747), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n884), .A2(new_n892), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n899), .B1(new_n884), .B2(new_n892), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n875), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n899), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n882), .A2(new_n883), .A3(new_n889), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n876), .B1(new_n886), .B2(new_n891), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n884), .A2(new_n892), .A3(new_n899), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n656), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n667), .A2(G162), .ZN(new_n912));
  INV_X1    g487(.A(G160), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n502), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n910), .A3(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n909), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n902), .A2(new_n921), .A3(new_n908), .ZN(new_n925));
  AND4_X1   g500(.A1(KEYINPUT100), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(G37), .B1(new_n909), .B2(new_n922), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT100), .B1(new_n927), .B2(new_n925), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(G395));
  XNOR2_X1  g506(.A(new_n579), .B(new_n860), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(new_n650), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  AND4_X1   g509(.A1(new_n596), .A2(new_n604), .A3(new_n637), .A4(new_n632), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n596), .A2(new_n604), .B1(new_n637), .B2(new_n632), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n639), .A2(new_n596), .A3(new_n604), .ZN(new_n938));
  NAND2_X1  g513(.A1(G299), .A2(new_n638), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT41), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n935), .A2(new_n936), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(new_n933), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT42), .Z(new_n945));
  XNOR2_X1  g520(.A(G290), .B(G305), .ZN(new_n946));
  XNOR2_X1  g521(.A(G303), .B(G288), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(KEYINPUT102), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n945), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(G868), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G868), .B2(new_n860), .ZN(G295));
  OAI21_X1  g527(.A(new_n951), .B1(G868), .B2(new_n860), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  INV_X1    g529(.A(new_n941), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT103), .B1(G168), .B2(G301), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n957));
  AOI211_X1 g532(.A(new_n957), .B(G171), .C1(new_n546), .C2(new_n561), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT78), .ZN(new_n960));
  NAND2_X1  g535(.A1(G168), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n546), .A2(KEYINPUT78), .A3(new_n561), .ZN(new_n962));
  AOI21_X1  g537(.A(G301), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n959), .A2(new_n963), .A3(new_n932), .ZN(new_n964));
  AOI22_X1  g539(.A1(G89), .A2(new_n553), .B1(new_n557), .B2(new_n558), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n560), .B1(new_n965), .B2(new_n552), .ZN(new_n966));
  AND4_X1   g541(.A1(new_n560), .A2(new_n552), .A3(new_n554), .A4(new_n559), .ZN(new_n967));
  OAI21_X1  g542(.A(G301), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n957), .ZN(new_n969));
  NAND3_X1  g544(.A1(G168), .A2(KEYINPUT103), .A3(G301), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(G171), .B1(new_n607), .B2(new_n608), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n868), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n955), .B1(new_n964), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n932), .B1(new_n959), .B2(new_n963), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n972), .B(new_n868), .C1(new_n956), .C2(new_n958), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(new_n943), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(KEYINPUT106), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n948), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n978), .B(new_n979), .C1(KEYINPUT106), .C2(new_n974), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n948), .A2(new_n974), .A3(new_n977), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n924), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n954), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n975), .A2(new_n943), .A3(new_n976), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n941), .B1(new_n975), .B2(new_n976), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n974), .A2(KEYINPUT104), .A3(new_n977), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n979), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n924), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT105), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(KEYINPUT105), .A3(new_n924), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n981), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n983), .B1(new_n994), .B2(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n981), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT105), .B1(new_n989), .B2(new_n924), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT107), .B1(new_n1001), .B2(new_n954), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n1003));
  AOI211_X1 g578(.A(new_n1003), .B(KEYINPUT44), .C1(new_n998), .C2(new_n1000), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n995), .B1(new_n1002), .B2(new_n1004), .ZN(G397));
  NAND2_X1  g580(.A1(G160), .A2(G40), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n878), .A2(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n811), .B(G1996), .ZN(new_n1012));
  INV_X1    g587(.A(G2067), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n777), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT109), .Z(new_n1017));
  XNOR2_X1  g592(.A(new_n747), .B(new_n751), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(G290), .B(G1986), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1011), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  AND2_X1   g598(.A1(G160), .A2(G40), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G164), .A2(G1384), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1009), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1008), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n787), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1007), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1024), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1023), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT51), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1031), .A2(G168), .A3(new_n1036), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(G8), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(G8), .ZN(new_n1042));
  AOI21_X1  g617(.A(G168), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1041), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT62), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1024), .A2(new_n1027), .A3(new_n783), .A4(new_n1029), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT53), .A3(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(G160), .B(G40), .C1(new_n1008), .C2(new_n1028), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n783), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  INV_X1    g631(.A(G1961), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1024), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1055), .A2(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1971), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1007), .A2(new_n1034), .ZN(new_n1063));
  OR3_X1    g638(.A1(new_n1006), .A2(KEYINPUT116), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT116), .B1(new_n1006), .B2(new_n1063), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1025), .A2(new_n1034), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(G2090), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G303), .A2(G8), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G288), .A2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT111), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1075), .A2(new_n1078), .A3(new_n1023), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n730), .A2(G1976), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1079), .B(new_n1080), .C1(KEYINPUT52), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1024), .A2(new_n1007), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1078), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n1080), .A4(G8), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1083), .A2(new_n1084), .A3(G8), .A4(new_n1081), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1075), .A2(new_n1023), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(G1981), .B1(new_n617), .B2(KEYINPUT113), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(new_n621), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT49), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1082), .A2(new_n1088), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1024), .A2(new_n759), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1062), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(G8), .A3(new_n1072), .ZN(new_n1102));
  AND4_X1   g677(.A1(new_n1060), .A2(new_n1074), .A3(new_n1099), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1041), .B(new_n1104), .C1(new_n1039), .C2(new_n1044), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1046), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(new_n1076), .A3(new_n730), .ZN(new_n1108));
  OR2_X1    g683(.A1(G305), .A2(G1981), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1090), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1099), .B(KEYINPUT115), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1102), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1037), .A2(new_n609), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1074), .A2(new_n1099), .A3(new_n1102), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1037), .A2(KEYINPUT63), .A3(new_n609), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1072), .B1(new_n1101), .B2(G8), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1118), .A2(new_n1112), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1088), .A2(new_n1082), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1122), .A2(KEYINPUT115), .A3(new_n1107), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1106), .A2(new_n1113), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(new_n1107), .A3(new_n1102), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1072), .B1(new_n1068), .B2(G8), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1056), .B1(KEYINPUT124), .B2(new_n783), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1010), .B(new_n1131), .C1(KEYINPUT124), .C2(new_n783), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1132), .A2(new_n1052), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1059), .A2(G301), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1060), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1051), .A2(G301), .A3(new_n1059), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1059), .A2(new_n1133), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1136), .B(KEYINPUT54), .C1(new_n1137), .C2(G301), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1045), .A2(new_n1129), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1956), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1067), .A2(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1142));
  NAND3_X1  g717(.A1(G299), .A2(KEYINPUT118), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(G299), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT118), .B1(G299), .B2(new_n1142), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT56), .B(G2072), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1054), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1141), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1147), .B1(new_n1141), .B2(new_n1149), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT120), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT61), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1058), .A2(new_n819), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1075), .A2(new_n1013), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OR3_X1    g732(.A1(new_n1157), .A2(KEYINPUT60), .A3(new_n638), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1157), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(new_n639), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT60), .B1(new_n1157), .B2(new_n638), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(KEYINPUT119), .B(G1996), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1054), .A2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(KEYINPUT58), .B(G1341), .Z(new_n1165));
  NAND2_X1  g740(.A1(new_n1083), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n579), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT59), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1162), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n1170));
  OAI211_X1 g745(.A(KEYINPUT120), .B(new_n1170), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1154), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1159), .A2(new_n638), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1152), .B1(new_n1150), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1139), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1022), .B1(new_n1126), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1011), .B1(new_n1015), .B2(new_n811), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT125), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1006), .A2(new_n1010), .A3(G1996), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT46), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT47), .Z(new_n1182));
  AND3_X1   g757(.A1(new_n1017), .A2(new_n751), .A3(new_n747), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n777), .A2(G2067), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1011), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(G290), .A2(G1986), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1011), .A2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g762(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1188));
  XNOR2_X1  g763(.A(new_n1187), .B(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1017), .A2(new_n1019), .A3(new_n1189), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1182), .A2(new_n1185), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1176), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  AOI21_X1  g768(.A(new_n999), .B1(new_n994), .B2(KEYINPUT43), .ZN(new_n1195));
  OR3_X1    g769(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G229), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g771(.A(new_n1197), .B1(new_n926), .B2(new_n928), .ZN(new_n1198));
  OAI21_X1  g772(.A(new_n1194), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g773(.A(new_n1197), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n927), .A2(new_n925), .ZN(new_n1201));
  INV_X1    g775(.A(KEYINPUT100), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g777(.A1(new_n927), .A2(KEYINPUT100), .A3(new_n925), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n1200), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g779(.A1(new_n1205), .A2(new_n1001), .A3(KEYINPUT127), .ZN(new_n1206));
  AND2_X1   g780(.A1(new_n1199), .A2(new_n1206), .ZN(G308));
  NAND2_X1  g781(.A1(new_n1199), .A2(new_n1206), .ZN(G225));
endmodule


