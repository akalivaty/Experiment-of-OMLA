//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n467), .A2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n473), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n464), .A2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n485), .B2(G124), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(G162));
  NAND4_X1  g062(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n466), .ZN(new_n488));
  OR2_X1    g063(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(KEYINPUT71), .B(KEYINPUT4), .Z(new_n491));
  NOR2_X1   g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(KEYINPUT70), .B2(G114), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT70), .A2(G114), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g082(.A(new_n507), .B(KEYINPUT72), .Z(new_n508));
  AOI22_X1  g083(.A1(new_n504), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  AND2_X1   g090(.A1(G76), .A2(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(KEYINPUT7), .B1(new_n516), .B2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n504), .A2(G63), .ZN(new_n518));
  NAND3_X1  g093(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n506), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n510), .A2(new_n511), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n504), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI211_X1 g098(.A(new_n517), .B(new_n520), .C1(G89), .C2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(G543), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT74), .B(G51), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n501), .A2(new_n503), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n523), .A2(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n527), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n534), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT76), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(G43), .B2(new_n528), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT77), .B(G81), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n523), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT78), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT80), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G188));
  XNOR2_X1  g137(.A(new_n522), .B(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G91), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(KEYINPUT81), .A2(KEYINPUT9), .ZN(new_n566));
  OR3_X1    g141(.A1(new_n527), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n506), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n566), .B1(new_n527), .B2(new_n565), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n564), .A2(new_n567), .A3(new_n569), .A4(new_n570), .ZN(G299));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n506), .B1(new_n534), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n563), .B2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n528), .A2(G49), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n563), .A2(G86), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n504), .A2(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n506), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n523), .A2(G85), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n506), .B2(new_n585), .C1(new_n586), .C2(new_n527), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n563), .A2(G92), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n506), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n528), .A2(G54), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n588), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n588), .B1(new_n595), .B2(G868), .ZN(G321));
  AND2_X1   g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G299), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT83), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(KEYINPUT83), .B2(new_n598), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(KEYINPUT83), .B2(new_n598), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n595), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n595), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n478), .A2(G135), .ZN(new_n611));
  NOR2_X1   g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(new_n485), .B2(G123), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT84), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2096), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2430), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT15), .B(G2435), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT87), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT86), .B(G2451), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n630), .B(new_n636), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XNOR2_X1  g214(.A(G2084), .B(G2090), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT88), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT17), .ZN(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n642), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n643), .B2(new_n646), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT89), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n644), .A2(new_n641), .A3(new_n646), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT90), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n642), .A2(new_n643), .A3(new_n646), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2096), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n660), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n667), .A2(KEYINPUT92), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n663), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1986), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1991), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n674), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G25), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n485), .A2(G119), .ZN(new_n682));
  OR2_X1    g257(.A1(G95), .A2(G2105), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n683), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT93), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n478), .A2(G131), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n681), .B1(new_n688), .B2(new_n680), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT35), .B(G1991), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G1986), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n694), .A2(G24), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G290), .B2(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n692), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n694), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1971), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(G23), .ZN(new_n701));
  INV_X1    g276(.A(G288), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n694), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT33), .Z(new_n704));
  AOI21_X1  g279(.A(new_n700), .B1(new_n704), .B2(G1976), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n694), .A2(G6), .ZN(new_n706));
  INV_X1    g281(.A(G305), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n694), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n705), .B(new_n710), .C1(G1976), .C2(new_n704), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT94), .B(KEYINPUT34), .Z(new_n712));
  AOI21_X1  g287(.A(new_n697), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n696), .A2(new_n693), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n713), .B(new_n714), .C1(new_n712), .C2(new_n711), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT36), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n694), .A2(G4), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n595), .B2(new_n694), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G1348), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n694), .A2(G19), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n553), .B2(new_n694), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n718), .A2(G1348), .B1(G1341), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G1341), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n680), .A2(G26), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n485), .A2(G128), .ZN(new_n725));
  OR2_X1    g300(.A1(G104), .A2(G2105), .ZN(new_n726));
  INV_X1    g301(.A(G116), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n469), .B1(new_n727), .B2(G2105), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n478), .A2(G140), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n724), .B1(new_n731), .B2(new_n680), .ZN(new_n732));
  MUX2_X1   g307(.A(new_n724), .B(new_n732), .S(KEYINPUT28), .Z(new_n733));
  AOI211_X1 g308(.A(new_n719), .B(new_n723), .C1(G2067), .C2(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(G2067), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT23), .B1(new_n600), .B2(new_n694), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n694), .A2(G20), .ZN(new_n737));
  MUX2_X1   g312(.A(KEYINPUT23), .B(new_n736), .S(new_n737), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G1956), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(G1956), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n734), .A2(new_n735), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n694), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n694), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT24), .A2(G34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(new_n680), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G160), .B2(new_n680), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT103), .B(G28), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT30), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n749), .A2(G2084), .B1(G29), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G21), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G168), .B2(G16), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G1966), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n752), .B(new_n755), .C1(G29), .C2(new_n616), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT102), .B(KEYINPUT31), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G11), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT99), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n485), .A2(G129), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n478), .A2(G141), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT97), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NAND3_X1  g340(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n761), .A2(new_n763), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(new_n680), .ZN(new_n768));
  NOR2_X1   g343(.A1(G29), .A2(G32), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n768), .A2(KEYINPUT98), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(KEYINPUT98), .B2(new_n768), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n756), .B(new_n758), .C1(new_n760), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n680), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n680), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT104), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G2078), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n754), .A2(G1966), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT101), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n772), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n771), .A2(new_n760), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n749), .A2(G2084), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G29), .B2(G33), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n782), .A2(G29), .A3(G33), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT25), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n478), .A2(G139), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n786), .B(new_n787), .C1(new_n466), .C2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n783), .B(new_n784), .C1(new_n790), .C2(new_n680), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2072), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n780), .A2(new_n781), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT100), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AND4_X1   g371(.A1(new_n745), .A2(new_n779), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT105), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n741), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n680), .A2(G35), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n680), .ZN(new_n801));
  MUX2_X1   g376(.A(new_n800), .B(new_n801), .S(KEYINPUT106), .Z(new_n802));
  XOR2_X1   g377(.A(KEYINPUT29), .B(G2090), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n797), .A2(new_n798), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n716), .A2(new_n799), .A3(new_n804), .A4(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  AOI22_X1  g382(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT107), .Z(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(new_n506), .ZN(new_n810));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  INV_X1    g386(.A(G93), .ZN(new_n812));
  OAI22_X1  g387(.A1(new_n527), .A2(new_n811), .B1(new_n812), .B2(new_n522), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT37), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n595), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n553), .A2(new_n815), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n552), .A2(new_n814), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT39), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n819), .B(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n817), .B1(new_n824), .B2(G860), .ZN(G145));
  XNOR2_X1  g400(.A(new_n790), .B(new_n730), .ZN(new_n826));
  INV_X1    g401(.A(new_n498), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n464), .A2(new_n828), .A3(G138), .A4(new_n466), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n488), .A2(new_n489), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT108), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT108), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n619), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n826), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n478), .A2(G142), .ZN(new_n836));
  NOR2_X1   g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n838));
  INV_X1    g413(.A(G130), .ZN(new_n839));
  OAI221_X1 g414(.A(new_n836), .B1(new_n837), .B2(new_n838), .C1(new_n484), .C2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n767), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n835), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n687), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n616), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G162), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n835), .A2(new_n841), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n835), .A2(new_n841), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n688), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n843), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT109), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(G37), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n843), .A2(new_n848), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n851), .B(new_n852), .C1(new_n845), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g430(.A1(new_n815), .A2(G868), .ZN(new_n856));
  XNOR2_X1  g431(.A(G288), .B(G290), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G303), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n707), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT42), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n595), .A2(new_n600), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n593), .A2(new_n594), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G299), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(KEYINPUT41), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT41), .B1(new_n861), .B2(new_n863), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n607), .B(new_n822), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n861), .A2(new_n863), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(new_n868), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n860), .B1(new_n871), .B2(KEYINPUT110), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(KEYINPUT110), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n872), .B(new_n873), .Z(new_n874));
  AOI21_X1  g449(.A(new_n856), .B1(new_n874), .B2(G868), .ZN(G295));
  AOI21_X1  g450(.A(new_n856), .B1(new_n874), .B2(G868), .ZN(G331));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n877));
  INV_X1    g452(.A(new_n859), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n870), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n820), .A2(G286), .A3(new_n821), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G286), .B1(new_n820), .B2(new_n821), .ZN(new_n883));
  OAI21_X1  g458(.A(G301), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n822), .A2(G168), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(G171), .A3(new_n881), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n880), .A2(new_n864), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n870), .A3(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n878), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT111), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n884), .A2(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n867), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT111), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n878), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n893), .A2(new_n878), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n877), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n891), .A2(new_n895), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n898), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(KEYINPUT44), .A3(new_n899), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n907), .ZN(G397));
  INV_X1    g483(.A(G1384), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT45), .B1(new_n833), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(KEYINPUT112), .B(G40), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n467), .A2(new_n476), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n767), .B(G1996), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n730), .B(G2067), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n691), .B2(new_n688), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n687), .A2(new_n690), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(new_n693), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n913), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT114), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n490), .B2(new_n492), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT108), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n498), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n924), .B1(new_n928), .B2(G1384), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n833), .A2(KEYINPUT114), .A3(new_n909), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G8), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n676), .ZN(new_n935));
  INV_X1    g510(.A(G86), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n578), .B1(new_n522), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT116), .ZN(new_n938));
  OAI21_X1  g513(.A(G1981), .B1(new_n938), .B2(new_n581), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n935), .A2(KEYINPUT49), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT49), .B1(new_n935), .B2(new_n939), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n934), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n943));
  INV_X1    g518(.A(G1976), .ZN(new_n944));
  NAND2_X1  g519(.A1(G288), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n702), .A2(G1976), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n933), .A2(new_n943), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n933), .A2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(new_n943), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n942), .B1(new_n949), .B2(KEYINPUT115), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT119), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT50), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n928), .A2(new_n924), .A3(G1384), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT114), .B1(new_n833), .B2(new_n909), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n909), .B1(new_n493), .B2(new_n498), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(new_n956), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n963), .A3(new_n913), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n964), .A2(G2090), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n833), .A2(KEYINPUT45), .A3(new_n909), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n966), .A2(new_n968), .A3(new_n913), .ZN(new_n969));
  INV_X1    g544(.A(G1971), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n932), .B1(new_n965), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G303), .A2(G8), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n975), .B(KEYINPUT55), .Z(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n955), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n929), .A2(KEYINPUT50), .A3(new_n930), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n979), .B(new_n913), .C1(KEYINPUT50), .C2(new_n960), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n971), .B1(new_n980), .B2(G2090), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n981), .A2(G8), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n976), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n953), .A2(new_n954), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n978), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n974), .A2(new_n976), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT63), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n974), .B2(new_n976), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n986), .A2(new_n988), .A3(new_n952), .A4(new_n950), .ZN(new_n989));
  INV_X1    g564(.A(G2084), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n959), .A2(new_n990), .A3(new_n963), .A4(new_n913), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n929), .A2(new_n967), .A3(new_n930), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n923), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1966), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT120), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(G1966), .C1(new_n993), .C2(new_n994), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n992), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n1000), .A2(new_n932), .A3(G286), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n989), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1956), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n980), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(G299), .B(KEYINPUT57), .Z(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT56), .B(G2072), .Z(new_n1006));
  OR2_X1    g581(.A1(new_n969), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n595), .ZN(new_n1009));
  AOI211_X1 g584(.A(G2067), .B(new_n923), .C1(new_n929), .C2(new_n930), .ZN(new_n1010));
  INV_X1    g585(.A(G1348), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n964), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1013));
  OAI22_X1  g588(.A1(new_n1009), .A2(new_n1012), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT58), .B(G1341), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT121), .B(G1996), .Z(new_n1016));
  OAI22_X1  g591(.A1(new_n931), .A2(new_n1015), .B1(new_n969), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT122), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  OAI221_X1 g594(.A(new_n1019), .B1(new_n969), .B2(new_n1016), .C1(new_n931), .C2(new_n1015), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n553), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1008), .A2(KEYINPUT61), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT61), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT123), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1018), .A2(new_n1020), .A3(KEYINPUT59), .A4(new_n553), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n595), .B1(new_n1012), .B2(KEYINPUT60), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT60), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1030), .B(new_n1010), .C1(new_n964), .C2(new_n1011), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n862), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1014), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G286), .A2(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT124), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT51), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1036), .B(new_n1039), .C1(new_n1000), .C2(new_n932), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n995), .A2(new_n996), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n998), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n995), .A2(KEYINPUT120), .A3(new_n996), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n991), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(G8), .A3(G286), .ZN(new_n1045));
  OAI211_X1 g620(.A(G8), .B(new_n1038), .C1(new_n1044), .C2(G286), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n969), .A2(G2078), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n964), .A2(new_n744), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G301), .B(KEYINPUT54), .ZN(new_n1051));
  INV_X1    g626(.A(G40), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n910), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n966), .A2(G160), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1054), .A2(new_n1049), .A3(G2078), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(KEYINPUT61), .B2(new_n1008), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n995), .A2(new_n1049), .A3(G2078), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1050), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1060), .B2(new_n1051), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1047), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1002), .B1(new_n1035), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1047), .A2(KEYINPUT62), .ZN(new_n1064));
  AOI21_X1  g639(.A(G301), .B1(new_n1050), .B2(new_n1059), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1040), .A2(new_n1046), .A3(new_n1066), .A4(new_n1045), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n985), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1001), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT63), .B1(new_n989), .B2(new_n1070), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n953), .A2(new_n977), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n933), .B(KEYINPUT117), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n942), .A2(G1976), .A3(G288), .ZN(new_n1074));
  XOR2_X1   g649(.A(new_n935), .B(KEYINPUT118), .Z(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1071), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n922), .B1(new_n1069), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n914), .A2(G1996), .ZN(new_n1081));
  NAND2_X1  g656(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n914), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n916), .B2(new_n767), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1083), .B(new_n1085), .C1(KEYINPUT125), .C2(KEYINPUT46), .ZN(new_n1086));
  XOR2_X1   g661(.A(new_n1086), .B(KEYINPUT47), .Z(new_n1087));
  OAI21_X1  g662(.A(new_n1084), .B1(new_n918), .B2(new_n919), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n914), .A2(G1986), .A3(G290), .ZN(new_n1089));
  XOR2_X1   g664(.A(new_n1089), .B(KEYINPUT48), .Z(new_n1090));
  AND2_X1   g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n730), .A2(G2067), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n917), .B2(new_n919), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(new_n914), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1087), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT126), .B1(new_n1080), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(new_n1002), .C1(new_n1035), .C2(new_n1062), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1078), .B1(new_n1100), .B2(new_n985), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1098), .B(new_n1095), .C1(new_n1101), .C2(new_n922), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1097), .A2(new_n1102), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g678(.A1(G401), .A2(G227), .ZN(new_n1105));
  INV_X1    g679(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g680(.A1(G229), .A2(new_n462), .ZN(new_n1107));
  NAND2_X1  g681(.A1(new_n854), .A2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g682(.A(new_n1106), .B(new_n1108), .C1(new_n906), .C2(new_n899), .ZN(G308));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n906), .B2(new_n899), .ZN(new_n1110));
  NAND3_X1  g684(.A1(new_n1110), .A2(new_n854), .A3(new_n1107), .ZN(G225));
endmodule


