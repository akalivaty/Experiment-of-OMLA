

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G168), .A2(n673), .ZN(n677) );
  XNOR2_X2 U550 ( .A(n719), .B(KEYINPUT32), .ZN(n733) );
  XNOR2_X1 U551 ( .A(n709), .B(KEYINPUT29), .ZN(n710) );
  INV_X2 U552 ( .A(G2105), .ZN(n514) );
  NOR2_X1 U553 ( .A1(G651), .A2(n612), .ZN(n632) );
  XNOR2_X2 U554 ( .A(n520), .B(n519), .ZN(n592) );
  INV_X1 U555 ( .A(KEYINPUT91), .ZN(n709) );
  NOR2_X1 U556 ( .A1(G1966), .A2(n760), .ZN(n721) );
  XNOR2_X1 U557 ( .A(n711), .B(n710), .ZN(n726) );
  AND2_X2 U558 ( .A1(n514), .A2(G2104), .ZN(n882) );
  INV_X1 U559 ( .A(KEYINPUT23), .ZN(n515) );
  NOR2_X1 U560 ( .A1(n612), .A2(n528), .ZN(n631) );
  XNOR2_X1 U561 ( .A(n516), .B(n515), .ZN(n517) );
  NOR2_X2 U562 ( .A1(n524), .A2(n523), .ZN(G160) );
  NOR2_X2 U563 ( .A1(G2104), .A2(n514), .ZN(n878) );
  NAND2_X1 U564 ( .A1(n878), .A2(G125), .ZN(n518) );
  NAND2_X1 U565 ( .A1(G101), .A2(n882), .ZN(n516) );
  NAND2_X1 U566 ( .A1(n518), .A2(n517), .ZN(n524) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U568 ( .A1(G113), .A2(n879), .ZN(n522) );
  XNOR2_X1 U569 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n520) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  NAND2_X1 U571 ( .A1(G137), .A2(n592), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n523) );
  INV_X1 U573 ( .A(G651), .ZN(n528) );
  NOR2_X1 U574 ( .A1(G543), .A2(n528), .ZN(n525) );
  XOR2_X1 U575 ( .A(KEYINPUT1), .B(n525), .Z(n628) );
  NAND2_X1 U576 ( .A1(G64), .A2(n628), .ZN(n527) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n612) );
  NAND2_X1 U578 ( .A1(G52), .A2(n632), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n533) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n627) );
  NAND2_X1 U581 ( .A1(G90), .A2(n627), .ZN(n530) );
  NAND2_X1 U582 ( .A1(G77), .A2(n631), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U584 ( .A(KEYINPUT9), .B(n531), .Z(n532) );
  NOR2_X1 U585 ( .A1(n533), .A2(n532), .ZN(G171) );
  AND2_X1 U586 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U587 ( .A(G132), .ZN(G219) );
  INV_X1 U588 ( .A(G82), .ZN(G220) );
  INV_X1 U589 ( .A(G69), .ZN(G235) );
  INV_X1 U590 ( .A(G57), .ZN(G237) );
  NAND2_X1 U591 ( .A1(G89), .A2(n627), .ZN(n534) );
  XOR2_X1 U592 ( .A(KEYINPUT4), .B(n534), .Z(n535) );
  XNOR2_X1 U593 ( .A(n535), .B(KEYINPUT71), .ZN(n537) );
  NAND2_X1 U594 ( .A1(G76), .A2(n631), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n538), .B(KEYINPUT5), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G63), .A2(n628), .ZN(n540) );
  NAND2_X1 U598 ( .A1(G51), .A2(n632), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U600 ( .A(KEYINPUT6), .B(n541), .Z(n542) );
  NAND2_X1 U601 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U602 ( .A(n544), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U604 ( .A1(G138), .A2(n592), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G102), .A2(n882), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G126), .A2(n878), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G114), .A2(n879), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U610 ( .A1(n550), .A2(n549), .ZN(G164) );
  NAND2_X1 U611 ( .A1(G91), .A2(n627), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G65), .A2(n628), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G78), .A2(n631), .ZN(n553) );
  XNOR2_X1 U615 ( .A(KEYINPUT67), .B(n553), .ZN(n554) );
  NOR2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n632), .A2(G53), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(G299) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n558) );
  XOR2_X1 U620 ( .A(n558), .B(KEYINPUT10), .Z(n916) );
  NAND2_X1 U621 ( .A1(n916), .A2(G567), .ZN(n559) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  NAND2_X1 U623 ( .A1(G56), .A2(n628), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT14), .B(n560), .Z(n566) );
  NAND2_X1 U625 ( .A1(n627), .A2(G81), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G68), .A2(n631), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT13), .B(n564), .Z(n565) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n632), .A2(G43), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n1008) );
  XOR2_X1 U633 ( .A(G860), .B(KEYINPUT68), .Z(n581) );
  NOR2_X1 U634 ( .A1(n1008), .A2(n581), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT69), .ZN(G153) );
  XOR2_X1 U636 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U637 ( .A1(G868), .A2(G301), .ZN(n578) );
  NAND2_X1 U638 ( .A1(G92), .A2(n627), .ZN(n571) );
  NAND2_X1 U639 ( .A1(G66), .A2(n628), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G79), .A2(n631), .ZN(n573) );
  NAND2_X1 U642 ( .A1(G54), .A2(n632), .ZN(n572) );
  NAND2_X1 U643 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U645 ( .A(KEYINPUT15), .B(n576), .ZN(n1005) );
  INV_X1 U646 ( .A(G868), .ZN(n646) );
  NAND2_X1 U647 ( .A1(n1005), .A2(n646), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(G284) );
  NOR2_X1 U649 ( .A1(G286), .A2(n646), .ZN(n580) );
  NOR2_X1 U650 ( .A1(G868), .A2(G299), .ZN(n579) );
  NOR2_X1 U651 ( .A1(n580), .A2(n579), .ZN(G297) );
  NAND2_X1 U652 ( .A1(n581), .A2(G559), .ZN(n582) );
  INV_X1 U653 ( .A(n1005), .ZN(n849) );
  NAND2_X1 U654 ( .A1(n582), .A2(n849), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT72), .ZN(n584) );
  XNOR2_X1 U656 ( .A(KEYINPUT16), .B(n584), .ZN(G148) );
  NOR2_X1 U657 ( .A1(G868), .A2(n1008), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G868), .A2(n849), .ZN(n585) );
  NOR2_X1 U659 ( .A1(G559), .A2(n585), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n587), .A2(n586), .ZN(G282) );
  NAND2_X1 U661 ( .A1(G123), .A2(n878), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n588), .B(KEYINPUT18), .ZN(n591) );
  NAND2_X1 U663 ( .A1(G99), .A2(n882), .ZN(n589) );
  XOR2_X1 U664 ( .A(KEYINPUT73), .B(n589), .Z(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G111), .A2(n879), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G135), .A2(n592), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n929) );
  XNOR2_X1 U670 ( .A(n929), .B(G2096), .ZN(n597) );
  INV_X1 U671 ( .A(G2100), .ZN(n827) );
  NAND2_X1 U672 ( .A1(n597), .A2(n827), .ZN(G156) );
  NAND2_X1 U673 ( .A1(G88), .A2(n627), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G62), .A2(n628), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G50), .A2(n632), .ZN(n600) );
  XNOR2_X1 U677 ( .A(KEYINPUT77), .B(n600), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n631), .A2(G75), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(G303) );
  NAND2_X1 U681 ( .A1(G86), .A2(n627), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G61), .A2(n628), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n631), .A2(G73), .ZN(n607) );
  XOR2_X1 U685 ( .A(KEYINPUT2), .B(n607), .Z(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n632), .A2(G48), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(G305) );
  NAND2_X1 U689 ( .A1(G49), .A2(n632), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G87), .A2(n612), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n628), .A2(n615), .ZN(n618) );
  NAND2_X1 U693 ( .A1(G74), .A2(G651), .ZN(n616) );
  XOR2_X1 U694 ( .A(KEYINPUT75), .B(n616), .Z(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U696 ( .A(KEYINPUT76), .B(n619), .ZN(G288) );
  NAND2_X1 U697 ( .A1(G60), .A2(n628), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G47), .A2(n632), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G85), .A2(n627), .ZN(n622) );
  XOR2_X1 U701 ( .A(KEYINPUT66), .B(n622), .Z(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n631), .A2(G72), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(G290) );
  XOR2_X1 U705 ( .A(G303), .B(G305), .Z(n643) );
  XNOR2_X1 U706 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n639) );
  NAND2_X1 U707 ( .A1(G93), .A2(n627), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G67), .A2(n628), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G80), .A2(n631), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G55), .A2(n632), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U713 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U714 ( .A(KEYINPUT74), .B(n637), .Z(n823) );
  XNOR2_X1 U715 ( .A(G290), .B(n823), .ZN(n638) );
  XNOR2_X1 U716 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U717 ( .A(G288), .B(n640), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n641), .B(G299), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n643), .B(n642), .ZN(n846) );
  NAND2_X1 U720 ( .A1(G559), .A2(n849), .ZN(n644) );
  XNOR2_X1 U721 ( .A(n1008), .B(n644), .ZN(n821) );
  XNOR2_X1 U722 ( .A(n846), .B(n821), .ZN(n645) );
  NOR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n648) );
  NOR2_X1 U724 ( .A1(n823), .A2(G868), .ZN(n647) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(G295) );
  NAND2_X1 U726 ( .A1(G2078), .A2(G2084), .ZN(n649) );
  XOR2_X1 U727 ( .A(KEYINPUT20), .B(n649), .Z(n650) );
  NAND2_X1 U728 ( .A1(G2090), .A2(n650), .ZN(n651) );
  XNOR2_X1 U729 ( .A(KEYINPUT21), .B(n651), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n652), .A2(G2072), .ZN(n653) );
  XOR2_X1 U731 ( .A(KEYINPUT79), .B(n653), .Z(G158) );
  XNOR2_X1 U732 ( .A(KEYINPUT80), .B(G44), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n654), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U734 ( .A1(G237), .A2(G235), .ZN(n655) );
  NAND2_X1 U735 ( .A1(G120), .A2(n655), .ZN(n656) );
  XNOR2_X1 U736 ( .A(KEYINPUT81), .B(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n657), .A2(G108), .ZN(n825) );
  NAND2_X1 U738 ( .A1(G567), .A2(n825), .ZN(n662) );
  NOR2_X1 U739 ( .A1(G220), .A2(G219), .ZN(n658) );
  XOR2_X1 U740 ( .A(KEYINPUT22), .B(n658), .Z(n659) );
  NOR2_X1 U741 ( .A1(G218), .A2(n659), .ZN(n660) );
  NAND2_X1 U742 ( .A1(G96), .A2(n660), .ZN(n824) );
  NAND2_X1 U743 ( .A1(G2106), .A2(n824), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U745 ( .A(KEYINPUT82), .B(n663), .ZN(n845) );
  NAND2_X1 U746 ( .A1(G661), .A2(G483), .ZN(n664) );
  NOR2_X1 U747 ( .A1(n845), .A2(n664), .ZN(n818) );
  NAND2_X1 U748 ( .A1(n818), .A2(G36), .ZN(G176) );
  INV_X1 U749 ( .A(G303), .ZN(G166) );
  INV_X1 U750 ( .A(G8), .ZN(n683) );
  NAND2_X1 U751 ( .A1(G160), .A2(G40), .ZN(n761) );
  INV_X1 U752 ( .A(n761), .ZN(n665) );
  NOR2_X1 U753 ( .A1(G164), .A2(G1384), .ZN(n762) );
  NAND2_X1 U754 ( .A1(n665), .A2(n762), .ZN(n666) );
  XNOR2_X2 U755 ( .A(n666), .B(KEYINPUT64), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n689), .A2(G2090), .ZN(n668) );
  NAND2_X1 U757 ( .A1(n689), .A2(G8), .ZN(n760) );
  NOR2_X1 U758 ( .A1(G1971), .A2(n760), .ZN(n667) );
  NOR2_X1 U759 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U760 ( .A1(n669), .A2(G303), .ZN(n679) );
  INV_X1 U761 ( .A(n679), .ZN(n670) );
  OR2_X1 U762 ( .A1(n670), .A2(G286), .ZN(n714) );
  INV_X1 U763 ( .A(n714), .ZN(n681) );
  NOR2_X1 U764 ( .A1(n689), .A2(G2084), .ZN(n720) );
  NOR2_X1 U765 ( .A1(n721), .A2(n720), .ZN(n671) );
  NAND2_X1 U766 ( .A1(n671), .A2(G8), .ZN(n672) );
  XNOR2_X1 U767 ( .A(n672), .B(KEYINPUT30), .ZN(n673) );
  XNOR2_X1 U768 ( .A(n689), .B(KEYINPUT87), .ZN(n698) );
  XNOR2_X1 U769 ( .A(G2078), .B(KEYINPUT25), .ZN(n975) );
  NAND2_X1 U770 ( .A1(n698), .A2(n975), .ZN(n675) );
  INV_X1 U771 ( .A(G1961), .ZN(n1009) );
  NAND2_X1 U772 ( .A1(n689), .A2(n1009), .ZN(n674) );
  NAND2_X1 U773 ( .A1(n675), .A2(n674), .ZN(n712) );
  NOR2_X1 U774 ( .A1(G171), .A2(n712), .ZN(n676) );
  NOR2_X1 U775 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U776 ( .A(KEYINPUT31), .B(n678), .Z(n727) );
  AND2_X1 U777 ( .A1(n727), .A2(n679), .ZN(n680) );
  OR2_X1 U778 ( .A1(n681), .A2(n680), .ZN(n682) );
  OR2_X2 U779 ( .A1(n683), .A2(n682), .ZN(n718) );
  INV_X1 U780 ( .A(G1996), .ZN(n981) );
  NOR2_X1 U781 ( .A1(n689), .A2(n981), .ZN(n684) );
  XOR2_X1 U782 ( .A(n684), .B(KEYINPUT26), .Z(n686) );
  NAND2_X1 U783 ( .A1(n689), .A2(G1341), .ZN(n685) );
  NAND2_X1 U784 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U785 ( .A1(n1008), .A2(n687), .ZN(n688) );
  OR2_X1 U786 ( .A1(n849), .A2(n688), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n849), .A2(n688), .ZN(n693) );
  NAND2_X1 U788 ( .A1(G2067), .A2(n698), .ZN(n691) );
  NAND2_X1 U789 ( .A1(n689), .A2(G1348), .ZN(n690) );
  NAND2_X1 U790 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U791 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U793 ( .A(KEYINPUT89), .B(n696), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G2072), .A2(n698), .ZN(n697) );
  XOR2_X1 U795 ( .A(KEYINPUT27), .B(n697), .Z(n701) );
  INV_X1 U796 ( .A(n698), .ZN(n699) );
  NAND2_X1 U797 ( .A1(n699), .A2(G1956), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U799 ( .A1(G299), .A2(n705), .ZN(n702) );
  XNOR2_X1 U800 ( .A(n702), .B(KEYINPUT90), .ZN(n703) );
  NOR2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U802 ( .A1(G299), .A2(n705), .ZN(n706) );
  XOR2_X1 U803 ( .A(KEYINPUT28), .B(n706), .Z(n707) );
  NOR2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U805 ( .A1(G171), .A2(n712), .ZN(n713) );
  XNOR2_X1 U806 ( .A(n713), .B(KEYINPUT88), .ZN(n724) );
  AND2_X1 U807 ( .A1(n724), .A2(n714), .ZN(n715) );
  AND2_X1 U808 ( .A1(n715), .A2(G8), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n726), .A2(n716), .ZN(n717) );
  AND2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n719) );
  AND2_X1 U811 ( .A1(G8), .A2(n720), .ZN(n722) );
  OR2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n728) );
  INV_X1 U813 ( .A(n728), .ZN(n723) );
  AND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n730) );
  OR2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U817 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U818 ( .A(n731), .B(KEYINPUT92), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n733), .A2(n732), .ZN(n743) );
  NAND2_X1 U820 ( .A1(G8), .A2(G166), .ZN(n734) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n734), .ZN(n735) );
  XNOR2_X1 U822 ( .A(n735), .B(KEYINPUT95), .ZN(n736) );
  NAND2_X1 U823 ( .A1(n743), .A2(n736), .ZN(n737) );
  XNOR2_X1 U824 ( .A(n737), .B(KEYINPUT96), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n738), .A2(n760), .ZN(n739) );
  XNOR2_X1 U826 ( .A(n739), .B(KEYINPUT97), .ZN(n756) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n747) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n740) );
  NOR2_X1 U829 ( .A1(n747), .A2(n740), .ZN(n1006) );
  INV_X1 U830 ( .A(KEYINPUT33), .ZN(n741) );
  AND2_X1 U831 ( .A1(n1006), .A2(n741), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n753) );
  XOR2_X1 U833 ( .A(G1981), .B(G305), .Z(n1000) );
  INV_X1 U834 ( .A(n760), .ZN(n745) );
  NAND2_X1 U835 ( .A1(G288), .A2(G1976), .ZN(n744) );
  XOR2_X1 U836 ( .A(KEYINPUT93), .B(n744), .Z(n996) );
  AND2_X1 U837 ( .A1(n745), .A2(n996), .ZN(n746) );
  NOR2_X1 U838 ( .A1(KEYINPUT33), .A2(n746), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n747), .A2(KEYINPUT33), .ZN(n748) );
  NOR2_X1 U840 ( .A1(n760), .A2(n748), .ZN(n749) );
  NOR2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X1 U842 ( .A1(n1000), .A2(n751), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U844 ( .A(KEYINPUT94), .B(n754), .Z(n755) );
  NOR2_X2 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U846 ( .A(n757), .B(KEYINPUT98), .ZN(n804) );
  NOR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n758) );
  XOR2_X1 U848 ( .A(n758), .B(KEYINPUT24), .Z(n759) );
  NOR2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n802) );
  NOR2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n807) );
  NAND2_X1 U851 ( .A1(G129), .A2(n878), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G141), .A2(n592), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n882), .A2(G105), .ZN(n765) );
  XOR2_X1 U855 ( .A(KEYINPUT38), .B(n765), .Z(n766) );
  NOR2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n879), .A2(G117), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U859 ( .A(KEYINPUT85), .B(n770), .Z(n875) );
  NOR2_X1 U860 ( .A1(G1996), .A2(n875), .ZN(n771) );
  XOR2_X1 U861 ( .A(KEYINPUT99), .B(n771), .Z(n924) );
  NAND2_X1 U862 ( .A1(G119), .A2(n878), .ZN(n773) );
  NAND2_X1 U863 ( .A1(G107), .A2(n879), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G95), .A2(n882), .ZN(n775) );
  NAND2_X1 U866 ( .A1(G131), .A2(n592), .ZN(n774) );
  NAND2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n776) );
  OR2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n865) );
  NAND2_X1 U869 ( .A1(G1991), .A2(n865), .ZN(n779) );
  NAND2_X1 U870 ( .A1(G1996), .A2(n875), .ZN(n778) );
  NAND2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n922) );
  NAND2_X1 U872 ( .A1(n807), .A2(n922), .ZN(n780) );
  XNOR2_X1 U873 ( .A(KEYINPUT86), .B(n780), .ZN(n806) );
  INV_X1 U874 ( .A(n806), .ZN(n783) );
  NOR2_X1 U875 ( .A1(G1986), .A2(G290), .ZN(n781) );
  NOR2_X1 U876 ( .A1(G1991), .A2(n865), .ZN(n930) );
  NOR2_X1 U877 ( .A1(n781), .A2(n930), .ZN(n782) );
  NOR2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U879 ( .A1(n924), .A2(n784), .ZN(n785) );
  XNOR2_X1 U880 ( .A(n785), .B(KEYINPUT39), .ZN(n797) );
  XNOR2_X1 U881 ( .A(KEYINPUT37), .B(G2067), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G104), .A2(n882), .ZN(n787) );
  NAND2_X1 U883 ( .A1(G140), .A2(n592), .ZN(n786) );
  NAND2_X1 U884 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n788), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n878), .A2(G128), .ZN(n789) );
  XNOR2_X1 U887 ( .A(KEYINPUT83), .B(n789), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n879), .A2(G116), .ZN(n790) );
  XOR2_X1 U889 ( .A(KEYINPUT84), .B(n790), .Z(n791) );
  NOR2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U891 ( .A(n793), .B(KEYINPUT35), .ZN(n794) );
  NOR2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n796), .ZN(n894) );
  NOR2_X1 U894 ( .A1(n798), .A2(n894), .ZN(n936) );
  NAND2_X1 U895 ( .A1(n807), .A2(n936), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n797), .A2(n805), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n798), .A2(n894), .ZN(n938) );
  NAND2_X1 U898 ( .A1(n799), .A2(n938), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n807), .A2(n800), .ZN(n801) );
  XOR2_X1 U900 ( .A(KEYINPUT100), .B(n801), .Z(n811) );
  NOR2_X1 U901 ( .A1(n802), .A2(n811), .ZN(n803) );
  NAND2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n809) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n995) );
  AND2_X1 U905 ( .A1(n995), .A2(n807), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  OR2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U909 ( .A(n814), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n916), .ZN(G217) );
  NAND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n816) );
  INV_X1 U912 ( .A(G661), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U914 ( .A(n817), .B(KEYINPUT103), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G1), .A2(G3), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n820), .B(KEYINPUT104), .ZN(G188) );
  XNOR2_X1 U918 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  XOR2_X1 U919 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  NOR2_X1 U921 ( .A1(G860), .A2(n821), .ZN(n822) );
  XOR2_X1 U922 ( .A(n823), .B(n822), .Z(G145) );
  INV_X1 U923 ( .A(G108), .ZN(G238) );
  NOR2_X1 U924 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U925 ( .A(n826), .B(KEYINPUT107), .Z(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U927 ( .A(n827), .B(G2096), .ZN(n829) );
  XNOR2_X1 U928 ( .A(KEYINPUT42), .B(G2678), .ZN(n828) );
  XNOR2_X1 U929 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U930 ( .A(KEYINPUT43), .B(G2090), .Z(n831) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U933 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2084), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(G227) );
  XOR2_X1 U936 ( .A(G1976), .B(G1971), .Z(n837) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1966), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U939 ( .A(n838), .B(KEYINPUT41), .Z(n840) );
  XOR2_X1 U940 ( .A(G1991), .B(n981), .Z(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n844) );
  XNOR2_X1 U942 ( .A(G2474), .B(n1009), .ZN(n842) );
  XNOR2_X1 U943 ( .A(G1981), .B(G1956), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(G229) );
  INV_X1 U946 ( .A(n845), .ZN(G319) );
  XNOR2_X1 U947 ( .A(G286), .B(n846), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n1008), .B(G171), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n849), .B(KEYINPUT115), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  NOR2_X1 U952 ( .A1(G37), .A2(n852), .ZN(G397) );
  NAND2_X1 U953 ( .A1(G100), .A2(n882), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G112), .A2(n879), .ZN(n853) );
  NAND2_X1 U955 ( .A1(n854), .A2(n853), .ZN(n861) );
  NAND2_X1 U956 ( .A1(G124), .A2(n878), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n855), .B(KEYINPUT108), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G136), .A2(n592), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U961 ( .A(KEYINPUT109), .B(n859), .Z(n860) );
  NOR2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U963 ( .A(KEYINPUT110), .B(n862), .ZN(G162) );
  XOR2_X1 U964 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n864) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n877) );
  NAND2_X1 U968 ( .A1(G103), .A2(n882), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G139), .A2(n592), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G127), .A2(n878), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G115), .A2(n879), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n871), .Z(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n917) );
  XOR2_X1 U976 ( .A(n929), .B(n917), .Z(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n893) );
  XNOR2_X1 U979 ( .A(G164), .B(G160), .ZN(n890) );
  NAND2_X1 U980 ( .A1(G130), .A2(n878), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G118), .A2(n879), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G106), .A2(n882), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G142), .A2(n592), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U986 ( .A(KEYINPUT45), .B(n885), .ZN(n886) );
  XNOR2_X1 U987 ( .A(KEYINPUT111), .B(n886), .ZN(n887) );
  NOR2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U990 ( .A(G162), .B(n891), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n895) );
  XOR2_X1 U992 ( .A(n895), .B(n894), .Z(n896) );
  NOR2_X1 U993 ( .A1(G37), .A2(n896), .ZN(n897) );
  XNOR2_X1 U994 ( .A(KEYINPUT114), .B(n897), .ZN(G395) );
  NOR2_X1 U995 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n912) );
  XNOR2_X1 U998 ( .A(G2454), .B(G2443), .ZN(n909) );
  XOR2_X1 U999 ( .A(G2430), .B(KEYINPUT102), .Z(n901) );
  XNOR2_X1 U1000 ( .A(G2446), .B(KEYINPUT101), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U1002 ( .A(G2451), .B(G2427), .Z(n903) );
  XNOR2_X1 U1003 ( .A(G1341), .B(G1348), .ZN(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1005 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1006 ( .A(G2435), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(n910), .A2(G14), .ZN(n915) );
  NAND2_X1 U1010 ( .A1(n915), .A2(G319), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G397), .A2(G395), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(n915), .ZN(G401) );
  INV_X1 U1016 ( .A(n916), .ZN(G223) );
  XNOR2_X1 U1017 ( .A(G164), .B(G2078), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G2072), .B(n917), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n918), .B(KEYINPUT120), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(KEYINPUT50), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n928) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1025 ( .A(KEYINPUT51), .B(n926), .Z(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n941) );
  XOR2_X1 U1027 ( .A(G160), .B(G2084), .Z(n933) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(KEYINPUT117), .B(n931), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1031 ( .A(KEYINPUT118), .B(n934), .Z(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1033 ( .A(KEYINPUT119), .B(n937), .Z(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n942), .ZN(n943) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n989) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n989), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(G29), .ZN(n1023) );
  XOR2_X1 U1040 ( .A(G16), .B(KEYINPUT126), .Z(n967) );
  XOR2_X1 U1041 ( .A(G1986), .B(G24), .Z(n948) );
  XNOR2_X1 U1042 ( .A(G1971), .B(G22), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G23), .B(G1976), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n950), .B(n949), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G21), .ZN(n952) );
  XOR2_X1 U1049 ( .A(n1009), .B(G5), .Z(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n964) );
  XOR2_X1 U1052 ( .A(G1348), .B(KEYINPUT59), .Z(n955) );
  XNOR2_X1 U1053 ( .A(G4), .B(n955), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G20), .B(G1956), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G1981), .B(G6), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(G19), .B(G1341), .ZN(n958) );
  NOR2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(KEYINPUT60), .B(n962), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(n965), .B(KEYINPUT61), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n968), .ZN(n1021) );
  XOR2_X1 U1065 ( .A(G2090), .B(G35), .Z(n971) );
  XOR2_X1 U1066 ( .A(KEYINPUT54), .B(G34), .Z(n969) );
  XNOR2_X1 U1067 ( .A(n969), .B(G2084), .ZN(n970) );
  NAND2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n987) );
  XNOR2_X1 U1069 ( .A(G1991), .B(G25), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(G26), .B(G2067), .ZN(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n980) );
  XOR2_X1 U1072 ( .A(G2072), .B(G33), .Z(n974) );
  NAND2_X1 U1073 ( .A1(n974), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(G27), .B(n975), .ZN(n976) );
  XNOR2_X1 U1075 ( .A(KEYINPUT121), .B(n976), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1078 ( .A(G32), .B(n981), .Z(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(KEYINPUT122), .B(n984), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(KEYINPUT53), .B(n985), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(n989), .B(n988), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(G29), .A2(n990), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(KEYINPUT123), .B(n991), .ZN(n1019) );
  XNOR2_X1 U1086 ( .A(G16), .B(KEYINPUT56), .ZN(n1017) );
  NAND2_X1 U1087 ( .A1(G1971), .A2(G303), .ZN(n993) );
  XOR2_X1 U1088 ( .A(G1956), .B(G299), .Z(n992) );
  NAND2_X1 U1089 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1090 ( .A1(n995), .A2(n994), .ZN(n997) );
  NAND2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n1002) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G168), .ZN(n998) );
  XNOR2_X1 U1094 ( .A(n998), .B(KEYINPUT124), .ZN(n999) );
  NAND2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1096 ( .A(n1002), .B(n1001), .Z(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1015) );
  XOR2_X1 U1098 ( .A(n1005), .B(G1348), .Z(n1007) );
  NAND2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(n1008), .B(G1341), .Z(n1011) );
  XOR2_X1 U1101 ( .A(G171), .B(n1009), .Z(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1024), .ZN(G150) );
  INV_X1 U1110 ( .A(G150), .ZN(G311) );
endmodule

