//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  OR2_X1    g001(.A1(G127gat), .A2(G134gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G127gat), .A2(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n205), .B1(new_n206), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT68), .B1(new_n207), .B2(G113gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(new_n209), .A3(G120gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n216), .A3(new_n208), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT69), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n214), .A2(new_n216), .A3(new_n219), .A4(new_n208), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT70), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n203), .A2(KEYINPUT70), .A3(new_n204), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT1), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n221), .A2(new_n222), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n221), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n213), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT27), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT27), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G183gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n233), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n230), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n232), .A2(new_n238), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT28), .A3(new_n235), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g042(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NOR2_X1   g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247));
  OAI22_X1  g046(.A1(new_n244), .A2(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT67), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n250));
  OAI221_X1 g049(.A(new_n250), .B1(new_n247), .B2(new_n246), .C1(new_n244), .C2(new_n245), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n246), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G183gat), .A2(G190gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n243), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(KEYINPUT24), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT24), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(G183gat), .A3(G190gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(G183gat), .B2(G190gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT64), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n267), .A2(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n264), .A2(new_n265), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n268), .ZN(new_n275));
  NOR3_X1   g074(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n276));
  OAI22_X1  g075(.A1(new_n275), .A2(new_n276), .B1(new_n244), .B2(new_n245), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n262), .B1(new_n256), .B2(new_n258), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT25), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n255), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT72), .B1(new_n229), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n221), .A2(new_n226), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n221), .A2(new_n226), .A3(new_n222), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n274), .A2(new_n279), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n240), .A2(new_n242), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n253), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n286), .A2(new_n289), .A3(new_n290), .A4(new_n213), .ZN(new_n291));
  NAND2_X1  g090(.A1(G227gat), .A2(G233gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n229), .A2(new_n281), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n282), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n294), .B(KEYINPUT34), .Z(new_n295));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n282), .A2(new_n291), .A3(new_n293), .ZN(new_n297));
  INV_X1    g096(.A(new_n292), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT33), .B1(new_n297), .B2(new_n298), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301));
  XNOR2_X1  g100(.A(G15gat), .B(G43gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G71gat), .B(G99gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NOR4_X1   g103(.A1(new_n299), .A2(new_n300), .A3(new_n301), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(new_n298), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT33), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(KEYINPUT32), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT73), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n304), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT33), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n316), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n295), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n306), .A2(new_n307), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n309), .A2(new_n320), .A3(new_n312), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n301), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n308), .A2(KEYINPUT73), .A3(new_n309), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n322), .A2(new_n318), .A3(new_n295), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n202), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G141gat), .B(G148gat), .Z(new_n327));
  OR2_X1    g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(KEYINPUT2), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n327), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G141gat), .B(G148gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n329), .B(new_n328), .C1(new_n333), .C2(KEYINPUT2), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  XOR2_X1   g135(.A(G211gat), .B(G218gat), .Z(new_n337));
  AOI21_X1  g136(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n338));
  INV_X1    g137(.A(G197gat), .ZN(new_n339));
  INV_X1    g138(.A(G204gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G197gat), .A2(G204gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT76), .B1(new_n348), .B2(new_n338), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n337), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n348), .A2(KEYINPUT76), .A3(new_n338), .ZN(new_n351));
  INV_X1    g150(.A(new_n337), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n336), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n335), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n342), .ZN(new_n357));
  INV_X1    g156(.A(new_n338), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n344), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n352), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n337), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n332), .A2(new_n334), .A3(new_n355), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(new_n336), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT82), .B1(new_n356), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n336), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT3), .B1(new_n362), .B2(new_n336), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(new_n335), .ZN(new_n371));
  INV_X1    g170(.A(G228gat), .ZN(new_n372));
  INV_X1    g171(.A(G233gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n365), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(KEYINPUT82), .B(new_n374), .C1(new_n356), .C2(new_n364), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(G22gat), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT31), .B(G50gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n376), .A2(new_n377), .ZN(new_n385));
  INV_X1    g184(.A(G22gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n378), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n387), .A2(KEYINPUT83), .A3(new_n378), .A4(new_n383), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G226gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n373), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(new_n289), .B2(KEYINPUT29), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n281), .B2(new_n393), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT78), .B(new_n394), .C1(new_n255), .C2(new_n280), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n362), .B(new_n395), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n281), .B2(new_n336), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n289), .B2(new_n394), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n281), .A2(KEYINPUT77), .A3(new_n393), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n404), .B2(new_n362), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n399), .B(new_n408), .C1(new_n404), .C2(new_n362), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(KEYINPUT30), .A3(new_n411), .ZN(new_n412));
  OR3_X1    g211(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n409), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT35), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT0), .ZN(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n335), .A2(new_n355), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n332), .A2(new_n334), .A3(new_n355), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n229), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n213), .B(new_n335), .C1(new_n227), .C2(new_n228), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n286), .A2(KEYINPUT4), .A3(new_n213), .A4(new_n335), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT79), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT79), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n428), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n432), .A3(new_n431), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n335), .B1(new_n286), .B2(new_n213), .ZN(new_n439));
  INV_X1    g238(.A(new_n429), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n422), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n438), .A2(new_n441), .A3(KEYINPUT5), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n420), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444));
  INV_X1    g243(.A(new_n428), .ZN(new_n445));
  INV_X1    g244(.A(new_n436), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n438), .A2(new_n441), .A3(KEYINPUT5), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n419), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n443), .A2(new_n444), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n419), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  INV_X1    g252(.A(new_n451), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n450), .A2(new_n451), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT86), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n415), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n322), .A2(new_n318), .A3(new_n323), .ZN(new_n460));
  INV_X1    g259(.A(new_n295), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(KEYINPUT87), .A3(new_n324), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n326), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n326), .A2(new_n459), .A3(KEYINPUT88), .A4(new_n463), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n460), .A2(new_n468), .A3(new_n461), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n460), .B2(new_n461), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT81), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n453), .B1(new_n457), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n451), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n473), .A2(new_n474), .B1(new_n453), .B2(new_n454), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n412), .A2(new_n413), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n391), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n325), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n471), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n466), .A2(new_n467), .B1(KEYINPUT35), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n389), .A2(KEYINPUT84), .A3(new_n390), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT84), .B1(new_n389), .B2(new_n390), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n475), .B2(new_n477), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n324), .A2(KEYINPUT36), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n469), .A2(new_n470), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT36), .B1(new_n462), .B2(new_n324), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n456), .A2(new_n458), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n405), .A2(KEYINPUT37), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n409), .B1(new_n405), .B2(KEYINPUT37), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n366), .B(new_n395), .C1(new_n397), .C2(new_n398), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(KEYINPUT37), .C1(new_n404), .C2(new_n366), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT38), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n494), .B(new_n411), .C1(new_n493), .C2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n229), .A2(new_n425), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n446), .B2(new_n447), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n422), .ZN(new_n503));
  OR3_X1    g302(.A1(new_n439), .A2(new_n440), .A3(new_n422), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT39), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT39), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n506), .A3(new_n422), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n419), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n505), .A2(KEYINPUT40), .A3(new_n419), .A4(new_n507), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n510), .A2(new_n443), .A3(new_n477), .A4(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n512), .A2(new_n391), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n490), .A2(KEYINPUT85), .B1(new_n500), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n486), .B(new_n515), .C1(new_n488), .C2(new_n489), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n482), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G36gat), .ZN(new_n519));
  AND2_X1   g318(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n527));
  XNOR2_X1  g326(.A(G43gat), .B(G50gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(KEYINPUT17), .B2(new_n531), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(G1gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G1gat), .B2(new_n535), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n531), .A2(new_n540), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT18), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n531), .B(new_n540), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n544), .A2(new_n545), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G169gat), .B(G197gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT12), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n546), .A2(new_n550), .A3(new_n551), .A4(new_n558), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n564), .B1(new_n531), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n534), .B2(new_n574), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT95), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n576), .B(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT94), .Z(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n579), .B(new_n583), .Z(new_n584));
  XOR2_X1   g383(.A(G57gat), .B(G64gat), .Z(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G71gat), .B(G78gat), .Z(new_n591));
  OR2_X1    g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  OAI21_X1  g397(.A(new_n540), .B1(new_n595), .B2(new_n594), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT93), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT92), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n600), .B(new_n607), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n584), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n573), .B(new_n594), .Z(new_n610));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT96), .Z(new_n614));
  OR2_X1    g413(.A1(new_n610), .A2(KEYINPUT10), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n573), .A2(KEYINPUT10), .A3(new_n593), .A4(new_n592), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n611), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n618), .B1(new_n617), .B2(new_n611), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G120gat), .B(G148gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT97), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n617), .A2(new_n611), .ZN(new_n628));
  INV_X1    g427(.A(new_n626), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n609), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n518), .A2(new_n562), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n475), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT99), .B(G1gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(G1324gat));
  INV_X1    g436(.A(new_n633), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n539), .B1(new_n638), .B2(new_n477), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT16), .B(G8gat), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n633), .A2(new_n476), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT42), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(KEYINPUT42), .B2(new_n641), .ZN(G1325gat));
  NOR2_X1   g442(.A1(new_n488), .A2(new_n489), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(G15gat), .B1(new_n633), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n326), .A2(new_n463), .ZN(new_n647));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n633), .B2(new_n649), .ZN(G1326gat));
  INV_X1    g449(.A(new_n485), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n633), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  INV_X1    g454(.A(new_n584), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n512), .B(new_n391), .C1(new_n491), .C2(new_n499), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n657), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n655), .B(new_n656), .C1(new_n482), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n490), .A2(KEYINPUT85), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n516), .A3(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n466), .A2(new_n467), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n584), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  OAI211_X1 g465(.A(KEYINPUT100), .B(new_n660), .C1(new_n666), .C2(new_n655), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n668), .B(KEYINPUT44), .C1(new_n517), .C2(new_n584), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n562), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(new_n608), .A3(new_n631), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674), .B2(new_n634), .ZN(new_n675));
  INV_X1    g474(.A(new_n666), .ZN(new_n676));
  INV_X1    g475(.A(new_n673), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n523), .A3(new_n475), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT45), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n675), .A2(new_n680), .ZN(G1328gat));
  NAND3_X1  g480(.A1(new_n678), .A2(new_n519), .A3(new_n477), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT46), .Z(new_n683));
  OAI21_X1  g482(.A(G36gat), .B1(new_n674), .B2(new_n476), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1329gat));
  NAND4_X1  g484(.A1(new_n667), .A2(new_n644), .A3(new_n669), .A4(new_n673), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(G43gat), .ZN(new_n687));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n666), .A2(new_n688), .A3(new_n647), .A4(new_n673), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(KEYINPUT47), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(KEYINPUT101), .Z(new_n691));
  AOI21_X1  g490(.A(KEYINPUT47), .B1(new_n691), .B2(new_n687), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n692), .A2(KEYINPUT102), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(KEYINPUT102), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(G1330gat));
  OAI211_X1 g494(.A(KEYINPUT48), .B(G50gat), .C1(new_n674), .C2(new_n391), .ZN(new_n696));
  NOR4_X1   g495(.A1(new_n676), .A2(G50gat), .A3(new_n651), .A4(new_n677), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n671), .A2(new_n485), .A3(new_n673), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n702), .A2(G50gat), .B1(new_n698), .B2(new_n697), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(KEYINPUT48), .B2(new_n703), .ZN(G1331gat));
  NAND2_X1  g503(.A1(new_n665), .A2(new_n658), .ZN(new_n705));
  INV_X1    g504(.A(new_n630), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n622), .B2(new_n626), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n609), .A2(new_n562), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n475), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(G57gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1332gat));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n477), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT49), .B(G64gat), .Z(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n714), .B2(new_n716), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n709), .B2(new_n645), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n647), .A2(new_n587), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1334gat));
  NAND2_X1  g521(.A1(new_n710), .A2(new_n485), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g523(.A1(new_n562), .A2(new_n608), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n656), .B(new_n725), .C1(new_n482), .C2(new_n659), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(new_n568), .A3(new_n475), .A4(new_n631), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n562), .A2(new_n608), .A3(new_n707), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n671), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT106), .B1(new_n731), .B2(new_n634), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G85gat), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n731), .A2(KEYINPUT106), .A3(new_n634), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n729), .B1(new_n733), .B2(new_n734), .ZN(G1336gat));
  OAI21_X1  g534(.A(G92gat), .B1(new_n731), .B2(new_n476), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n707), .A2(G92gat), .A3(new_n476), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT52), .B1(new_n728), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT108), .B1(new_n726), .B2(KEYINPUT107), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(new_n727), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n740), .A2(new_n727), .B1(new_n726), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n737), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n736), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n731), .B2(new_n645), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n707), .A2(G99gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n728), .A2(new_n647), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1338gat));
  NAND4_X1  g551(.A1(new_n667), .A2(new_n485), .A3(new_n669), .A4(new_n730), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G106gat), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n707), .A2(G106gat), .A3(new_n391), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n744), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT53), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n667), .A2(new_n479), .A3(new_n669), .A4(new_n730), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G106gat), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n762), .A2(KEYINPUT53), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(KEYINPUT53), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n728), .A2(new_n755), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n760), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n761), .B1(new_n760), .B2(new_n765), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n758), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n758), .B(KEYINPUT111), .C1(new_n766), .C2(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1339gat));
  INV_X1    g571(.A(new_n608), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n774), .A2(KEYINPUT113), .B1(new_n547), .B2(new_n549), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n557), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n631), .A2(new_n561), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n628), .A2(KEYINPUT98), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n619), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n617), .B2(new_n611), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n615), .A2(new_n612), .A3(new_n616), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n629), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(KEYINPUT55), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n630), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(new_n781), .B2(new_n784), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n778), .B1(new_n792), .B2(new_n672), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n584), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n561), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n792), .A2(new_n584), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n773), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n632), .A2(new_n672), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n799), .A2(new_n471), .A3(new_n480), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n634), .A2(new_n477), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT114), .Z(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n209), .A3(new_n562), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n485), .B1(new_n797), .B2(new_n798), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n805), .A2(new_n647), .A3(new_n801), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n672), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(G1340gat));
  NAND3_X1  g608(.A1(new_n803), .A2(new_n207), .A3(new_n631), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n207), .B1(new_n806), .B2(new_n631), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT115), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1341gat));
  OAI21_X1  g612(.A(G127gat), .B1(new_n807), .B2(new_n773), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n773), .A2(G127gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n802), .B2(new_n815), .ZN(G1342gat));
  NAND2_X1  g615(.A1(new_n656), .A2(new_n476), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n634), .A3(G134gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT56), .Z(new_n820));
  OAI21_X1  g619(.A(G134gat), .B1(new_n807), .B2(new_n584), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1343gat));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n799), .A2(new_n823), .A3(new_n479), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n644), .A2(new_n634), .A3(new_n477), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n631), .A2(new_n826), .A3(new_n561), .A4(new_n777), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT116), .B1(new_n795), .B2(new_n707), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n786), .B2(new_n788), .ZN(new_n831));
  INV_X1    g630(.A(new_n788), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n832), .A2(KEYINPUT117), .A3(new_n630), .A4(new_n785), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n833), .A3(new_n562), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n656), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n773), .B1(new_n835), .B2(new_n796), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n651), .B1(new_n836), .B2(new_n798), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n824), .B(new_n825), .C1(new_n823), .C2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G141gat), .B1(new_n838), .B2(new_n672), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n839), .B2(KEYINPUT119), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n391), .B1(new_n797), .B2(new_n798), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n825), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n672), .A2(G141gat), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT118), .Z(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n840), .B(new_n846), .Z(G1344gat));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n848), .B(G148gat), .C1(new_n838), .C2(new_n707), .ZN(new_n849));
  INV_X1    g648(.A(new_n837), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n851), .A3(new_n823), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n841), .A2(KEYINPUT57), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT120), .B1(new_n837), .B2(KEYINPUT57), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n825), .A2(new_n631), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G148gat), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT121), .B1(new_n858), .B2(KEYINPUT59), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n860), .B(new_n848), .C1(new_n857), .C2(G148gat), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n849), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(G148gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n842), .A2(new_n863), .A3(new_n631), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1345gat));
  OAI21_X1  g664(.A(G155gat), .B1(new_n838), .B2(new_n773), .ZN(new_n866));
  INV_X1    g665(.A(G155gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n842), .A2(new_n867), .A3(new_n608), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n838), .B2(new_n584), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n817), .A2(new_n634), .A3(G162gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n841), .A2(new_n645), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n475), .A2(new_n476), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n800), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(G169gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n562), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT123), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n805), .A2(new_n647), .A3(new_n875), .ZN(new_n880));
  OAI21_X1  g679(.A(G169gat), .B1(new_n880), .B2(new_n672), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1348gat));
  INV_X1    g681(.A(G176gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n876), .A2(new_n883), .A3(new_n631), .ZN(new_n884));
  OAI21_X1  g683(.A(G176gat), .B1(new_n880), .B2(new_n707), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1349gat));
  NAND3_X1  g685(.A1(new_n876), .A2(new_n241), .A3(new_n608), .ZN(new_n887));
  OAI21_X1  g686(.A(G183gat), .B1(new_n880), .B2(new_n773), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n876), .A2(new_n235), .A3(new_n656), .ZN(new_n891));
  OAI21_X1  g690(.A(G190gat), .B1(new_n880), .B2(new_n584), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(KEYINPUT61), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(KEYINPUT61), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT124), .ZN(G1351gat));
  NAND2_X1  g695(.A1(new_n645), .A2(new_n875), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n841), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(G197gat), .B1(new_n899), .B2(new_n562), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n855), .A2(new_n898), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n672), .A2(new_n339), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(G1352gat));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n340), .A3(new_n631), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT62), .Z(new_n906));
  OAI21_X1  g705(.A(G204gat), .B1(new_n901), .B2(new_n707), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1353gat));
  INV_X1    g707(.A(G211gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n899), .A2(new_n909), .A3(new_n608), .ZN(new_n910));
  OAI21_X1  g709(.A(G211gat), .B1(new_n901), .B2(new_n773), .ZN(new_n911));
  NOR2_X1   g710(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n911), .A2(new_n912), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(G1354gat));
  AOI21_X1  g716(.A(G218gat), .B1(new_n899), .B2(new_n656), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n656), .A2(G218gat), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT127), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n902), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n901), .A2(KEYINPUT126), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(G1355gat));
endmodule


