//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n205), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT29), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT3), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT74), .ZN(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(G155gat), .B2(G162gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G155gat), .B(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n218), .A2(KEYINPUT2), .ZN(new_n227));
  INV_X1    g026(.A(G141gat), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n224), .A3(new_n219), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n204), .B1(new_n217), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n215), .B(KEYINPUT71), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n232), .A2(new_n224), .A3(new_n219), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n224), .B1(new_n232), .B2(new_n219), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n216), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n235), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n238), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT76), .B1(new_n226), .B2(new_n233), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT29), .B1(new_n213), .B2(new_n214), .ZN(new_n246));
  OAI22_X1  g045(.A1(new_n244), .A2(new_n245), .B1(KEYINPUT3), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI221_X1 g048(.A(KEYINPUT78), .B1(new_n246), .B2(KEYINPUT3), .C1(new_n244), .C2(new_n245), .ZN(new_n250));
  INV_X1    g049(.A(new_n215), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT3), .B1(new_n226), .B2(new_n233), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(KEYINPUT29), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT79), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n241), .A2(new_n255), .A3(new_n251), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n249), .A2(new_n250), .A3(new_n254), .A4(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n203), .B(KEYINPUT77), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n242), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G22gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n202), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT31), .B(G50gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n257), .A2(new_n258), .ZN(new_n266));
  INV_X1    g065(.A(new_n242), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n260), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI211_X1 g067(.A(G22gat), .B(new_n242), .C1(new_n257), .C2(new_n258), .ZN(new_n269));
  OAI22_X1  g068(.A1(new_n261), .A2(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n267), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G22gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n259), .A2(new_n260), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n202), .A3(new_n273), .A4(new_n264), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276));
  AND2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT24), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n277), .A2(new_n278), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT24), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT23), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n279), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n285), .B2(KEYINPUT23), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n290), .B(KEYINPUT67), .C1(G169gat), .C2(G176gat), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT25), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n280), .A2(KEYINPUT27), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G183gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n296), .A3(new_n281), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT68), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n277), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G169gat), .ZN(new_n301));
  INV_X1    g100(.A(G176gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT69), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT26), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n285), .A2(KEYINPUT69), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n281), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n300), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n307), .B1(new_n283), .B2(KEYINPUT24), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n277), .A2(new_n278), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(new_n282), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT65), .B(G169gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT23), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n289), .A2(new_n291), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n315), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n293), .A2(new_n312), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n293), .A2(new_n312), .A3(new_n323), .A4(KEYINPUT73), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n276), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n276), .B(KEYINPUT72), .Z(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n324), .B2(new_n216), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n236), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n329), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n322), .A2(new_n284), .A3(new_n279), .A4(new_n286), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n316), .A2(new_n317), .A3(new_n290), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n334), .A2(new_n319), .B1(new_n289), .B2(new_n291), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n279), .A2(new_n284), .A3(new_n321), .ZN(new_n336));
  AOI22_X1  g135(.A1(KEYINPUT25), .A2(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n332), .B1(new_n337), .B2(new_n312), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n251), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n326), .B2(new_n327), .ZN(new_n340));
  INV_X1    g139(.A(new_n276), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  NAND3_X1  g144(.A1(new_n331), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n331), .A2(new_n342), .A3(KEYINPUT30), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n342), .ZN(new_n350));
  INV_X1    g149(.A(new_n345), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n348), .A2(new_n352), .A3(KEYINPUT81), .A4(new_n349), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G15gat), .B(G43gat), .Z(new_n358));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT64), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n364));
  INV_X1    g163(.A(G113gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(G120gat), .ZN(new_n366));
  INV_X1    g165(.A(G120gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(G113gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n364), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G127gat), .B(G134gat), .Z(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n372), .B(new_n364), .C1(new_n366), .C2(new_n368), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n324), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n374), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n376), .A2(new_n293), .A3(new_n312), .A4(new_n323), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n363), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n360), .B1(new_n378), .B2(KEYINPUT33), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT32), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n375), .A2(new_n377), .ZN(new_n383));
  AOI221_X4 g182(.A(new_n380), .B1(KEYINPUT33), .B2(new_n360), .C1(new_n383), .C2(new_n362), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n375), .A2(new_n363), .A3(new_n377), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT70), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT34), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n382), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n376), .B1(new_n337), .B2(new_n312), .ZN(new_n390));
  AND4_X1   g189(.A1(new_n376), .A2(new_n293), .A3(new_n312), .A4(new_n323), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n362), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT32), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT33), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n395), .A3(new_n360), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n389), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI22_X1  g197(.A1(new_n388), .A2(new_n398), .B1(new_n386), .B2(new_n385), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n387), .B1(new_n382), .B2(new_n384), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n385), .A2(new_n386), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n389), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n275), .A2(new_n357), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n376), .A2(new_n234), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n374), .B1(new_n226), .B2(new_n233), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n243), .B1(new_n238), .B2(new_n239), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n226), .A2(new_n233), .A3(KEYINPUT76), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n376), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n413), .A2(new_n415), .B1(new_n409), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n226), .A2(new_n233), .A3(KEYINPUT3), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n240), .A2(new_n418), .A3(new_n374), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n406), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT5), .B(new_n410), .C1(new_n417), .C2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n376), .A2(new_n234), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT4), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n411), .A2(new_n412), .A3(new_n376), .A4(new_n414), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT0), .ZN(new_n430));
  XNOR2_X1  g229(.A(G57gat), .B(G85gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT6), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n428), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n421), .A2(new_n427), .A3(new_n435), .A4(new_n432), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT35), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n353), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n275), .A2(new_n441), .A3(new_n404), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n405), .A2(new_n440), .B1(new_n442), .B2(KEYINPUT35), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT36), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n401), .B1(new_n400), .B2(new_n402), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n399), .A2(KEYINPUT36), .A3(new_n403), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(new_n448), .C1(new_n275), .C2(new_n441), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT37), .ZN(new_n451));
  INV_X1    g250(.A(new_n338), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n340), .B2(new_n341), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n251), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n328), .A2(new_n330), .ZN(new_n455));
  INV_X1    g254(.A(new_n236), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n451), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(KEYINPUT82), .B(KEYINPUT37), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n331), .A2(new_n342), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n345), .A2(KEYINPUT38), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n437), .A2(new_n438), .A3(new_n346), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n450), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n453), .A2(new_n251), .B1(new_n455), .B2(new_n456), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n461), .B(new_n462), .C1(new_n467), .C2(new_n451), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n439), .A2(new_n468), .A3(KEYINPUT83), .A4(new_n346), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n350), .A2(KEYINPUT37), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(new_n351), .A3(new_n461), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT38), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n408), .A2(new_n409), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n475), .B2(new_n406), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n418), .A2(new_n374), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n424), .A2(new_n425), .B1(new_n477), .B2(new_n240), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n478), .B2(new_n406), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n426), .A2(new_n419), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n474), .A3(new_n407), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n481), .A3(new_n433), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT40), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT40), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n479), .A2(new_n481), .A3(new_n484), .A4(new_n433), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n483), .A2(new_n485), .B1(new_n428), .B2(new_n432), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n355), .A2(new_n356), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n473), .A2(new_n275), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n449), .B1(new_n488), .B2(KEYINPUT84), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n473), .A2(new_n490), .A3(new_n275), .A4(new_n487), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n443), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT88), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G1gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(KEYINPUT89), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT16), .B1(new_n498), .B2(G1gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n493), .B(KEYINPUT88), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n496), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n505), .A3(G8gat), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n500), .B(new_n504), .C1(new_n501), .C2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G36gat), .ZN(new_n510));
  AND2_X1   g309(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522));
  INV_X1    g321(.A(G43gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(KEYINPUT86), .A3(G50gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n525), .A2(new_n518), .A3(new_n516), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n519), .B1(new_n526), .B2(KEYINPUT87), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n518), .A3(new_n516), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n509), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT13), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT91), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n527), .A2(KEYINPUT17), .A3(new_n530), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n509), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n506), .A2(new_n508), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n531), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n540), .A2(KEYINPUT18), .A3(new_n533), .A4(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n541), .B(new_n531), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n534), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G197gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT11), .B(G169gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT12), .Z(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n540), .A2(new_n542), .ZN(new_n554));
  INV_X1    g353(.A(new_n533), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n547), .A2(new_n552), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n547), .A2(KEYINPUT92), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n536), .A2(new_n560), .A3(new_n543), .A4(new_n546), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n552), .B(KEYINPUT85), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n558), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G127gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n509), .B1(new_n572), .B2(new_n571), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G155gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT94), .B1(G99gat), .B2(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT8), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT94), .A2(G99gat), .A3(G106gat), .ZN(new_n593));
  AND3_X1   g392(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(new_n592), .A2(new_n593), .B1(KEYINPUT7), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT7), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT95), .B(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n595), .B1(new_n599), .B2(new_n594), .ZN(new_n600));
  XOR2_X1   g399(.A(G99gat), .B(G106gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n530), .B2(new_n527), .ZN(new_n603));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n603), .B1(KEYINPUT41), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n538), .A2(new_n539), .A3(new_n602), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n589), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  AOI211_X1 g410(.A(new_n609), .B(new_n588), .C1(new_n605), .C2(new_n606), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n611), .B2(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n566), .B1(new_n587), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n586), .A2(KEYINPUT97), .A3(new_n620), .ZN(new_n623));
  INV_X1    g422(.A(G230gat), .ZN(new_n624));
  INV_X1    g423(.A(G233gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n571), .B1(new_n628), .B2(new_n600), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n602), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n602), .A2(new_n629), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT10), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n602), .A2(new_n633), .A3(new_n571), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n627), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(new_n631), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n635), .B1(new_n627), .B2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G120gat), .B(G148gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT99), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  OR2_X1    g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n622), .A2(new_n623), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n492), .A2(new_n565), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n439), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n650), .A2(KEYINPUT100), .A3(new_n357), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT100), .B1(new_n650), .B2(new_n357), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(G8gat), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n357), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT16), .B(G8gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT101), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n647), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT102), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n656), .B1(new_n651), .B2(new_n652), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n653), .B(new_n660), .C1(new_n661), .C2(KEYINPUT42), .ZN(G1325gat));
  AOI21_X1  g461(.A(G15gat), .B1(new_n647), .B2(new_n404), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n447), .A2(new_n448), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT103), .Z(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n647), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT104), .ZN(G1326gat));
  INV_X1    g467(.A(new_n275), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n647), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT105), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  AND3_X1   g472(.A1(new_n466), .A2(new_n469), .A3(new_n472), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n487), .A2(new_n275), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT84), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n270), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT80), .A4(new_n265), .ZN(new_n678));
  OAI22_X1  g477(.A1(new_n677), .A2(new_n678), .B1(new_n439), .B2(new_n353), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n679), .A2(new_n448), .A3(new_n447), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n676), .A2(new_n491), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n405), .A2(new_n440), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n442), .A2(KEYINPUT35), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n620), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n565), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n586), .A2(new_n644), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n514), .A3(new_n439), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT45), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n620), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n617), .A2(KEYINPUT107), .A3(new_n619), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n693), .ZN(new_n699));
  OAI22_X1  g498(.A1(new_n685), .A2(new_n693), .B1(new_n492), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n689), .B(KEYINPUT106), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n439), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n700), .A2(KEYINPUT108), .A3(new_n701), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n692), .B1(new_n709), .B2(new_n514), .ZN(G1328gat));
  NAND2_X1  g509(.A1(new_n681), .A2(new_n684), .ZN(new_n711));
  AND4_X1   g510(.A1(new_n510), .A2(new_n688), .A3(new_n654), .A4(new_n621), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n687), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT46), .Z(new_n714));
  NOR3_X1   g513(.A1(new_n705), .A2(new_n357), .A3(new_n708), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n510), .ZN(G1329gat));
  INV_X1    g515(.A(new_n404), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(G43gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n690), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n664), .A3(new_n701), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G43gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT47), .B(new_n719), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n704), .A2(new_n707), .A3(new_n664), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n726), .A2(G43gat), .B1(new_n690), .B2(new_n718), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n727), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  OAI21_X1  g528(.A(G50gat), .B1(new_n702), .B2(new_n275), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n686), .A2(G50gat), .A3(new_n275), .A4(new_n689), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n729), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n704), .A2(new_n707), .A3(new_n669), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n729), .A3(G50gat), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n731), .B1(new_n732), .B2(KEYINPUT48), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(G1331gat));
  AND4_X1   g537(.A1(new_n565), .A2(new_n622), .A3(new_n623), .A4(new_n644), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n711), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n439), .B(KEYINPUT111), .Z(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT113), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(G57gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n741), .A2(KEYINPUT114), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n357), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT115), .Z(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n753), .B(new_n754), .Z(G1333gat));
  NOR3_X1   g554(.A1(new_n740), .A2(G71gat), .A3(new_n717), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n747), .A2(new_n664), .A3(new_n749), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(G71gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g558(.A1(new_n750), .A2(new_n669), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g560(.A1(new_n687), .A2(new_n586), .ZN(new_n762));
  AND4_X1   g561(.A1(KEYINPUT51), .A2(new_n711), .A3(new_n621), .A4(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT51), .B1(new_n685), .B2(new_n762), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n645), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(new_n439), .A3(new_n597), .ZN(new_n768));
  INV_X1    g567(.A(new_n762), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n645), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n700), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n706), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n597), .B2(new_n772), .ZN(G1336gat));
  NOR2_X1   g572(.A1(new_n771), .A2(new_n357), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT117), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n771), .B2(new_n357), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(G92gat), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n357), .A2(G92gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n598), .B2(new_n774), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1337gat));
  XOR2_X1   g584(.A(KEYINPUT118), .B(G99gat), .Z(new_n786));
  INV_X1    g585(.A(new_n664), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n771), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n767), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n717), .A2(new_n786), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(G1338gat));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n645), .A2(G106gat), .A3(new_n275), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n763), .B2(new_n765), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n693), .B1(new_n711), .B2(new_n621), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n492), .A2(new_n699), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n669), .B(new_n770), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n792), .B(new_n794), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n794), .A2(KEYINPUT119), .B1(new_n797), .B2(G106gat), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(new_n793), .C1(new_n763), .C2(new_n765), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n803), .B(new_n792), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n794), .A2(KEYINPUT119), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n797), .A2(G106gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT120), .B1(new_n810), .B2(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n802), .B1(new_n807), .B2(new_n811), .ZN(G1339gat));
  NAND4_X1  g611(.A1(new_n622), .A2(new_n565), .A3(new_n623), .A4(new_n645), .ZN(new_n813));
  INV_X1    g612(.A(new_n641), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n636), .A2(new_n633), .ZN(new_n815));
  INV_X1    g614(.A(new_n634), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n626), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n626), .A3(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n635), .A3(KEYINPUT54), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n642), .ZN(new_n823));
  INV_X1    g622(.A(new_n547), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n557), .A2(new_n552), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n554), .A2(new_n555), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n544), .B2(new_n534), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n551), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n819), .A2(new_n821), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n823), .A2(new_n826), .A3(new_n829), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n697), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n826), .A2(new_n644), .A3(new_n829), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n823), .A2(new_n832), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n565), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n834), .B1(new_n837), .B2(new_n697), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n813), .B1(new_n838), .B2(new_n586), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n839), .A2(new_n405), .A3(new_n742), .ZN(new_n840));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n687), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n839), .A2(new_n275), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n654), .A2(new_n717), .A3(new_n706), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n565), .A2(new_n365), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n841), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n840), .B2(new_n644), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n645), .A2(new_n367), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n845), .B2(new_n849), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n844), .B2(new_n587), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n840), .A2(new_n576), .A3(new_n586), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1342gat));
  INV_X1    g652(.A(G134gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n840), .A2(new_n854), .A3(new_n621), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n844), .B2(new_n620), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(KEYINPUT56), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(G1343gat));
  AND2_X1   g658(.A1(new_n839), .A2(new_n742), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n664), .A2(new_n275), .A3(new_n654), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n228), .B1(new_n862), .B2(new_n565), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n664), .A2(new_n706), .A3(new_n654), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n565), .A2(new_n228), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n839), .B2(new_n669), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n275), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n832), .A2(KEYINPUT122), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n830), .A2(new_n871), .A3(new_n831), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n557), .B1(new_n547), .B2(KEYINPUT92), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n563), .B1(new_n874), .B2(new_n561), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n873), .B(new_n823), .C1(new_n875), .C2(new_n558), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n621), .B1(new_n876), .B2(new_n835), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n587), .B1(new_n877), .B2(new_n834), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n869), .B1(new_n878), .B2(new_n813), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n863), .A2(KEYINPUT58), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1344gat));
  OAI21_X1  g684(.A(new_n864), .B1(new_n866), .B2(new_n879), .ZN(new_n886));
  OR3_X1    g685(.A1(new_n886), .A2(KEYINPUT59), .A3(new_n645), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT59), .B1(new_n862), .B2(new_n645), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n229), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n833), .A2(new_n620), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n823), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n835), .B1(new_n891), .B2(new_n565), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n892), .B2(new_n620), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n813), .B1(new_n893), .B2(new_n586), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n669), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n839), .A2(new_n868), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n897), .A2(new_n644), .A3(new_n864), .ZN(new_n898));
  NAND2_X1  g697(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n887), .B(new_n889), .C1(new_n898), .C2(new_n899), .ZN(G1345gat));
  OAI211_X1 g699(.A(new_n586), .B(new_n864), .C1(new_n866), .C2(new_n879), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G155gat), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n587), .A2(G155gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n860), .A2(new_n861), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n902), .A2(new_n904), .A3(KEYINPUT123), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1346gat));
  NOR2_X1   g708(.A1(new_n620), .A2(G162gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n860), .A2(new_n861), .A3(new_n910), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT124), .Z(new_n912));
  OAI21_X1  g711(.A(G162gat), .B1(new_n886), .B2(new_n697), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1347gat));
  OR2_X1    g713(.A1(new_n742), .A2(new_n357), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n717), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n842), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n565), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n357), .A2(new_n439), .ZN(new_n919));
  AND4_X1   g718(.A1(new_n275), .A2(new_n839), .A3(new_n404), .A4(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n319), .A3(new_n687), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n921), .ZN(G1348gat));
  NOR3_X1   g721(.A1(new_n917), .A2(new_n318), .A3(new_n645), .ZN(new_n923));
  AOI21_X1  g722(.A(G176gat), .B1(new_n920), .B2(new_n644), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(G1349gat));
  OAI21_X1  g724(.A(G183gat), .B1(new_n917), .B2(new_n587), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n920), .A2(new_n309), .A3(new_n586), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n920), .A2(new_n281), .A3(new_n698), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n842), .A2(new_n621), .A3(new_n916), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n935));
  AND4_X1   g734(.A1(KEYINPUT125), .A2(new_n934), .A3(new_n935), .A4(G190gat), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n281), .B1(new_n937), .B2(KEYINPUT61), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n934), .A2(new_n938), .B1(KEYINPUT125), .B2(new_n935), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n933), .B1(new_n936), .B2(new_n939), .ZN(G1351gat));
  AND2_X1   g739(.A1(new_n839), .A2(new_n919), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n664), .A2(new_n275), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT126), .B(G197gat), .Z(new_n944));
  NAND3_X1  g743(.A1(new_n943), .A2(new_n687), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n915), .A2(new_n664), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n897), .A2(new_n687), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n948), .B2(new_n944), .ZN(G1352gat));
  NOR2_X1   g748(.A1(new_n645), .A2(G204gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n644), .B(new_n946), .C1(new_n895), .C2(new_n896), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n943), .A2(new_n207), .A3(new_n586), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n586), .B(new_n946), .C1(new_n895), .C2(new_n896), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n943), .B2(new_n698), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n897), .A2(new_n946), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n621), .A2(G218gat), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT127), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n963), .B2(new_n965), .ZN(G1355gat));
endmodule


