//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156, new_n1157, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  AOI22_X1  g039(.A1(new_n462), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n474), .B(new_n481), .C1(G136), .C2(new_n462), .ZN(G162));
  OR2_X1    g057(.A1(new_n475), .A2(G114), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n479), .A2(G126), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n459), .B2(new_n460), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n487), .B1(new_n490), .B2(KEYINPUT68), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n487), .A2(KEYINPUT67), .A3(KEYINPUT68), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(KEYINPUT67), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n486), .A2(new_n491), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT69), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n512));
  OAI221_X1 g087(.A(new_n512), .B1(new_n508), .B2(new_n509), .C1(new_n507), .C2(new_n506), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n511), .A2(new_n513), .B1(G651), .B2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n508), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n505), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n517), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n502), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n503), .B2(new_n504), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n506), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n531), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n502), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT70), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n533), .A2(G43), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT71), .B(G81), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n506), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n540), .B2(KEYINPUT70), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n533), .A2(G53), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT73), .B1(new_n554), .B2(KEYINPUT72), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n555), .B1(KEYINPUT73), .B2(new_n554), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n553), .B(KEYINPUT73), .C1(KEYINPUT72), .C2(new_n554), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n517), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  INV_X1    g137(.A(new_n506), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G91), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n557), .A2(new_n558), .A3(new_n562), .A4(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  NAND2_X1  g141(.A1(new_n511), .A2(new_n513), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n519), .A2(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G303));
  NAND2_X1  g144(.A1(new_n563), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n533), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  AND3_X1   g148(.A1(KEYINPUT74), .A2(G73), .A3(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT74), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n517), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(G48), .B2(new_n533), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n500), .A2(new_n505), .A3(G86), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n500), .A2(new_n505), .A3(KEYINPUT75), .A4(G86), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n517), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n502), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(new_n588), .B2(new_n587), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n563), .A2(G85), .B1(G47), .B2(new_n533), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NOR2_X1   g168(.A1(G301), .A2(new_n593), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n500), .A2(new_n505), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n508), .A2(KEYINPUT78), .ZN(new_n600));
  INV_X1    g175(.A(G54), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n508), .B2(KEYINPUT78), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n517), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n600), .A2(new_n602), .B1(G651), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n597), .A2(new_n598), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n607), .A2(KEYINPUT79), .A3(new_n608), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n594), .B1(new_n613), .B2(new_n593), .ZN(G284));
  AOI21_X1  g189(.A(new_n594), .B1(new_n613), .B2(new_n593), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  XNOR2_X1  g193(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT81), .Z(G148));
  NAND3_X1  g197(.A1(new_n611), .A2(new_n620), .A3(new_n612), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n492), .A2(new_n464), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n462), .A2(G135), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n635), .A2(KEYINPUT83), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(KEYINPUT83), .B2(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n479), .A2(G123), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n634), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT84), .Z(G156));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(G401));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT17), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n667), .B(new_n664), .C1(new_n660), .C2(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n660), .A3(new_n662), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n692), .A2(G23), .ZN(new_n693));
  NAND2_X1  g268(.A1(G288), .A2(KEYINPUT91), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n695));
  NAND4_X1  g270(.A1(new_n570), .A2(new_n695), .A3(new_n571), .A4(new_n572), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n693), .B1(new_n697), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(G22), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT92), .Z(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n692), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n698), .A2(new_n700), .B1(new_n703), .B2(G1971), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G1971), .B2(new_n703), .ZN(new_n705));
  MUX2_X1   g280(.A(G6), .B(G305), .S(G16), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT32), .B(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n698), .A2(new_n700), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n462), .A2(G131), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n479), .A2(G119), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n475), .A2(G107), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n714), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G25), .B(new_n718), .S(G29), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT35), .B(G1991), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT87), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT88), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n719), .B(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G24), .B(G290), .S(G16), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1986), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n723), .B1(new_n725), .B2(KEYINPUT89), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(KEYINPUT89), .B2(new_n725), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n712), .A2(new_n713), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT36), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n692), .A2(G19), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n547), .B2(new_n692), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1341), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n692), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n692), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G33), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT25), .ZN(new_n739));
  NAND2_X1  g314(.A1(G103), .A2(G2104), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G2105), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n475), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n462), .A2(G139), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n475), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n640), .A2(new_n737), .ZN(new_n749));
  INV_X1    g324(.A(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n751));
  AOI21_X1  g326(.A(G29), .B1(new_n750), .B2(KEYINPUT30), .ZN(new_n752));
  OR2_X1    g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  NAND2_X1  g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n751), .A2(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n736), .A2(new_n748), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n462), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n479), .A2(G128), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n475), .A2(G116), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n737), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT93), .B(G2067), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n737), .A2(G27), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT97), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n737), .ZN(new_n770));
  INV_X1    g345(.A(G2078), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G34), .ZN(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n773), .B2(KEYINPUT24), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(KEYINPUT24), .B2(new_n773), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n470), .B2(new_n737), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2084), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n767), .A2(new_n772), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n692), .A2(G20), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT23), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n617), .B2(new_n692), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1956), .ZN(new_n782));
  OR4_X1    g357(.A1(new_n732), .A2(new_n756), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n692), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n613), .B2(new_n692), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1348), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n737), .A2(G35), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G162), .B2(new_n737), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT29), .Z(new_n789));
  INV_X1    g364(.A(G2090), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT96), .B(G1966), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n692), .A2(G21), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G168), .B2(new_n692), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT95), .Z(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n737), .A2(G32), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n462), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n479), .A2(G129), .ZN(new_n801));
  NAND3_X1  g376(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT26), .Z(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n737), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT27), .Z(new_n807));
  AOI22_X1  g382(.A1(new_n807), .A2(G1996), .B1(new_n797), .B2(new_n793), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n746), .A2(new_n747), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT94), .Z(new_n810));
  OAI211_X1 g385(.A(new_n808), .B(new_n810), .C1(G1996), .C2(new_n807), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n783), .A2(new_n786), .A3(new_n798), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n729), .A2(new_n812), .ZN(G150));
  INV_X1    g388(.A(G150), .ZN(G311));
  NAND2_X1  g389(.A1(new_n533), .A2(G55), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n506), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT98), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(new_n502), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT99), .B(G860), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT100), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT37), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n613), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n821), .B(new_n546), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT39), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n822), .ZN(G145));
  XNOR2_X1  g407(.A(G164), .B(new_n761), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n479), .A2(G130), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n475), .A2(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G142), .B2(new_n462), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n833), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n745), .B(new_n804), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n718), .B(new_n629), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n839), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G162), .B(new_n470), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n640), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT101), .B(G37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g424(.A(new_n609), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n617), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n609), .A2(G299), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT41), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(KEYINPUT41), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n623), .A2(new_n829), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n611), .A2(new_n828), .A3(new_n620), .A4(new_n612), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n855), .A2(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n853), .A3(new_n858), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT42), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n855), .A2(new_n856), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n857), .A2(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G303), .B(G305), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n697), .B(G290), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(KEYINPUT102), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(KEYINPUT102), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n862), .A2(new_n867), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G868), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n879));
  INV_X1    g454(.A(new_n821), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(G868), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n593), .B1(new_n874), .B2(new_n876), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT103), .B1(new_n884), .B2(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G295));
  NAND2_X1  g461(.A1(new_n878), .A2(new_n882), .ZN(G331));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n888));
  XNOR2_X1  g463(.A(G301), .B(G286), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n828), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(G301), .B(G168), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n880), .A2(new_n547), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n821), .A2(new_n546), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(KEYINPUT104), .A3(new_n894), .ZN(new_n895));
  OR3_X1    g470(.A1(new_n828), .A2(KEYINPUT104), .A3(new_n889), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n863), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n890), .A2(new_n899), .A3(new_n894), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n828), .A2(KEYINPUT105), .A3(new_n889), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n853), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n873), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n904), .B(new_n873), .C1(new_n863), .C2(new_n897), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n888), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n906), .A2(new_n847), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n855), .A2(new_n856), .A3(new_n901), .A4(new_n900), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n897), .A2(new_n903), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n911), .B1(new_n914), .B2(new_n875), .ZN(new_n915));
  AOI211_X1 g490(.A(KEYINPUT106), .B(new_n873), .C1(new_n912), .C2(new_n913), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n909), .B1(new_n917), .B2(new_n888), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT44), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n905), .B2(new_n908), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n917), .B2(KEYINPUT43), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n923), .ZN(G397));
  XNOR2_X1  g499(.A(KEYINPUT107), .B(G1384), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT45), .B1(new_n496), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n465), .A2(G40), .A3(new_n469), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G2067), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n761), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n931), .B2(new_n805), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT124), .Z(new_n933));
  NOR2_X1   g508(.A1(new_n929), .A2(G1996), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT46), .Z(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT47), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n805), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT108), .Z(new_n939));
  INV_X1    g514(.A(new_n929), .ZN(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n931), .B1(new_n805), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n939), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n718), .B(new_n721), .Z(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(new_n929), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n929), .A2(G1986), .A3(G290), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  XOR2_X1   g522(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n948));
  XNOR2_X1  g523(.A(new_n947), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n937), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n761), .A2(G2067), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n718), .A2(new_n721), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n943), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT123), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n929), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G8), .ZN(new_n958));
  NOR2_X1   g533(.A1(G168), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT51), .B1(new_n960), .B2(KEYINPUT120), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  OAI211_X1 g538(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n483), .A2(new_n485), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n495), .A2(new_n494), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n475), .A2(G138), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n477), .B2(new_n478), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT68), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT4), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT110), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n496), .A2(new_n974), .A3(new_n963), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n927), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(G2084), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n972), .B2(new_n975), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT115), .B1(new_n980), .B2(new_n927), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n971), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n496), .A2(new_n974), .A3(new_n963), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n974), .B1(new_n496), .B2(new_n963), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n928), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n981), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n979), .B1(new_n990), .B2(new_n793), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n960), .B(new_n962), .C1(new_n991), .C2(new_n958), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n793), .ZN(new_n993));
  INV_X1    g568(.A(new_n979), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n959), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n958), .B(new_n962), .C1(new_n991), .C2(G168), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT62), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(G8), .B(new_n961), .C1(new_n995), .C2(G286), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n996), .A4(new_n992), .ZN(new_n1002));
  NAND3_X1  g577(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(G166), .B2(new_n958), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT109), .B(G1971), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n927), .B1(new_n971), .B2(new_n982), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n925), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n928), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n972), .A2(new_n975), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1011), .B1(new_n1014), .B2(new_n790), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1007), .B1(new_n1015), .B2(new_n958), .ZN(new_n1016));
  INV_X1    g591(.A(G1981), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n579), .A2(new_n1017), .A3(new_n582), .A4(new_n583), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n577), .B1(new_n498), .B2(new_n499), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G73), .A2(G543), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT74), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(KEYINPUT74), .A2(G73), .A3(G543), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(G651), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n533), .A2(G48), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n580), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(G1981), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1018), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1027), .B2(G1981), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT112), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1031), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(new_n1018), .A4(new_n1029), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1018), .A3(new_n1029), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT113), .B1(new_n1038), .B2(new_n1033), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1032), .A2(new_n1036), .A3(KEYINPUT113), .A4(new_n1033), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n972), .A2(new_n975), .A3(new_n928), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n958), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1046));
  OAI22_X1  g621(.A1(new_n978), .A2(G2090), .B1(new_n1046), .B2(new_n1008), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(G8), .A3(new_n1006), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n694), .A2(G1976), .A3(new_n696), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1042), .A2(G8), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT52), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1042), .A2(G8), .A3(new_n1049), .A4(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1016), .A2(new_n1045), .A3(new_n1048), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(G2078), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n981), .A2(new_n989), .A3(new_n984), .A4(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1009), .A2(new_n771), .A3(new_n1010), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n978), .A2(new_n735), .B1(new_n1061), .B2(new_n1058), .ZN(new_n1062));
  AOI21_X1  g637(.A(G301), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n999), .A2(new_n1002), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT63), .ZN(new_n1066));
  INV_X1    g641(.A(new_n793), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n927), .B1(new_n1013), .B2(new_n982), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n983), .B1(new_n1068), .B2(new_n988), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1069), .B2(new_n981), .ZN(new_n1070));
  OAI211_X1 g645(.A(G8), .B(G168), .C1(new_n1070), .C2(new_n979), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1071), .B2(new_n1056), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT116), .B(new_n1066), .C1(new_n1071), .C2(new_n1056), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1071), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1045), .A2(new_n1048), .A3(new_n1055), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1047), .A2(G8), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1066), .B1(new_n1078), .B2(new_n1007), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1074), .A2(new_n1075), .A3(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1046), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1956), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n973), .B1(new_n972), .B2(new_n975), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1012), .ZN(new_n1086));
  AND3_X1   g661(.A1(G299), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1083), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1348), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n978), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1043), .A2(new_n930), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n609), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1089), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT118), .B(new_n1090), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1090), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(new_n1095), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1089), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(KEYINPUT61), .A3(new_n1090), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n1093), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1348), .B1(new_n976), .B2(new_n977), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1042), .A2(G2067), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n850), .A3(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1092), .A2(new_n1093), .A3(KEYINPUT60), .A4(new_n609), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(KEYINPUT119), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1046), .A2(new_n941), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT58), .B(G1341), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n1042), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1117), .B1(new_n1121), .B2(new_n547), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n546), .B(new_n1116), .C1(new_n1118), .C2(new_n1120), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1113), .B(new_n1114), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1098), .B(new_n1099), .C1(new_n1107), .C2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1000), .A2(new_n996), .A3(new_n992), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n1128));
  INV_X1    g703(.A(new_n926), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n928), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n927), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1010), .B(new_n1059), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1062), .A2(G301), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1127), .B1(new_n1063), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1060), .A2(G301), .A3(new_n1062), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1062), .A2(new_n1132), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1135), .B(KEYINPUT54), .C1(new_n1136), .C2(G301), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1125), .A2(new_n1126), .A3(new_n1138), .A4(new_n1057), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G288), .A2(G1976), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT114), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1045), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1018), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1045), .A2(new_n1055), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1048), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1143), .A2(new_n1044), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1065), .A2(new_n1081), .A3(new_n1139), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n1148));
  XNOR2_X1  g723(.A(G290), .B(G1986), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n945), .B1(new_n940), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n957), .B1(new_n1151), .B2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g728(.A(G319), .ZN(new_n1155));
  NOR3_X1   g729(.A1(new_n658), .A2(G227), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n690), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g731(.A(new_n1157), .B(KEYINPUT127), .ZN(new_n1158));
  AND3_X1   g732(.A1(new_n1158), .A2(new_n921), .A3(new_n848), .ZN(G308));
  NAND3_X1  g733(.A1(new_n1158), .A2(new_n921), .A3(new_n848), .ZN(G225));
endmodule


