//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G119), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n189), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NOR3_X1   g012(.A1(KEYINPUT64), .A2(KEYINPUT2), .A3(G113), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n200));
  INV_X1    g014(.A(G113), .ZN(new_n201));
  OAI22_X1  g015(.A1(new_n198), .A2(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n188), .B1(new_n196), .B2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT65), .B(G116), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n194), .B1(new_n204), .B2(G119), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n200), .A3(new_n201), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n207), .A2(new_n197), .B1(KEYINPUT2), .B2(G113), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(KEYINPUT66), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT3), .A3(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT77), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n214), .B2(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n212), .A2(KEYINPUT77), .A3(G107), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n216), .A2(new_n217), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n212), .B2(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n212), .A2(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n214), .A2(KEYINPUT78), .A3(G104), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n201), .B1(new_n194), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n196), .B2(new_n230), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n210), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n203), .A2(new_n209), .B1(new_n202), .B2(new_n196), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n214), .A2(KEYINPUT3), .A3(G104), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT3), .B1(new_n214), .B2(G104), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n219), .B(new_n220), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G101), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n240), .A3(G101), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n233), .B1(new_n234), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G110), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n233), .B(new_n244), .C1(new_n234), .C2(new_n242), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT6), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n249), .A3(new_n245), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(G146), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  OAI211_X1 g069(.A(G128), .B(new_n252), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G125), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(G146), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n258), .B(new_n259), .C1(KEYINPUT1), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n256), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G143), .B(G146), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G128), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n262), .B1(new_n257), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n268), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n248), .A2(new_n250), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n268), .A2(KEYINPUT82), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(KEYINPUT82), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n274), .A2(KEYINPUT82), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n268), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n247), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n244), .B(KEYINPUT8), .ZN(new_n282));
  INV_X1    g096(.A(new_n233), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n229), .B1(new_n210), .B2(new_n232), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n287), .B(KEYINPUT83), .Z(new_n288));
  AND3_X1   g102(.A1(new_n272), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n272), .B2(new_n286), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G214), .B1(G237), .B2(G902), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n187), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n292), .ZN(new_n294));
  NOR4_X1   g108(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT84), .A4(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n297));
  INV_X1    g111(.A(G119), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(G128), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n260), .A2(KEYINPUT23), .A3(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(G128), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G110), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT71), .ZN(new_n304));
  XNOR2_X1  g118(.A(G125), .B(G140), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(KEYINPUT16), .ZN(new_n306));
  INV_X1    g120(.A(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G125), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT16), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n254), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n305), .B2(KEYINPUT16), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G146), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT24), .B(G110), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n298), .B2(G128), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n260), .A2(KEYINPUT70), .A3(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n301), .A3(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n304), .B(new_n313), .C1(new_n314), .C2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n257), .A2(G140), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n307), .A2(G125), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n320), .A2(new_n321), .A3(G146), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n311), .B2(G146), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(new_n318), .B2(new_n314), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n324), .A3(new_n314), .ZN(new_n326));
  INV_X1    g140(.A(G110), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n299), .A2(new_n300), .A3(new_n327), .A4(new_n301), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n323), .B(KEYINPUT73), .C1(new_n325), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n318), .A2(new_n314), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT72), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n328), .A3(new_n326), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT73), .B1(new_n334), .B2(new_n323), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n319), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G137), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G902), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n323), .B1(new_n329), .B2(new_n325), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT73), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n330), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n319), .A3(new_n339), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n341), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT25), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n341), .A2(new_n347), .A3(new_n350), .A4(new_n342), .ZN(new_n351));
  INV_X1    g165(.A(G217), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(G234), .B2(new_n342), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(G902), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n341), .A2(new_n347), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n354), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n196), .A2(new_n202), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n196), .A2(new_n202), .A3(new_n188), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT66), .B1(new_n205), .B2(new_n208), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT11), .ZN(new_n366));
  INV_X1    g180(.A(G134), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(G137), .ZN(new_n368));
  INV_X1    g182(.A(G137), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT11), .A3(G134), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(G137), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G131), .ZN(new_n373));
  INV_X1    g187(.A(G131), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n368), .A2(new_n370), .A3(new_n374), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n267), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n367), .A2(G137), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n369), .A2(G134), .ZN(new_n380));
  OAI21_X1  g194(.A(G131), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n256), .A2(new_n375), .A3(new_n381), .A4(new_n261), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n365), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n210), .A2(new_n362), .A3(new_n378), .A4(new_n382), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n361), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n383), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT28), .B1(new_n387), .B2(new_n234), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT68), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n365), .A2(new_n383), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n210), .A2(new_n362), .B1(new_n378), .B2(new_n382), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT28), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT68), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(G237), .A2(G953), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G210), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT27), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT26), .B(G101), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n389), .A2(new_n394), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n267), .B1(new_n375), .B2(new_n373), .ZN(new_n403));
  AND4_X1   g217(.A1(new_n375), .A2(new_n256), .A3(new_n261), .A4(new_n381), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT30), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n378), .B2(new_n382), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n365), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n385), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n409), .B2(new_n400), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT69), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT69), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n386), .A2(new_n388), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n401), .A2(KEYINPUT29), .ZN(new_n416));
  AOI21_X1  g230(.A(G902), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G472), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n389), .A2(new_n394), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n400), .B1(KEYINPUT67), .B2(KEYINPUT31), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n408), .A2(new_n385), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(KEYINPUT67), .A2(KEYINPUT31), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT30), .B1(new_n403), .B2(new_n404), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n378), .A2(new_n406), .A3(new_n382), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n234), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(new_n390), .ZN(new_n428));
  INV_X1    g242(.A(new_n423), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n421), .A3(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n420), .A2(new_n400), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(G472), .A2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT32), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n385), .A2(new_n361), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n393), .B1(new_n392), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n386), .A2(KEYINPUT68), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n400), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n424), .A2(new_n430), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT32), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n432), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n434), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n360), .B1(new_n419), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT9), .B(G234), .ZN(new_n445));
  OAI21_X1  g259(.A(G221), .B1(new_n445), .B2(G902), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT75), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT79), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n256), .A2(new_n261), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n228), .B2(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n256), .A2(new_n261), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n451), .A2(KEYINPUT79), .A3(new_n221), .A4(new_n227), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n228), .A2(new_n449), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n376), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT12), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n457), .A3(new_n376), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT10), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n450), .A2(new_n452), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n376), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n229), .A2(KEYINPUT10), .A3(new_n451), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n239), .A2(new_n377), .A3(new_n241), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n456), .A2(new_n458), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n269), .A2(G227), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT76), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G140), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT80), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n450), .A2(new_n459), .A3(new_n452), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n463), .A2(new_n462), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n376), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n469), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n464), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n471), .B1(new_n470), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n342), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G469), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  AND4_X1   g295(.A1(new_n458), .A2(new_n456), .A3(new_n464), .A4(new_n475), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n475), .B1(new_n474), .B2(new_n464), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n481), .B(new_n342), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT81), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n463), .A2(new_n462), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n461), .B1(new_n487), .B2(new_n460), .ZN(new_n488));
  INV_X1    g302(.A(new_n464), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n469), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n456), .A2(new_n458), .A3(new_n464), .A4(new_n475), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT81), .A3(new_n481), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n447), .B1(new_n480), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G237), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n269), .A3(G214), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n251), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n395), .A2(G143), .A3(G214), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT17), .A3(G131), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n310), .A2(new_n312), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(G131), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n374), .A3(new_n499), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n507), .A2(KEYINPUT17), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT89), .A4(new_n501), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AND4_X1   g324(.A1(G143), .A2(new_n496), .A3(new_n269), .A4(G214), .ZN(new_n511));
  AOI21_X1  g325(.A(G143), .B1(new_n395), .B2(G214), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(KEYINPUT18), .A2(G131), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n305), .A2(new_n254), .ZN(new_n515));
  OAI21_X1  g329(.A(G146), .B1(new_n320), .B2(new_n321), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n518));
  INV_X1    g332(.A(new_n514), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n500), .B2(new_n519), .ZN(new_n520));
  AOI211_X1 g334(.A(KEYINPUT85), .B(new_n514), .C1(new_n498), .C2(new_n499), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n517), .B(KEYINPUT86), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G113), .B(G122), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(new_n212), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n510), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n510), .B2(new_n526), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n342), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G475), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT19), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT87), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n305), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n538), .B(new_n254), .C1(new_n305), .C2(new_n537), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n507), .A2(new_n312), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n524), .B2(new_n525), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT88), .B1(new_n541), .B2(new_n528), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n507), .A2(new_n539), .A3(new_n312), .ZN(new_n543));
  INV_X1    g357(.A(new_n525), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n519), .B1(new_n511), .B2(new_n512), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT85), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n500), .A2(new_n518), .A3(new_n519), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT86), .B1(new_n548), .B2(new_n517), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n543), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT88), .ZN(new_n551));
  INV_X1    g365(.A(new_n528), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n542), .A2(new_n553), .A3(new_n529), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT20), .ZN(new_n555));
  NOR2_X1   g369(.A1(G475), .A2(G902), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n533), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G478), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n445), .A2(new_n352), .A3(G953), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT92), .Z(new_n563));
  INV_X1    g377(.A(G122), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G116), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT90), .B1(new_n204), .B2(G122), .ZN(new_n566));
  AND4_X1   g380(.A1(KEYINPUT90), .A2(new_n190), .A3(new_n192), .A4(G122), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n214), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n251), .A2(G128), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n260), .A2(G143), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n367), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n570), .A3(G134), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT14), .B1(new_n566), .B2(new_n567), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n190), .A2(new_n192), .A3(G122), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n204), .A2(KEYINPUT90), .A3(G122), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT14), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n576), .A2(new_n565), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n575), .B1(G107), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(G134), .A3(new_n570), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n572), .A3(new_n573), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n585), .A2(G134), .A3(new_n569), .A4(new_n570), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G107), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n591), .B2(new_n568), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n563), .B1(new_n584), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n583), .A2(G107), .ZN(new_n594));
  INV_X1    g408(.A(new_n575), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n563), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n591), .A2(new_n568), .ZN(new_n598));
  INV_X1    g412(.A(new_n589), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n593), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(KEYINPUT93), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n604), .B(G902), .C1(new_n593), .C2(new_n601), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n561), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n605), .A2(new_n561), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(G234), .A2(G237), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n609), .A2(G952), .A3(new_n269), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n609), .A2(G902), .A3(G953), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT21), .B(G898), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n559), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n296), .A2(new_n444), .A3(new_n495), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n431), .B2(new_n433), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n431), .B2(G902), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n617), .B(G472), .C1(new_n431), .C2(G902), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n360), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n495), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n625), .B(KEYINPUT95), .Z(new_n626));
  INV_X1    g440(.A(new_n613), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n291), .A2(new_n627), .A3(new_n292), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n597), .B1(new_n596), .B2(new_n600), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n584), .A2(new_n563), .A3(new_n592), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(KEYINPUT96), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n593), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g451(.A(KEYINPUT97), .B(new_n563), .C1(new_n584), .C2(new_n592), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT33), .A4(new_n601), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n560), .A2(G902), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n634), .A2(new_n635), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n602), .A2(G478), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n559), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n628), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n626), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n554), .A2(new_n556), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT20), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n650), .A2(new_n651), .B1(G475), .B2(new_n532), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n608), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n628), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n626), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  NAND2_X1  g471(.A1(new_n336), .A2(KEYINPUT98), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n340), .A2(KEYINPUT36), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n346), .A2(new_n660), .A3(new_n319), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n659), .B1(new_n658), .B2(new_n661), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n355), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n354), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n354), .A2(new_n664), .A3(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n296), .A2(new_n614), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n623), .A2(new_n495), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT37), .B(G110), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AOI22_X1  g488(.A1(new_n419), .A2(new_n443), .B1(new_n667), .B2(new_n668), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n650), .A2(new_n651), .ZN(new_n676));
  INV_X1    g490(.A(new_n610), .ZN(new_n677));
  INV_X1    g491(.A(new_n611), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n677), .B1(new_n678), .B2(G900), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT100), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n608), .A2(new_n676), .A3(new_n533), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n291), .A2(new_n292), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n675), .A2(new_n495), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(new_n680), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n495), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n291), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n428), .A2(new_n400), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n384), .A2(new_n385), .A3(new_n400), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n342), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n443), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n443), .A2(KEYINPUT102), .A3(new_n695), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n691), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n668), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT99), .B1(new_n354), .B2(new_n664), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n559), .A2(new_n608), .A3(new_n292), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT103), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n559), .A2(new_n608), .A3(new_n292), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n706), .B1(new_n669), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT40), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n495), .A2(new_n710), .A3(new_n687), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n689), .A2(new_n700), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND3_X1  g527(.A1(new_n559), .A2(new_n643), .A3(new_n681), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n683), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n675), .A2(new_n495), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  INV_X1    g531(.A(new_n447), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n492), .A2(new_n481), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n494), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n494), .A2(KEYINPUT104), .A3(new_n718), .A4(new_n719), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n444), .A3(new_n645), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n654), .A2(new_n722), .A3(new_n444), .A4(new_n723), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NOR2_X1   g542(.A1(new_n720), .A2(new_n683), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n675), .A3(new_n614), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n400), .B1(new_n386), .B2(new_n388), .ZN(new_n733));
  AOI211_X1 g547(.A(new_n732), .B(new_n433), .C1(new_n439), .C2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n429), .B1(new_n428), .B2(new_n421), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n385), .A2(new_n408), .A3(new_n421), .A4(new_n429), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT105), .B1(new_n737), .B2(new_n432), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  AOI21_X1  g554(.A(G902), .B1(new_n438), .B2(new_n439), .ZN(new_n741));
  INV_X1    g555(.A(G472), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT106), .B(G472), .C1(new_n431), .C2(G902), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n739), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n559), .A2(new_n291), .A3(new_n608), .A4(new_n292), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n746), .A3(new_n624), .A4(new_n627), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n722), .A2(new_n723), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n564), .ZN(G24));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n714), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n559), .A2(new_n643), .A3(KEYINPUT107), .A4(new_n681), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n739), .A2(new_n743), .A3(new_n744), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n703), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n729), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(new_n417), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n411), .B2(KEYINPUT69), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n742), .B1(new_n760), .B2(new_n414), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(KEYINPUT111), .B2(new_n443), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n443), .A2(KEYINPUT111), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n360), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n470), .B2(new_n476), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT108), .B1(new_n465), .B2(new_n469), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n342), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n768), .A2(G469), .B1(new_n486), .B2(new_n493), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n447), .A2(new_n294), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n289), .B2(new_n290), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT109), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n773));
  INV_X1    g587(.A(new_n771), .ZN(new_n774));
  INV_X1    g588(.A(new_n767), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n474), .A2(new_n464), .A3(new_n475), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n465), .B2(new_n469), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n775), .B1(new_n777), .B2(new_n765), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n481), .B1(new_n778), .B2(new_n342), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n484), .A2(new_n485), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT81), .B1(new_n492), .B2(new_n481), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n773), .B(new_n774), .C1(new_n779), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n772), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n764), .A2(new_n784), .A3(KEYINPUT42), .A4(new_n754), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n784), .A2(new_n786), .A3(new_n754), .A4(new_n444), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n434), .A2(new_n442), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n624), .B1(new_n790), .B2(new_n761), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n772), .B2(new_n783), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n786), .B1(new_n792), .B2(new_n754), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n785), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G131), .ZN(G33));
  INV_X1    g609(.A(new_n682), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  NOR2_X1   g612(.A1(new_n766), .A2(new_n767), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n481), .B1(new_n799), .B2(KEYINPUT45), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n477), .B2(new_n478), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n800), .A2(new_n802), .B1(G469), .B2(G902), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT112), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n782), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n802), .B(G469), .C1(new_n801), .C2(new_n778), .ZN(new_n806));
  NAND2_X1  g620(.A1(G469), .A2(G902), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT46), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(new_n805), .A3(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(new_n718), .A3(new_n687), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n652), .A2(new_n643), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT43), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT43), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n652), .A2(new_n817), .A3(new_n643), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n622), .A2(new_n669), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n814), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n292), .B1(new_n289), .B2(new_n290), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n819), .A2(new_n820), .A3(new_n814), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n813), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G137), .ZN(G39));
  INV_X1    g642(.A(new_n714), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n624), .A2(new_n822), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n443), .A4(new_n419), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n812), .A2(KEYINPUT47), .A3(new_n718), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT47), .B1(new_n812), .B2(new_n718), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  NAND3_X1  g651(.A1(new_n816), .A2(new_n610), .A3(new_n818), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n360), .A3(new_n755), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n729), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT120), .Z(new_n841));
  NOR3_X1   g655(.A1(new_n838), .A2(new_n720), .A3(new_n822), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n764), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT48), .ZN(new_n844));
  INV_X1    g658(.A(G952), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n720), .A2(new_n822), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n360), .A2(new_n677), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n698), .A2(new_n846), .A3(new_n699), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n644), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n845), .B(G953), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n841), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n691), .A2(new_n294), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n720), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n839), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT50), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n839), .A2(KEYINPUT50), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n842), .A2(KEYINPUT117), .A3(new_n756), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n846), .A2(new_n610), .A3(new_n816), .A4(new_n818), .ZN(new_n861));
  INV_X1    g675(.A(new_n756), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n559), .A2(new_n643), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n859), .A2(new_n863), .B1(new_n848), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n858), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n859), .A2(new_n863), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n848), .A2(new_n864), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n868), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT119), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n869), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n865), .A2(new_n866), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n858), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n834), .A2(new_n835), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n494), .A2(new_n719), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n718), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n839), .A2(new_n823), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT115), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n878), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n851), .B1(new_n877), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n883), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n880), .A2(new_n718), .ZN(new_n887));
  INV_X1    g701(.A(new_n835), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n833), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n858), .A2(new_n865), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n878), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n768), .A2(G469), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n494), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n665), .A2(new_n447), .A3(new_n680), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n746), .A2(new_n696), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n716), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n901), .A2(KEYINPUT52), .A3(new_n685), .A4(new_n757), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n745), .A2(new_n669), .A3(new_n752), .A4(new_n753), .ZN(new_n904));
  INV_X1    g718(.A(new_n729), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n685), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n716), .A2(new_n900), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT114), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT114), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n902), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n615), .B(new_n730), .C1(new_n671), .C2(new_n670), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n653), .A2(new_n644), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n296), .A2(new_n627), .A3(new_n915), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n625), .A2(new_n916), .B1(new_n747), .B2(new_n748), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n727), .A2(new_n724), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n784), .A2(new_n756), .A3(new_n754), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n822), .A2(new_n559), .A3(new_n608), .A4(new_n680), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n675), .A2(new_n921), .A3(new_n495), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n797), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n794), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT53), .B1(new_n913), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n909), .A2(new_n794), .A3(new_n919), .A4(new_n923), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT53), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT54), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n913), .A2(KEYINPUT53), .A3(new_n924), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n927), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  OAI22_X1  g748(.A1(new_n896), .A2(new_n934), .B1(G952), .B2(G953), .ZN(new_n935));
  INV_X1    g749(.A(new_n815), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n624), .A2(new_n770), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n691), .B(new_n936), .C1(KEYINPUT113), .C2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(KEYINPUT113), .B2(new_n937), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n880), .B(KEYINPUT49), .Z(new_n940));
  NAND4_X1  g754(.A1(new_n939), .A2(new_n698), .A3(new_n699), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n935), .A2(new_n941), .ZN(G75));
  NAND2_X1  g756(.A1(new_n930), .A2(new_n932), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(G902), .A3(new_n288), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT56), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n248), .A2(new_n250), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n271), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n944), .B2(new_n945), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n845), .A2(G953), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT121), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n949), .A2(new_n950), .A3(new_n953), .ZN(G51));
  XOR2_X1   g768(.A(new_n807), .B(KEYINPUT57), .Z(new_n955));
  AND3_X1   g769(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n490), .A2(new_n491), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n943), .A2(G902), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n961), .A2(new_n806), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n952), .B1(new_n960), .B2(new_n962), .ZN(G54));
  NAND2_X1  g777(.A1(KEYINPUT58), .A2(G475), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n554), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n554), .ZN(new_n966));
  INV_X1    g780(.A(new_n964), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n943), .A2(G902), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n952), .B1(new_n965), .B2(new_n968), .ZN(G60));
  AND3_X1   g783(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(new_n970));
  NAND2_X1  g784(.A1(G478), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT59), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n970), .B(new_n972), .C1(new_n956), .C2(new_n957), .ZN(new_n973));
  INV_X1    g787(.A(new_n953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n934), .B2(new_n972), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G63));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n662), .A2(new_n663), .ZN(new_n979));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT60), .Z(new_n981));
  NAND3_X1  g795(.A1(new_n943), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n974), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n943), .A2(new_n981), .B1(new_n347), .B2(new_n341), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n978), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n943), .A2(new_n981), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n341), .A2(new_n347), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n974), .A4(new_n982), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n985), .A2(new_n989), .ZN(G66));
  INV_X1    g804(.A(G224), .ZN(new_n991));
  OAI21_X1  g805(.A(G953), .B1(new_n612), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n919), .B2(G953), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n946), .B1(G898), .B2(new_n269), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT123), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n993), .B(new_n995), .ZN(G69));
  NAND2_X1  g810(.A1(G900), .A2(G953), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n405), .A2(new_n407), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n538), .B1(new_n305), .B2(new_n537), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n716), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n906), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n797), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(new_n813), .B2(new_n826), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n813), .A2(new_n746), .A3(new_n764), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1004), .A2(new_n794), .A3(new_n836), .A4(new_n1005), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n997), .B(new_n1000), .C1(new_n1006), .C2(G953), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n689), .A2(new_n700), .A3(new_n709), .A4(new_n711), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n757), .A2(new_n685), .A3(new_n716), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1002), .A2(KEYINPUT62), .A3(new_n712), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n444), .A2(new_n823), .A3(new_n915), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1014), .A2(new_n688), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n813), .B2(new_n826), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1013), .A2(new_n836), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT125), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1013), .A2(new_n836), .A3(KEYINPUT125), .A4(new_n1016), .ZN(new_n1020));
  AOI21_X1  g834(.A(G953), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1000), .B(KEYINPUT124), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1007), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(G72));
  NAND3_X1  g839(.A1(new_n1019), .A2(new_n919), .A3(new_n1020), .ZN(new_n1026));
  XNOR2_X1  g840(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n692), .ZN(new_n1031));
  INV_X1    g845(.A(new_n919), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1029), .B1(new_n1006), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n409), .A2(new_n401), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n952), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1034), .ZN(new_n1036));
  INV_X1    g850(.A(new_n692), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1036), .A2(new_n1037), .A3(new_n1029), .ZN(new_n1038));
  INV_X1    g852(.A(new_n912), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n911), .B1(new_n902), .B2(new_n908), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n794), .A2(new_n919), .A3(new_n923), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n927), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n928), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1038), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1045), .A2(KEYINPUT127), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT127), .ZN(new_n1047));
  AOI211_X1 g861(.A(new_n1047), .B(new_n1038), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1048));
  OAI211_X1 g862(.A(new_n1031), .B(new_n1035), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1049), .ZN(G57));
endmodule


