//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT13), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(new_n190), .ZN(new_n195));
  OAI21_X1  g009(.A(G134), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(new_n193), .A3(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT77), .B(G107), .ZN(new_n199));
  XNOR2_X1  g013(.A(G116), .B(G122), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n200), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n196), .B(new_n198), .C1(new_n201), .C2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT14), .A3(G122), .ZN(new_n206));
  INV_X1    g020(.A(new_n200), .ZN(new_n207));
  OAI211_X1 g021(.A(G107), .B(new_n206), .C1(new_n207), .C2(KEYINPUT14), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n189), .A2(new_n193), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n198), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n211), .A3(new_n202), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n204), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT9), .B(G234), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(G217), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n187), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(KEYINPUT91), .A3(new_n218), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n214), .A2(KEYINPUT90), .A3(new_n219), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n213), .B2(new_n218), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  INV_X1    g042(.A(G478), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n227), .B(new_n228), .C1(KEYINPUT15), .C2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(KEYINPUT15), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n220), .A2(new_n221), .B1(new_n223), .B2(new_n225), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G902), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G125), .B(G140), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT16), .ZN(new_n237));
  INV_X1    g051(.A(G140), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G125), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n239), .A2(KEYINPUT16), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(G146), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(G146), .B1(new_n237), .B2(new_n240), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n217), .A3(G214), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n188), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n245), .A2(new_n217), .A3(G143), .A4(G214), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT17), .A3(G131), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(G131), .ZN(new_n251));
  INV_X1    g065(.A(G131), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n252), .A3(new_n248), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n244), .B(new_n250), .C1(KEYINPUT17), .C2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G113), .B(G122), .ZN(new_n256));
  INV_X1    g070(.A(G104), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G125), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G140), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n239), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(G146), .B1(new_n261), .B2(KEYINPUT74), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(KEYINPUT74), .B2(new_n261), .ZN(new_n263));
  INV_X1    g077(.A(G146), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n236), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT86), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n247), .A2(new_n266), .A3(new_n248), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT18), .A2(G131), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n265), .A2(new_n269), .A3(KEYINPUT87), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT87), .B1(new_n265), .B2(new_n269), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n255), .B(new_n258), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n269), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT87), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n265), .A2(new_n269), .A3(KEYINPUT87), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT74), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT88), .B1(new_n236), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT19), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT88), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT74), .B1(new_n280), .B2(new_n279), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n278), .A2(new_n279), .B1(new_n236), .B2(new_n281), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n282), .A2(G146), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n242), .B1(new_n251), .B2(new_n253), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n275), .A2(new_n276), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n272), .B1(new_n285), .B2(new_n258), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G475), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n228), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT20), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT20), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n286), .A2(new_n291), .A3(new_n288), .A4(new_n228), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(G234), .A2(G237), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(G952), .A3(new_n217), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n295), .B(KEYINPUT92), .Z(new_n296));
  AND3_X1   g110(.A1(new_n294), .A2(G902), .A3(G953), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT21), .B(G898), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n255), .B1(new_n270), .B2(new_n271), .ZN(new_n302));
  INV_X1    g116(.A(new_n258), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT89), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n304), .A2(new_n305), .A3(new_n272), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n228), .B1(new_n304), .B2(new_n305), .ZN(new_n307));
  OAI21_X1  g121(.A(G475), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n235), .A2(new_n293), .A3(new_n301), .A4(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  OAI21_X1  g125(.A(G210), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT5), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(G116), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT69), .B1(new_n205), .B2(G119), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT69), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n314), .A3(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n205), .A2(G119), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(G113), .B(new_n315), .C1(new_n320), .C2(new_n313), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT2), .B(G113), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n257), .A2(G107), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G101), .B1(new_n257), .B2(G107), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(KEYINPUT76), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AND4_X1   g148(.A1(KEYINPUT78), .A2(new_n334), .A3(new_n199), .A4(G104), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n257), .B1(new_n331), .B2(new_n333), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT78), .B1(new_n336), .B2(new_n199), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n329), .B(new_n330), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n199), .A2(G104), .ZN(new_n339));
  OAI21_X1  g153(.A(G101), .B1(new_n339), .B2(new_n326), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n338), .A2(KEYINPUT80), .A3(new_n340), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n325), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  INV_X1    g161(.A(G101), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n334), .A2(new_n199), .A3(G104), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n336), .A2(KEYINPUT78), .A3(new_n199), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n328), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n257), .A2(G107), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n338), .A2(KEYINPUT4), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT79), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n353), .B2(new_n330), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n329), .B(new_n354), .C1(new_n335), .C2(new_n337), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G101), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n320), .A2(new_n322), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n324), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT70), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n358), .A3(G101), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n346), .B(new_n347), .C1(new_n365), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n347), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n357), .B2(new_n363), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(new_n345), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(KEYINPUT6), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n264), .A2(G143), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n188), .A2(G146), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT1), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G128), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT65), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n188), .A2(KEYINPUT65), .A3(G146), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n384), .A2(new_n385), .B1(G143), .B2(new_n264), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n192), .B1(new_n378), .B2(KEYINPUT1), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n259), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT0), .A2(G128), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NOR3_X1   g207(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n378), .A2(new_n379), .ZN(new_n396));
  OAI22_X1  g210(.A1(new_n386), .A2(new_n395), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G125), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n377), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n377), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G224), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n402), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n407), .B(new_n373), .C1(new_n374), .C2(new_n345), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n376), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n390), .A2(new_n398), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT85), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n411), .A2(KEYINPUT7), .A3(new_n405), .A4(new_n400), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(KEYINPUT7), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n399), .B2(new_n401), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n338), .A2(new_n340), .ZN(new_n416));
  INV_X1    g230(.A(new_n325), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n346), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n347), .B(KEYINPUT8), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n420), .B2(new_n371), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n312), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n409), .A2(new_n421), .A3(new_n312), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n310), .B(new_n311), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G221), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n426), .B1(new_n216), .B2(new_n228), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G137), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT11), .B1(new_n429), .B2(G134), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n429), .B2(G134), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(KEYINPUT11), .A3(G134), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n433), .A2(new_n429), .A3(KEYINPUT11), .A4(G134), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G131), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n438), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n430), .B(KEYINPUT67), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n252), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n338), .A2(KEYINPUT80), .A3(new_n340), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT80), .B1(new_n338), .B2(new_n340), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n447), .A2(new_n448), .A3(new_n388), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n382), .B1(new_n380), .B2(new_n387), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n416), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n446), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT12), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n343), .A2(new_n389), .A3(new_n344), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n416), .A2(new_n450), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n455), .A3(new_n446), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT10), .ZN(new_n463));
  AND4_X1   g277(.A1(new_n463), .A2(new_n338), .A3(new_n340), .A4(new_n450), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n389), .B1(new_n343), .B2(new_n344), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n465), .B1(new_n466), .B2(new_n463), .ZN(new_n467));
  INV_X1    g281(.A(new_n397), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n369), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n364), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n443), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G140), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n217), .A2(G227), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n462), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n388), .B1(new_n447), .B2(new_n448), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n464), .B1(new_n479), .B2(KEYINPUT10), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n469), .B1(new_n357), .B2(new_n363), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n480), .A2(new_n443), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n472), .B1(new_n467), .B2(new_n471), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n476), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT83), .B(G469), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n228), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n477), .B1(new_n462), .B2(new_n473), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n443), .B1(new_n480), .B2(new_n481), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n490), .A2(new_n473), .A3(new_n477), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT82), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n455), .B1(new_n460), .B2(new_n446), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n456), .B(new_n445), .C1(new_n458), .C2(new_n459), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n476), .B1(new_n495), .B2(new_n482), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n473), .A3(new_n477), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G469), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n488), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n314), .B2(G128), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n505), .C1(G119), .C2(new_n192), .ZN(new_n506));
  XNOR2_X1  g320(.A(G119), .B(G128), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  AOI22_X1  g322(.A1(new_n506), .A2(G110), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n242), .B2(new_n243), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n506), .A2(G110), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n263), .A2(new_n511), .A3(new_n241), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT22), .B(G137), .ZN(new_n514));
  INV_X1    g328(.A(G234), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n426), .A2(new_n515), .A3(G953), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n514), .B(new_n516), .Z(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(new_n512), .A3(new_n517), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n228), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n523), .A2(KEYINPUT75), .ZN(new_n524));
  OAI21_X1  g338(.A(G217), .B1(new_n515), .B2(G902), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT73), .ZN(new_n526));
  INV_X1    g340(.A(new_n523), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT75), .B1(new_n521), .B2(new_n522), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n524), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n519), .A2(new_n520), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n515), .B2(G217), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n397), .B1(new_n439), .B2(new_n442), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n197), .A2(G137), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n429), .A2(G134), .ZN(new_n537));
  OAI21_X1  g351(.A(G131), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n442), .A2(new_n388), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(KEYINPUT30), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n442), .A2(new_n388), .A3(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n468), .A2(KEYINPUT66), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT66), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n439), .A2(new_n442), .B1(new_n397), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n540), .B(new_n368), .C1(new_n545), .C2(KEYINPUT30), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n367), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n535), .A2(new_n548), .A3(new_n539), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n245), .A2(new_n217), .A3(G210), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n550), .B(KEYINPUT27), .Z(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT26), .B(G101), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(KEYINPUT71), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n546), .A2(KEYINPUT31), .A3(new_n549), .A4(new_n554), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n549), .A2(KEYINPUT28), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT28), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n541), .A2(new_n534), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(new_n548), .ZN(new_n562));
  OAI22_X1  g376(.A1(new_n559), .A2(new_n562), .B1(new_n548), .B2(new_n545), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n557), .A2(new_n558), .B1(new_n563), .B2(new_n553), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n368), .B1(new_n541), .B2(new_n534), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n559), .B2(new_n562), .ZN(new_n569));
  INV_X1    g383(.A(new_n553), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT29), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n228), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n570), .B1(new_n561), .B2(new_n548), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n563), .A2(new_n570), .B1(new_n546), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n573), .B1(new_n575), .B2(KEYINPUT29), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n567), .A2(KEYINPUT32), .B1(new_n576), .B2(G472), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n564), .B2(new_n566), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n533), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n425), .A2(new_n428), .A3(new_n502), .A4(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT93), .B(G101), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(G3));
  INV_X1    g397(.A(new_n533), .ZN(new_n584));
  OAI21_X1  g398(.A(G472), .B1(new_n564), .B2(G902), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n557), .A2(new_n558), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n563), .A2(new_n553), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n565), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n502), .A2(new_n428), .A3(new_n584), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n219), .A2(KEYINPUT95), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT33), .B1(new_n213), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n213), .B2(new_n593), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(new_n227), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n229), .A2(G902), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n227), .A2(new_n228), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT96), .B(G478), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n597), .A2(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n300), .B(new_n601), .C1(new_n293), .C2(new_n308), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n409), .A2(new_n421), .A3(new_n603), .A4(new_n312), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n311), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n423), .A2(new_n422), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n606), .B2(KEYINPUT94), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n592), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  NAND2_X1  g424(.A1(new_n293), .A2(new_n308), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n611), .A2(new_n300), .A3(new_n235), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n592), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G107), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NAND2_X1  g430(.A1(new_n409), .A2(new_n421), .ZN(new_n617));
  INV_X1    g431(.A(new_n312), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n409), .A2(new_n421), .A3(new_n312), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n518), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n513), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n531), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n529), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n309), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n621), .A2(new_n311), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n428), .A3(new_n502), .A4(new_n590), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  NAND3_X1  g446(.A1(new_n588), .A2(KEYINPUT32), .A3(new_n565), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n563), .A2(new_n570), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n546), .A2(new_n574), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT29), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G472), .B1(new_n636), .B2(new_n572), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n633), .A2(new_n579), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n293), .A2(new_n308), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n234), .ZN(new_n640));
  INV_X1    g454(.A(new_n296), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(new_n297), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n619), .A2(KEYINPUT94), .A3(new_n620), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n604), .A2(new_n311), .ZN(new_n646));
  AND4_X1   g460(.A1(new_n638), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n502), .A2(new_n428), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n625), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XOR2_X1   g464(.A(new_n643), .B(KEYINPUT39), .Z(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n639), .A2(new_n235), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n311), .A3(new_n626), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(G472), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n546), .A2(new_n549), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n570), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n574), .B2(new_n568), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n633), .B(new_n579), .C1(new_n659), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n656), .A2(new_n657), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n658), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n606), .B(KEYINPUT38), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n653), .A2(new_n654), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  INV_X1    g484(.A(new_n601), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n611), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n643), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n638), .A2(new_n645), .A3(new_n646), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n648), .A2(new_n625), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  AOI21_X1  g490(.A(G902), .B1(new_n478), .B2(new_n484), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n501), .ZN(new_n678));
  AOI211_X1 g492(.A(G902), .B(new_n486), .C1(new_n478), .C2(new_n484), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n678), .A2(new_n679), .A3(new_n427), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n607), .A2(new_n580), .A3(new_n602), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND4_X1  g497(.A1(new_n607), .A2(new_n580), .A3(new_n612), .A4(new_n680), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  NAND2_X1  g499(.A1(new_n627), .A2(new_n638), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n645), .A2(new_n646), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n488), .B(new_n428), .C1(new_n501), .C2(new_n677), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT99), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT99), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n680), .A2(new_n690), .A3(new_n645), .A4(new_n646), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n686), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT100), .B(G119), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G21));
  NAND2_X1  g508(.A1(new_n569), .A2(new_n553), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n586), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n565), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n585), .A2(new_n697), .A3(new_n584), .A4(new_n301), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n688), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n607), .A3(new_n655), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT101), .B(G122), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G24));
  AND2_X1   g516(.A1(new_n585), .A2(new_n697), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n673), .A2(new_n703), .A3(new_n625), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n690), .B1(new_n607), .B2(new_n680), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n687), .A2(KEYINPUT99), .A3(new_n688), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n496), .A2(new_n498), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n501), .B1(new_n710), .B2(new_n228), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n711), .B2(new_n679), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n489), .A2(new_n491), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n713), .B2(G902), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(KEYINPUT102), .A3(new_n488), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n311), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n427), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n619), .A2(new_n620), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n716), .A2(new_n720), .A3(new_n580), .A4(new_n673), .ZN(new_n721));
  XOR2_X1   g535(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT104), .B1(new_n567), .B2(KEYINPUT32), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT32), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n589), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n577), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n584), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n719), .B1(new_n712), .B2(new_n715), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n731), .A3(KEYINPUT42), .A4(new_n673), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n723), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NAND3_X1  g548(.A1(new_n731), .A2(new_n580), .A3(new_n644), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  NAND2_X1  g550(.A1(new_n651), .A2(new_n428), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n501), .A2(new_n228), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n492), .A2(new_n499), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n501), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n744), .A2(KEYINPUT105), .B1(KEYINPUT45), .B2(new_n713), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n492), .B2(new_n499), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(new_n747), .B2(new_n501), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT106), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n489), .A2(new_n491), .A3(KEYINPUT82), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n497), .B1(new_n496), .B2(new_n498), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n743), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT105), .A3(G469), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n713), .A2(KEYINPUT45), .ZN(new_n754));
  AND4_X1   g568(.A1(KEYINPUT106), .A2(new_n753), .A3(new_n748), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n741), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n488), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n748), .A3(new_n754), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n753), .A2(new_n748), .A3(KEYINPUT106), .A4(new_n754), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n739), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT46), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n738), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n739), .B1(new_n760), .B2(new_n761), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n756), .B(new_n488), .C1(new_n768), .C2(KEYINPUT46), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(KEYINPUT107), .A3(new_n738), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n639), .A2(new_n671), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n625), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n590), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(KEYINPUT44), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(KEYINPUT44), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n619), .A2(new_n311), .A3(new_n620), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n767), .A2(new_n770), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT108), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  OAI21_X1  g596(.A(new_n428), .B1(new_n757), .B2(new_n764), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n769), .A2(new_n785), .A3(new_n428), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n673), .A2(new_n533), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n787), .A2(new_n638), .A3(new_n778), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  AND4_X1   g604(.A1(new_n584), .A2(new_n773), .A3(new_n641), .A4(new_n703), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n717), .A3(new_n667), .A4(new_n680), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n678), .A2(new_n679), .A3(new_n296), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n720), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n533), .A3(new_n664), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n639), .A3(new_n601), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n773), .A2(new_n720), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n703), .A2(new_n625), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n801), .A3(KEYINPUT116), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n798), .A2(new_n801), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AND4_X1   g619(.A1(KEYINPUT51), .A2(new_n794), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n678), .A2(new_n679), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n427), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n784), .B2(new_n786), .ZN(new_n810));
  INV_X1    g624(.A(new_n778), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n791), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(G952), .ZN(new_n814));
  INV_X1    g628(.A(new_n672), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n814), .B(G953), .C1(new_n797), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n799), .A2(new_n729), .ZN(new_n817));
  AND2_X1   g631(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n816), .B(new_n819), .C1(new_n817), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n689), .A2(new_n691), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n791), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n794), .A2(new_n801), .A3(new_n798), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n808), .B(KEYINPUT115), .Z(new_n827));
  OAI21_X1  g641(.A(new_n763), .B1(new_n749), .B2(new_n755), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n740), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n679), .B1(new_n762), .B2(new_n741), .ZN(new_n830));
  AOI211_X1 g644(.A(KEYINPUT47), .B(new_n427), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n785), .B1(new_n769), .B2(new_n428), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n812), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n826), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n813), .B(new_n825), .C1(new_n835), .C2(KEYINPUT51), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n648), .B(new_n625), .C1(new_n647), .C2(new_n674), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n687), .A2(new_n235), .A3(new_n639), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n625), .A2(new_n427), .A3(new_n643), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n664), .A3(new_n716), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n707), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n707), .A2(new_n837), .A3(new_n840), .A4(KEYINPUT52), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n681), .A2(new_n684), .A3(new_n700), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n692), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n847), .A2(new_n733), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n621), .A2(new_n311), .A3(new_n602), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT110), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n621), .A2(new_n311), .A3(new_n612), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT111), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n717), .B1(new_n619), .B2(new_n620), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT111), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n612), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n591), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n611), .A2(new_n234), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n626), .A2(new_n643), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n638), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n428), .A3(new_n502), .A4(new_n811), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n731), .A2(new_n704), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n735), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n630), .A2(new_n581), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n857), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n848), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT53), .B1(new_n845), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n848), .A2(new_n865), .A3(KEYINPUT112), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n735), .A2(new_n861), .A3(new_n862), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n849), .A2(KEYINPUT110), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT110), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n853), .B2(new_n602), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n852), .B(new_n855), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n592), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n630), .A2(new_n581), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n870), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n847), .A2(new_n733), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n869), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n868), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n843), .A2(KEYINPUT113), .A3(new_n844), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n841), .A2(new_n883), .A3(new_n842), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n867), .B(KEYINPUT54), .C1(new_n881), .C2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n880), .B1(new_n845), .B2(new_n866), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT114), .B1(new_n847), .B2(new_n733), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n870), .A2(new_n875), .A3(new_n876), .A4(KEYINPUT53), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n847), .A2(KEYINPUT114), .A3(new_n733), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n882), .A3(new_n884), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT118), .B1(new_n836), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n886), .A2(new_n894), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n784), .A2(new_n786), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n812), .B1(new_n900), .B2(new_n827), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n901), .B2(new_n826), .ZN(new_n902));
  INV_X1    g716(.A(new_n825), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n808), .B1(new_n831), .B2(new_n832), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n834), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n905), .B2(new_n806), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n897), .A2(new_n898), .A3(new_n902), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n814), .A2(new_n217), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n896), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n639), .A2(new_n584), .A3(new_n671), .A4(new_n718), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT109), .Z(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n664), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT49), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n807), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT49), .B1(new_n678), .B2(new_n679), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n912), .A2(new_n667), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n909), .A2(new_n916), .ZN(G75));
  AOI21_X1  g731(.A(new_n228), .B1(new_n887), .B2(new_n892), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n918), .A2(G210), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n376), .A2(new_n408), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n406), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n217), .A2(G952), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n919), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n924), .A2(new_n929), .ZN(G51));
  AOI211_X1 g744(.A(new_n228), .B(new_n762), .C1(new_n887), .C2(new_n892), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n739), .B(KEYINPUT57), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n887), .A2(new_n892), .A3(new_n893), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n893), .B1(new_n887), .B2(new_n892), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n931), .B1(new_n935), .B2(new_n485), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT120), .B1(new_n936), .B2(new_n925), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  INV_X1    g752(.A(new_n485), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT114), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n878), .A2(new_n940), .ZN(new_n941));
  NOR4_X1   g755(.A1(new_n857), .A2(new_n863), .A3(new_n880), .A4(new_n864), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n942), .A3(new_n891), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n885), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n877), .A2(new_n878), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n843), .A2(new_n844), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT53), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT54), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n894), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n939), .B1(new_n949), .B2(new_n932), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n938), .B(new_n926), .C1(new_n950), .C2(new_n931), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n937), .A2(new_n951), .ZN(G54));
  NAND3_X1  g766(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n953), .A2(new_n287), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n287), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n925), .ZN(G60));
  XNOR2_X1  g770(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n229), .A2(new_n228), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n957), .B(new_n958), .Z(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n886), .B2(new_n894), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n926), .B1(new_n960), .B2(new_n597), .ZN(new_n961));
  INV_X1    g775(.A(new_n959), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n597), .B(new_n962), .C1(new_n933), .C2(new_n934), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n887), .B2(new_n892), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n925), .B1(new_n970), .B2(new_n623), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n530), .B(KEYINPUT123), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G66));
  NOR2_X1   g790(.A1(new_n857), .A2(new_n864), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n847), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n217), .ZN(new_n979));
  OAI21_X1  g793(.A(G953), .B1(new_n298), .B2(new_n403), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(KEYINPUT124), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(KEYINPUT124), .B2(new_n979), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n921), .B1(G898), .B2(new_n217), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(G69));
  INV_X1    g798(.A(new_n640), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n580), .B1(new_n815), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n652), .A2(new_n778), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n669), .A2(new_n707), .A3(new_n837), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n669), .A2(KEYINPUT62), .A3(new_n707), .A4(new_n837), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n780), .A3(new_n789), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n217), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n540), .B1(new_n545), .B2(KEYINPUT30), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(new_n282), .Z(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n996), .B1(G900), .B2(G953), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n838), .A2(new_n730), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n767), .A2(new_n770), .A3(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n733), .A2(new_n707), .A3(new_n735), .A4(new_n837), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n780), .A2(new_n789), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n999), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n997), .A2(new_n998), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n217), .B1(G227), .B2(G900), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1007), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n997), .A2(new_n998), .A3(new_n1009), .A4(new_n1005), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n993), .B2(new_n978), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n570), .A3(new_n660), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n661), .A2(new_n635), .A3(new_n1013), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n867), .B(new_n1016), .C1(new_n881), .C2(new_n885), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n766), .B(new_n737), .C1(new_n829), .C2(new_n830), .ZN(new_n1021));
  AOI21_X1  g835(.A(KEYINPUT107), .B1(new_n769), .B2(new_n738), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1002), .B1(new_n1023), .B2(new_n779), .ZN(new_n1024));
  INV_X1    g838(.A(new_n978), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1024), .A2(new_n789), .A3(new_n1025), .A4(new_n1001), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n635), .B1(new_n1026), .B2(new_n1013), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1020), .B1(new_n1027), .B2(new_n925), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1013), .B1(new_n1004), .B2(new_n978), .ZN(new_n1029));
  INV_X1    g843(.A(new_n635), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1031), .A2(KEYINPUT126), .A3(new_n926), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1019), .B1(new_n1028), .B2(new_n1032), .ZN(G57));
endmodule


