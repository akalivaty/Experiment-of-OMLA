//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G110), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT72), .B1(new_n196), .B2(G119), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT72), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(new_n193), .A3(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(G119), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT24), .B(G110), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n198), .A2(new_n199), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT73), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT16), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n215), .A2(new_n207), .A3(new_n208), .A4(G125), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n210), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n210), .A2(new_n214), .A3(G146), .A4(new_n216), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n206), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G125), .B(G140), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n218), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n198), .A2(new_n199), .B1(new_n204), .B2(new_n205), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n191), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT74), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n204), .ZN(new_n230));
  INV_X1    g044(.A(new_n205), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n230), .A2(new_n231), .B1(G110), .B2(new_n232), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n212), .A2(KEYINPUT16), .A3(G140), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n222), .A2(KEYINPUT16), .B1(new_n234), .B2(new_n215), .ZN(new_n235));
  AOI21_X1  g049(.A(G146), .B1(new_n235), .B2(new_n210), .ZN(new_n236));
  INV_X1    g050(.A(new_n220), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n230), .A2(new_n231), .B1(G110), .B2(new_n232), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n220), .A3(new_n223), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT74), .A3(new_n191), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n229), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n240), .A3(new_n190), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT75), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT75), .A4(new_n190), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT76), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n250));
  AOI21_X1  g064(.A(G902), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n243), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n253), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n243), .A2(new_n248), .A3(new_n255), .A4(new_n251), .ZN(new_n256));
  INV_X1    g070(.A(G217), .ZN(new_n257));
  INV_X1    g071(.A(G902), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n257), .B1(G234), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n254), .A2(KEYINPUT77), .A3(new_n256), .A4(new_n259), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n243), .A2(new_n248), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n259), .A2(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n269));
  NOR2_X1   g083(.A1(G472), .A2(G902), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT64), .B(G131), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G137), .ZN(new_n277));
  INV_X1    g091(.A(G137), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(G137), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n274), .A2(new_n277), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n280), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n276), .A2(G137), .ZN(new_n283));
  OAI21_X1  g097(.A(G131), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n218), .A2(G143), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT1), .ZN(new_n286));
  XNOR2_X1  g100(.A(G143), .B(G146), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(G128), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n218), .A2(G143), .ZN(new_n290));
  INV_X1    g104(.A(G143), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G146), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n281), .B(new_n284), .C1(new_n288), .C2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n290), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT0), .B(G128), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n287), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G131), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n281), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n295), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI211_X1 g118(.A(KEYINPUT65), .B(new_n299), .C1(new_n281), .C2(new_n301), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n273), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n193), .A2(G116), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G119), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT2), .B(G113), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n299), .A2(KEYINPUT66), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n297), .B(new_n314), .C1(new_n287), .C2(new_n298), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n301), .A2(new_n281), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT30), .A3(new_n295), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n306), .A2(new_n312), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n306), .A2(KEYINPUT67), .A3(new_n312), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT68), .B(G237), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n325), .A2(new_n188), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G210), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT27), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT27), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n329), .A3(G210), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G101), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n328), .B2(new_n330), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n312), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n318), .A2(new_n335), .A3(new_n295), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n272), .B1(new_n324), .B2(new_n338), .ZN(new_n339));
  AOI211_X1 g153(.A(KEYINPUT31), .B(new_n337), .C1(new_n322), .C2(new_n323), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n318), .A2(new_n295), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT69), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n312), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n318), .A2(KEYINPUT69), .A3(new_n295), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT28), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n304), .A2(new_n305), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n336), .B1(new_n348), .B2(new_n335), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT28), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n334), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n271), .B1(new_n341), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n269), .B1(new_n354), .B2(KEYINPUT32), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n324), .A2(new_n338), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT31), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n324), .A2(new_n272), .A3(new_n338), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n270), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(KEYINPUT70), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n334), .B1(new_n347), .B2(new_n350), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n339), .A2(new_n340), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n271), .A2(new_n361), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT71), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n351), .A2(new_n334), .ZN(new_n369));
  INV_X1    g183(.A(new_n336), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n322), .B2(new_n323), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n352), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n342), .A2(new_n312), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n336), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT28), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n347), .A2(KEYINPUT29), .A3(new_n334), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n258), .ZN(new_n378));
  OAI21_X1  g192(.A(G472), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT71), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n359), .A2(new_n380), .A3(new_n366), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n368), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n268), .B1(new_n363), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  XNOR2_X1  g198(.A(G116), .B(G122), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n385), .A2(new_n386), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(G116), .B(G122), .Z(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT92), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n387), .A3(G107), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n291), .A2(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n196), .A2(G143), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n390), .A2(new_n393), .B1(new_n276), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT13), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT93), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n394), .B2(new_n398), .ZN(new_n400));
  AOI211_X1 g214(.A(KEYINPUT93), .B(KEYINPUT13), .C1(new_n291), .C2(G128), .ZN(new_n401));
  OAI221_X1 g215(.A(new_n395), .B1(new_n398), .B2(new_n394), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n402), .A2(KEYINPUT94), .A3(G134), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT94), .B1(new_n402), .B2(G134), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT95), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n397), .B(KEYINPUT95), .C1(new_n403), .C2(new_n404), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n396), .B(new_n276), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n308), .A2(KEYINPUT14), .A3(G122), .ZN(new_n410));
  OAI211_X1 g224(.A(G107), .B(new_n410), .C1(new_n391), .C2(KEYINPUT14), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n390), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT9), .B(G234), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n413), .A2(new_n257), .A3(G953), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n407), .A2(new_n408), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT96), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n408), .A3(new_n412), .ZN(new_n418));
  INV_X1    g232(.A(new_n414), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n412), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n405), .B2(new_n406), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n422), .A2(KEYINPUT96), .A3(new_n408), .A4(new_n414), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n258), .ZN(new_n425));
  INV_X1    g239(.A(G478), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(KEYINPUT15), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n427), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(G475), .A2(G902), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT91), .Z(new_n432));
  NAND3_X1  g246(.A1(new_n325), .A2(G214), .A3(new_n188), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n291), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n325), .A2(G143), .A3(G214), .A4(new_n188), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n274), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n236), .A2(new_n237), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n437), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(new_n274), .A3(new_n435), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n438), .B(new_n439), .C1(new_n442), .C2(KEYINPUT17), .ZN(new_n443));
  XNOR2_X1  g257(.A(G113), .B(G122), .ZN(new_n444));
  INV_X1    g258(.A(G104), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(KEYINPUT18), .A2(G131), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n222), .A2(new_n218), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n436), .A2(new_n447), .B1(new_n223), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n436), .B2(new_n447), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n443), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n222), .B(KEYINPUT19), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n218), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT90), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(KEYINPUT90), .A3(new_n218), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n442), .A2(new_n220), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n446), .B1(new_n457), .B2(new_n450), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n432), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT20), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n443), .A2(new_n446), .A3(new_n450), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n457), .A2(new_n450), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n446), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n432), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n446), .B1(new_n443), .B2(new_n450), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n258), .B1(new_n451), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G475), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G234), .ZN(new_n471));
  INV_X1    g285(.A(G237), .ZN(new_n472));
  OAI211_X1 g286(.A(G902), .B(G953), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT97), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(G898), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n188), .A2(G952), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n471), .B2(new_n472), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n430), .A2(new_n470), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n290), .A2(new_n292), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n484), .A2(new_n196), .B1(KEYINPUT1), .B2(new_n285), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n293), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n212), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n212), .B2(new_n299), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n188), .A2(G224), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT86), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n488), .B(new_n491), .Z(new_n492));
  XNOR2_X1  g306(.A(G110), .B(G122), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n493), .B(KEYINPUT8), .Z(new_n494));
  NAND3_X1  g308(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT5), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G113), .B1(new_n307), .B2(KEYINPUT5), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n310), .A2(new_n311), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT3), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT78), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(KEYINPUT78), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n384), .A2(G104), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G101), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n445), .A2(G107), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT78), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT3), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n445), .A2(G107), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT79), .B1(new_n384), .B2(G104), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n504), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n507), .A2(KEYINPUT79), .ZN(new_n515));
  OAI21_X1  g329(.A(G101), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n494), .B1(new_n500), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n497), .B1(new_n495), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n496), .A2(KEYINPUT88), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n499), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n518), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n492), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT81), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n512), .A2(new_n527), .A3(new_n516), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n512), .B2(new_n516), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n500), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n508), .A2(KEYINPUT3), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n509), .B1(new_n510), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n507), .B1(new_n502), .B2(new_n504), .ZN(new_n533));
  OAI21_X1  g347(.A(G101), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT4), .A3(new_n512), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n384), .A2(G104), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n509), .B2(new_n510), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n506), .B1(new_n537), .B2(new_n505), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n535), .A2(new_n312), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n530), .A2(new_n493), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n530), .A2(KEYINPUT85), .A3(new_n493), .A4(new_n541), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n526), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n530), .A2(new_n541), .ZN(new_n549));
  INV_X1    g363(.A(new_n493), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n548), .A3(new_n550), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n488), .B(new_n490), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n553), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n546), .B2(new_n551), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT87), .B1(new_n559), .B2(new_n554), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n547), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n555), .A2(new_n556), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n559), .A2(KEYINPUT87), .A3(new_n554), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n562), .A3(new_n547), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n483), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G221), .B1(new_n413), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G140), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n188), .A2(G227), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n572), .B(new_n573), .Z(new_n574));
  INV_X1    g388(.A(KEYINPUT80), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n293), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n287), .A2(KEYINPUT80), .A3(new_n289), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n485), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n517), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n486), .B1(new_n512), .B2(new_n516), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n317), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(KEYINPUT12), .B(new_n317), .C1(new_n579), .C2(new_n580), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n485), .B2(new_n293), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n528), .B2(new_n529), .ZN(new_n587));
  INV_X1    g401(.A(new_n317), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n585), .B1(new_n578), .B2(new_n517), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n316), .A2(new_n535), .A3(new_n540), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n313), .A2(new_n315), .B1(new_n538), .B2(new_n539), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n485), .A2(new_n576), .A3(new_n577), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n512), .A3(new_n516), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n535), .A2(new_n594), .B1(new_n596), .B2(new_n585), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(KEYINPUT82), .A3(new_n588), .A4(new_n587), .ZN(new_n598));
  AOI221_X4 g412(.A(new_n574), .B1(new_n583), .B2(new_n584), .C1(new_n593), .C2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n574), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n593), .A2(new_n598), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n587), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n317), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n571), .B(new_n258), .C1(new_n599), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT84), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n574), .B1(new_n593), .B2(new_n598), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n583), .A2(new_n584), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n593), .A2(new_n598), .B1(new_n602), .B2(new_n317), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n600), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT84), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n571), .A4(new_n258), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n601), .A2(new_n608), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n615), .A2(new_n574), .B1(new_n607), .B2(new_n603), .ZN(new_n616));
  OAI21_X1  g430(.A(G469), .B1(new_n616), .B2(G902), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n601), .A2(new_n603), .A3(new_n600), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n593), .A2(new_n598), .B1(new_n584), .B2(new_n583), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n620), .B1(new_n600), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n571), .B1(new_n622), .B2(new_n258), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT83), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n614), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n481), .A2(new_n569), .A3(new_n570), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n383), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT98), .B(G101), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G3));
  INV_X1    g443(.A(new_n570), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n623), .B(new_n618), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n631), .B2(new_n614), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n359), .A2(new_n258), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n634), .A2(new_n360), .A3(new_n268), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n564), .A2(new_n637), .A3(new_n568), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n424), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n420), .A2(KEYINPUT33), .A3(new_n415), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n426), .A2(G902), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n425), .A2(new_n426), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n645), .A2(new_n470), .A3(new_n479), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n562), .B1(new_n567), .B2(new_n547), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n483), .B1(new_n647), .B2(KEYINPUT99), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n638), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n636), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT34), .B(G104), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  INV_X1    g466(.A(new_n470), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n430), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n479), .B(KEYINPUT100), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n638), .A2(new_n648), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n632), .A2(new_n658), .A3(new_n635), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NAND2_X1  g476(.A1(new_n634), .A2(new_n360), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n632), .A2(new_n569), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n241), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n265), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n262), .A2(new_n263), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n262), .A2(new_n671), .A3(new_n263), .A4(new_n668), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n481), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n665), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  AND3_X1   g491(.A1(new_n673), .A2(new_n570), .A3(new_n625), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n365), .A2(KEYINPUT71), .A3(new_n367), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n380), .B1(new_n359), .B2(new_n366), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n355), .A3(new_n362), .A4(new_n379), .ZN(new_n682));
  INV_X1    g496(.A(new_n478), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n683), .B1(new_n474), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n430), .A2(new_n653), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n678), .A2(new_n659), .A3(new_n682), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XOR2_X1   g504(.A(new_n685), .B(KEYINPUT39), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n632), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT40), .Z(new_n693));
  AOI21_X1  g507(.A(new_n653), .B1(new_n429), .B2(new_n428), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n482), .A3(new_n670), .A4(new_n672), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n371), .A2(new_n352), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n258), .B1(new_n375), .B2(new_n334), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n681), .A2(new_n355), .A3(new_n362), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n564), .A2(new_n568), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n693), .A2(new_n696), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  AOI221_X4 g519(.A(new_n685), .B1(new_n466), .B2(new_n469), .C1(new_n643), .C2(new_n644), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n678), .A2(new_n659), .A3(new_n682), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT104), .B(G146), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G48));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  INV_X1    g524(.A(new_n614), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n601), .A2(new_n603), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n574), .ZN(new_n713));
  AOI21_X1  g527(.A(G902), .B1(new_n713), .B2(new_n609), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n571), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n711), .A2(new_n630), .A3(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n716), .B(new_n268), .C1(new_n363), .C2(new_n382), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n710), .B1(new_n717), .B2(new_n649), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT70), .B1(new_n360), .B2(new_n361), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n269), .B(KEYINPUT32), .C1(new_n359), .C2(new_n270), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n382), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n267), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n649), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT105), .A4(new_n716), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT41), .B(G113), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n723), .A2(new_n658), .A3(new_n659), .A4(new_n716), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NAND4_X1  g544(.A1(new_n674), .A2(new_n682), .A3(new_n659), .A4(new_n716), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  XNOR2_X1  g546(.A(new_n267), .B(KEYINPUT107), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n375), .A2(KEYINPUT28), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n734), .B1(new_n735), .B2(new_n346), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n347), .A2(KEYINPUT106), .A3(new_n376), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n352), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n341), .A2(new_n738), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n633), .A2(G472), .B1(new_n739), .B2(new_n270), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n733), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n715), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n614), .A2(new_n742), .A3(new_n570), .A4(new_n656), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n638), .A2(new_n648), .A3(new_n694), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  AND3_X1   g562(.A1(new_n673), .A2(new_n706), .A3(new_n740), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n659), .A3(new_n716), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  OAI221_X1 g565(.A(new_n379), .B1(new_n365), .B2(new_n367), .C1(new_n354), .C2(KEYINPUT32), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(new_n733), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n706), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n612), .B1(new_n714), .B2(new_n571), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n605), .A2(KEYINPUT84), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n617), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT108), .A3(new_n570), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n564), .A2(new_n482), .A3(new_n568), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n623), .B1(new_n606), .B2(new_n613), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n630), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT42), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n383), .A2(new_n763), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n706), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(G131), .Z(G33));
  NAND3_X1  g583(.A1(new_n564), .A2(new_n482), .A3(new_n568), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n757), .A2(new_n570), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n760), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n723), .A2(new_n688), .A3(new_n772), .A4(new_n758), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(new_n645), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT43), .B1(new_n775), .B2(new_n470), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n645), .A2(new_n777), .A3(new_n653), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n776), .A2(new_n663), .A3(new_n673), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n759), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(G469), .B1(new_n616), .B2(KEYINPUT45), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n786), .A2(KEYINPUT109), .B1(KEYINPUT45), .B2(new_n616), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(KEYINPUT109), .B2(new_n786), .ZN(new_n788));
  NAND2_X1  g602(.A1(G469), .A2(G902), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT46), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n711), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(KEYINPUT46), .A3(new_n789), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n630), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(new_n691), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n781), .A2(new_n782), .A3(KEYINPUT110), .A4(new_n759), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n785), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  XOR2_X1   g611(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n798));
  OR2_X1    g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n793), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n759), .A2(new_n267), .A3(new_n706), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n682), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT112), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n799), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n262), .A2(new_n263), .A3(new_n668), .A4(new_n686), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n761), .A2(new_n630), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n746), .A2(new_n700), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n368), .A2(new_n381), .A3(new_n699), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n810), .B1(new_n363), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT119), .B1(new_n813), .B2(new_n745), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n689), .A2(new_n707), .A3(new_n750), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT52), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n689), .A2(new_n707), .A3(new_n750), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n811), .A2(new_n814), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n673), .A2(new_n706), .A3(new_n740), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n763), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n772), .A2(new_n749), .A3(KEYINPUT115), .A4(new_n758), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n430), .A2(new_n470), .A3(new_n685), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n678), .A2(new_n682), .A3(new_n759), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n773), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n823), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n826), .A2(new_n827), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(KEYINPUT116), .A3(new_n773), .A4(new_n830), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n768), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n674), .A2(new_n665), .B1(new_n744), .B2(new_n746), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n658), .A2(new_n632), .A3(new_n569), .A4(new_n635), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n729), .A3(new_n731), .A4(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n645), .A2(new_n470), .A3(new_n656), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n632), .A2(new_n569), .A3(new_n635), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n383), .B2(new_n626), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n840), .B(KEYINPUT114), .C1(new_n383), .C2(new_n626), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n838), .A2(new_n845), .A3(new_n726), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n822), .A2(new_n835), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n689), .A2(new_n750), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n689), .A2(KEYINPUT118), .A3(new_n750), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n707), .A3(new_n820), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n817), .B1(KEYINPUT52), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n846), .A4(new_n835), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n849), .A2(new_n850), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n847), .A2(new_n848), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n835), .A2(new_n846), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n835), .A2(new_n846), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n864), .A3(new_n856), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n865), .B2(new_n848), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n859), .B1(new_n866), .B2(new_n850), .ZN(new_n867));
  INV_X1    g681(.A(new_n716), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n776), .A2(new_n778), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n868), .A2(new_n869), .A3(new_n478), .A4(new_n770), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n753), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT48), .Z(new_n872));
  NOR3_X1   g686(.A1(new_n741), .A2(new_n869), .A3(new_n478), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n659), .A3(new_n716), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n775), .A2(new_n653), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n700), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n267), .A2(new_n478), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n716), .A3(new_n759), .A4(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n874), .B(new_n477), .C1(new_n876), .C2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n873), .A2(new_n759), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n799), .A2(new_n802), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n711), .A2(new_n715), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n630), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n882), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n870), .A2(new_n673), .A3(new_n740), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n775), .A2(new_n653), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n703), .A2(new_n868), .A3(new_n482), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n889), .A2(KEYINPUT50), .A3(new_n873), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT50), .B1(new_n889), .B2(new_n873), .ZN(new_n891));
  OAI221_X1 g705(.A(new_n887), .B1(new_n879), .B2(new_n888), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n881), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n872), .B(new_n880), .C1(new_n893), .C2(KEYINPUT51), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(KEYINPUT51), .B2(new_n893), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n867), .A2(new_n895), .B1(G952), .B2(G953), .ZN(new_n896));
  NOR4_X1   g710(.A1(new_n775), .A2(new_n470), .A3(new_n630), .A4(new_n483), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT49), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n897), .B(new_n733), .C1(new_n898), .C2(new_n884), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT113), .Z(new_n900));
  AOI21_X1  g714(.A(new_n703), .B1(new_n898), .B2(new_n884), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n877), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n896), .A2(new_n902), .ZN(G75));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n188), .A2(G952), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n258), .B1(new_n849), .B2(new_n857), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT56), .B1(new_n907), .B2(G210), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n559), .B(new_n554), .Z(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT55), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n906), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(G210), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n913), .B(new_n258), .C1(new_n849), .C2(new_n857), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n914), .A2(KEYINPUT56), .A3(new_n910), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n904), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n908), .A2(new_n911), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n910), .B1(new_n914), .B2(KEYINPUT56), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT121), .A4(new_n906), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(G51));
  XOR2_X1   g734(.A(new_n789), .B(KEYINPUT57), .Z(new_n921));
  AOI21_X1  g735(.A(new_n850), .B1(new_n849), .B2(new_n857), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n858), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(KEYINPUT122), .B(new_n921), .C1(new_n858), .C2(new_n922), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n611), .A3(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n907), .B(new_n787), .C1(KEYINPUT109), .C2(new_n786), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n905), .B1(new_n927), .B2(new_n928), .ZN(G54));
  AND3_X1   g743(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n906), .B1(new_n930), .B2(new_n463), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n463), .B2(new_n930), .ZN(G60));
  NOR2_X1   g746(.A1(new_n858), .A2(new_n922), .ZN(new_n933));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT59), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n640), .A2(new_n641), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n906), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n867), .A2(new_n935), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n640), .A2(new_n641), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n849), .B2(new_n857), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n906), .B1(new_n943), .B2(new_n264), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n667), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n947), .ZN(new_n951));
  INV_X1    g765(.A(new_n948), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n950), .B(new_n951), .C1(new_n952), .C2(new_n944), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n949), .A2(new_n953), .ZN(G66));
  NOR2_X1   g768(.A1(new_n846), .A2(G953), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT124), .Z(new_n956));
  INV_X1    g770(.A(G224), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n475), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n559), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(G898), .B2(new_n188), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(G69));
  NAND2_X1  g777(.A1(new_n306), .A2(new_n319), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT126), .Z(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(new_n452), .Z(new_n966));
  AND3_X1   g780(.A1(new_n853), .A2(new_n707), .A3(new_n854), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n704), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n770), .B1(new_n876), .B2(new_n654), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(new_n723), .A3(new_n632), .A4(new_n691), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n806), .A2(new_n796), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n969), .A2(new_n973), .A3(new_n976), .A4(new_n970), .ZN(new_n977));
  AOI211_X1 g791(.A(G953), .B(new_n966), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n966), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n794), .A2(new_n746), .A3(new_n753), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n764), .A2(new_n980), .A3(new_n767), .A4(new_n773), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n796), .A2(new_n981), .A3(new_n806), .A4(new_n967), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n188), .ZN(new_n983));
  NAND2_X1  g797(.A1(G900), .A2(G953), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n978), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n983), .A2(new_n984), .ZN(new_n988));
  NAND2_X1  g802(.A1(G227), .A2(G900), .ZN(new_n989));
  AND4_X1   g803(.A1(G953), .A2(new_n988), .A3(new_n989), .A4(new_n966), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n987), .A2(new_n990), .ZN(G72));
  INV_X1    g805(.A(new_n697), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n975), .A2(new_n846), .A3(new_n977), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n995), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n982), .B2(new_n846), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n906), .B1(new_n998), .B2(new_n372), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n992), .A2(new_n372), .A3(new_n995), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n866), .A2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n996), .A2(new_n999), .A3(new_n1001), .ZN(G57));
endmodule


