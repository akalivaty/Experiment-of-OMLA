//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944;
  XOR2_X1   g000(.A(KEYINPUT24), .B(G110), .Z(new_n187));
  XNOR2_X1  g001(.A(G119), .B(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT82), .Z(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT83), .B1(new_n191), .B2(G128), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n192), .A2(KEYINPUT23), .B1(new_n191), .B2(G128), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(KEYINPUT23), .B2(new_n192), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G110), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G125), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n198), .B1(new_n202), .B2(new_n196), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(G146), .B(new_n198), .C1(new_n202), .C2(new_n196), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n190), .A2(new_n195), .A3(new_n207), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n194), .A2(G110), .B1(new_n188), .B2(new_n187), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n209), .B(new_n206), .C1(G146), .C2(new_n202), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(G221), .A3(G234), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n213), .B(KEYINPUT22), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n214), .B(G137), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n211), .B(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT25), .B1(new_n217), .B2(G902), .ZN(new_n218));
  INV_X1    g032(.A(G217), .ZN(new_n219));
  INV_X1    g033(.A(G902), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(G234), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n217), .A2(G902), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(KEYINPUT25), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n217), .B(KEYINPUT84), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n221), .A2(G902), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n224), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(G475), .A2(G902), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT95), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT95), .A2(G143), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G237), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n212), .A3(G214), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(G237), .A2(G953), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n233), .A2(G214), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT18), .A2(G131), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n240), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n233), .A2(new_n234), .B1(new_n239), .B2(G214), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT18), .B(G131), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT96), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n202), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G125), .B(G140), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT96), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n247), .A2(new_n249), .A3(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n202), .A2(G146), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n242), .B(new_n245), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G113), .B(G122), .ZN(new_n253));
  INV_X1    g067(.A(G104), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(G131), .B1(new_n243), .B2(new_n244), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n238), .A2(new_n257), .A3(new_n240), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT17), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT17), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n205), .B(new_n206), .C1(new_n256), .C2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n252), .B(new_n255), .C1(new_n260), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT19), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n202), .A2(KEYINPUT19), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n204), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n259), .A3(new_n206), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n255), .B1(new_n267), .B2(new_n252), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT97), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n263), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI211_X1 g084(.A(KEYINPUT97), .B(new_n255), .C1(new_n267), .C2(new_n252), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n230), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT20), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT20), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(new_n230), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G478), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(KEYINPUT15), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G116), .B(G122), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT14), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G107), .ZN(new_n283));
  INV_X1    g097(.A(G122), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G116), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n285), .B2(KEYINPUT14), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n282), .A2(new_n286), .B1(new_n283), .B2(new_n280), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT100), .ZN(new_n288));
  INV_X1    g102(.A(G128), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(G143), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n232), .A2(KEYINPUT100), .A3(G128), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n289), .A2(G143), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G134), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n292), .A2(G134), .A3(new_n293), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n280), .B(G107), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT98), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n280), .B(new_n283), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT98), .ZN(new_n303));
  INV_X1    g117(.A(new_n297), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT99), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n292), .B1(KEYINPUT13), .B2(new_n293), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n295), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n298), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n311), .A2(new_n219), .A3(G953), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n298), .B(new_n312), .C1(new_n305), .C2(new_n309), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n279), .B1(new_n316), .B2(new_n220), .ZN(new_n317));
  AOI211_X1 g131(.A(G902), .B(new_n278), .C1(new_n314), .C2(new_n315), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n212), .A2(G952), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(G234), .B2(G237), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT21), .B(G898), .Z(new_n323));
  NAND2_X1  g137(.A1(G234), .A2(G237), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n324), .A2(G902), .A3(G953), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n252), .B1(new_n260), .B2(new_n262), .ZN(new_n328));
  INV_X1    g142(.A(new_n255), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n263), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n220), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G475), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n276), .A2(new_n319), .A3(new_n327), .A4(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT101), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n273), .A2(new_n275), .B1(G475), .B2(new_n332), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n337), .A2(KEYINPUT101), .A3(new_n327), .A4(new_n319), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT0), .B(G128), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT64), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n204), .A2(G143), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n232), .A2(G146), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G143), .B(G146), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT64), .B1(new_n348), .B2(new_n341), .ZN(new_n349));
  AND2_X1   g163(.A1(KEYINPUT0), .A2(G128), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n347), .A2(new_n349), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT3), .B1(new_n254), .B2(G107), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n283), .A3(G104), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n254), .A2(G107), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G101), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT85), .B(G101), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(new_n353), .A3(new_n356), .A4(new_n355), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n352), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT4), .B1(new_n357), .B2(G101), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n351), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT86), .B1(new_n254), .B2(G107), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n356), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n254), .A2(KEYINPUT86), .A3(G107), .ZN(new_n366));
  OAI21_X1  g180(.A(G101), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n367), .A2(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT69), .ZN(new_n369));
  AOI21_X1  g183(.A(G128), .B1(new_n344), .B2(new_n345), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n232), .A2(KEYINPUT1), .A3(G146), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n369), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(KEYINPUT69), .B(new_n371), .C1(new_n348), .C2(G128), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n348), .A2(new_n375), .A3(G128), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n368), .A2(new_n377), .A3(KEYINPUT10), .ZN(new_n378));
  INV_X1    g192(.A(new_n376), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n371), .B1(new_n348), .B2(G128), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n367), .B(new_n360), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n363), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n295), .A2(G137), .ZN(new_n385));
  INV_X1    g199(.A(G137), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT65), .B1(new_n386), .B2(G134), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT11), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT65), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n390), .B1(new_n295), .B2(G137), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT11), .ZN(new_n392));
  OAI21_X1  g206(.A(G131), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(KEYINPUT11), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n387), .A2(new_n388), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n257), .A4(new_n385), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(KEYINPUT66), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT66), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n398), .B(G131), .C1(new_n389), .C2(new_n392), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n384), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n363), .A2(new_n378), .A3(new_n383), .A4(new_n400), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT88), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n384), .A2(new_n405), .A3(new_n401), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G140), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n212), .A2(G227), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n381), .B1(new_n368), .B2(new_n377), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n401), .A2(new_n411), .B1(KEYINPUT87), .B2(KEYINPUT12), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(KEYINPUT87), .B2(KEYINPUT12), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT12), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n401), .A2(new_n411), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n403), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n410), .B1(new_n417), .B2(new_n409), .ZN(new_n418));
  INV_X1    g232(.A(G469), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n220), .ZN(new_n420));
  INV_X1    g234(.A(new_n409), .ZN(new_n421));
  INV_X1    g235(.A(new_n404), .ZN(new_n422));
  INV_X1    g236(.A(new_n406), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n409), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(G469), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n419), .A2(new_n220), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT2), .B(G113), .Z(new_n432));
  XNOR2_X1  g246(.A(G116), .B(G119), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(KEYINPUT5), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n191), .A3(G116), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(G113), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n368), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n432), .A2(new_n433), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n434), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n361), .B2(new_n362), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G122), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT89), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n439), .A2(new_n442), .A3(new_n447), .A4(new_n444), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n443), .A2(new_n445), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n449), .B2(KEYINPUT90), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n443), .A2(new_n453), .A3(KEYINPUT6), .A4(new_n445), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  MUX2_X1   g269(.A(new_n377), .B(new_n351), .S(G125), .Z(new_n456));
  NAND2_X1  g270(.A1(new_n212), .A2(G224), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT91), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n377), .A2(G125), .ZN(new_n461));
  NAND2_X1  g275(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n461), .B(new_n462), .C1(new_n200), .C2(new_n351), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(KEYINPUT7), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n456), .A2(new_n464), .A3(new_n462), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n439), .A2(KEYINPUT92), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n438), .A2(new_n434), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n367), .A2(new_n360), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OR3_X1    g285(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT92), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n444), .B(KEYINPUT8), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n466), .A2(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n446), .A2(new_n448), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G210), .B1(G237), .B2(G902), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n460), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n460), .A2(new_n477), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n478), .B(KEYINPUT94), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G214), .B1(G237), .B2(G902), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n340), .A2(new_n431), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G472), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT67), .B1(new_n295), .B2(G137), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT67), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n386), .A3(G134), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n491), .A3(new_n385), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G131), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(KEYINPUT68), .A3(G131), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n396), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT70), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n495), .A2(KEYINPUT70), .A3(new_n396), .A4(new_n496), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n377), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n397), .A2(new_n351), .A3(new_n399), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n488), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n377), .A2(new_n396), .A3(new_n496), .A4(new_n495), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n502), .A2(new_n504), .A3(new_n488), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n441), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n441), .B(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n501), .A2(new_n507), .A3(new_n502), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(G101), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT73), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n239), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n516), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n510), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT74), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT74), .B1(new_n517), .B2(new_n519), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n508), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT75), .B(KEYINPUT28), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n502), .A2(new_n504), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n441), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n508), .B2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n525), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n522), .A2(KEYINPUT29), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n521), .A2(new_n527), .A3(KEYINPUT29), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n501), .A2(new_n502), .ZN(new_n538));
  INV_X1    g352(.A(new_n507), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n508), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n541), .B2(KEYINPUT28), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n501), .A2(new_n507), .A3(new_n502), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n507), .B1(new_n501), .B2(new_n502), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n537), .B(KEYINPUT28), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n536), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT28), .B1(new_n543), .B2(new_n544), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT79), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n535), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT80), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n220), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n534), .B1(new_n554), .B2(KEYINPUT81), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT81), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n548), .A2(new_n553), .A3(new_n556), .A4(new_n220), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n487), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n505), .B1(new_n538), .B2(KEYINPUT30), .ZN(new_n559));
  INV_X1    g373(.A(new_n441), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n521), .B(new_n508), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT31), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n525), .B1(new_n528), .B2(new_n532), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n506), .A2(new_n564), .A3(new_n521), .A4(new_n508), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT76), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n562), .A2(new_n563), .A3(new_n568), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(G472), .A2(G902), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT77), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n572), .B1(new_n567), .B2(new_n569), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT78), .B(KEYINPUT32), .Z(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n229), .B(new_n486), .C1(new_n558), .C2(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n578), .B(new_n359), .Z(G3));
  NAND2_X1  g393(.A1(new_n570), .A2(new_n220), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n580), .B2(G472), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n228), .A2(new_n431), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n460), .A2(new_n477), .A3(new_n478), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n478), .B1(new_n460), .B2(new_n477), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n484), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(KEYINPUT102), .B(new_n484), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT33), .B1(new_n312), .B2(KEYINPUT103), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n316), .B(new_n591), .Z(new_n592));
  NOR2_X1   g406(.A1(new_n277), .A2(G902), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n316), .A2(new_n220), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n277), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n276), .A2(new_n333), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n590), .A2(new_n327), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n583), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  NOR2_X1   g418(.A1(new_n598), .A2(new_n319), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n590), .A2(new_n327), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n583), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT35), .B(G107), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  NOR2_X1   g424(.A1(new_n216), .A2(KEYINPUT36), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n211), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n226), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n613), .B(KEYINPUT104), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n224), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n486), .A2(new_n581), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT37), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT105), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G110), .ZN(G12));
  AOI21_X1  g433(.A(new_n576), .B1(new_n570), .B2(new_n573), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT32), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n621), .B(new_n572), .C1(new_n567), .C2(new_n569), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n220), .B1(new_n551), .B2(new_n552), .ZN(new_n624));
  AOI211_X1 g438(.A(KEYINPUT80), .B(new_n535), .C1(new_n550), .C2(new_n545), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT81), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n534), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n557), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G472), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n326), .A2(G900), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n322), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n598), .A2(new_n319), .A3(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n634), .A2(new_n430), .A3(new_n429), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(new_n588), .A3(new_n589), .A4(new_n615), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n630), .A2(KEYINPUT106), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  INV_X1    g457(.A(new_n431), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n632), .B(KEYINPUT39), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT40), .Z(new_n647));
  INV_X1    g461(.A(new_n561), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n525), .B2(new_n541), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n649), .B2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n623), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n483), .B(KEYINPUT38), .Z(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n484), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n615), .A2(new_n319), .A3(new_n337), .A4(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n647), .A2(new_n651), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G143), .ZN(G45));
  AOI21_X1  g471(.A(new_n431), .B1(new_n623), .B2(new_n629), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n599), .A2(new_n633), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n588), .A2(new_n589), .A3(new_n615), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT107), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  AOI21_X1  g479(.A(new_n228), .B1(new_n623), .B2(new_n629), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n418), .A2(new_n220), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n420), .ZN(new_n669));
  INV_X1    g483(.A(new_n430), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n601), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT41), .B(G113), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  NOR2_X1   g490(.A1(new_n672), .A2(new_n606), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(G116), .Z(G18));
  NAND2_X1  g492(.A1(new_n671), .A2(new_n339), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n661), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(new_n558), .B2(new_n577), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G119), .ZN(G21));
  NOR2_X1   g496(.A1(new_n337), .A2(new_n319), .ZN(new_n683));
  AND4_X1   g497(.A1(new_n430), .A2(new_n683), .A3(new_n668), .A4(new_n420), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n327), .A2(new_n684), .A3(new_n588), .A4(new_n589), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n528), .B1(new_n550), .B2(new_n545), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n686), .A2(new_n523), .A3(new_n524), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n562), .A2(new_n565), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n580), .A2(G472), .B1(new_n689), .B2(new_n573), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n685), .A2(new_n690), .A3(new_n229), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  NAND4_X1  g506(.A1(new_n659), .A2(new_n671), .A3(new_n588), .A4(new_n589), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n573), .B1(new_n687), .B2(new_n688), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n567), .B2(new_n569), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n694), .B(new_n615), .C1(new_n695), .C2(new_n487), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n200), .ZN(G27));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n483), .A2(new_n670), .A3(new_n654), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n424), .A2(new_n425), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT108), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n425), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(G469), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n420), .A3(new_n428), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n229), .B(new_n708), .C1(new_n558), .C2(new_n577), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n699), .B1(new_n709), .B2(new_n660), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n707), .A2(new_n660), .A3(new_n699), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n575), .B(KEYINPUT32), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n711), .B(new_n229), .C1(new_n558), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G131), .ZN(G33));
  AOI211_X1 g529(.A(new_n228), .B(new_n707), .C1(new_n623), .C2(new_n629), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n634), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G134), .ZN(G36));
  XNOR2_X1  g532(.A(new_n598), .B(KEYINPUT109), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(KEYINPUT43), .A3(new_n597), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n721));
  INV_X1    g535(.A(new_n597), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(new_n598), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT110), .ZN(new_n725));
  INV_X1    g539(.A(new_n581), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n615), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n725), .A2(KEYINPUT44), .A3(new_n726), .A4(new_n615), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n483), .A2(new_n654), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n702), .A2(KEYINPUT45), .A3(new_n704), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n419), .B1(new_n701), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n427), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n420), .B1(new_n736), .B2(KEYINPUT46), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n430), .B(new_n645), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n729), .A2(new_n730), .A3(new_n731), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT111), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n386), .ZN(G39));
  OAI21_X1  g557(.A(new_n430), .B1(new_n737), .B2(new_n738), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n630), .ZN(new_n748));
  INV_X1    g562(.A(new_n731), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n660), .A2(new_n749), .A3(new_n229), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n747), .A2(KEYINPUT112), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n745), .A2(new_n746), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n754), .B1(new_n755), .B2(new_n751), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G140), .ZN(G42));
  NOR2_X1   g572(.A1(G952), .A2(G953), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n712), .A2(new_n558), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n322), .B1(new_n720), .B2(new_n723), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n671), .A3(new_n731), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n760), .A2(new_n762), .A3(new_n228), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT48), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n671), .A2(new_n731), .A3(new_n229), .A4(new_n321), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n651), .A2(new_n765), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n320), .B(new_n764), .C1(new_n600), .C2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n229), .A3(new_n690), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n590), .A3(new_n671), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT118), .Z(new_n771));
  NOR2_X1   g585(.A1(new_n669), .A2(new_n430), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n731), .B(new_n769), .C1(new_n747), .C2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n671), .A2(new_n654), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT114), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n652), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n774), .B1(new_n777), .B2(new_n768), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT50), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(KEYINPUT51), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n766), .A2(new_n337), .A3(new_n722), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n762), .A2(new_n696), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT117), .Z(new_n784));
  OAI211_X1 g598(.A(new_n767), .B(new_n771), .C1(new_n780), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n773), .A2(new_n782), .A3(new_n781), .ZN(new_n787));
  INV_X1    g601(.A(new_n779), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT116), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n785), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n319), .A2(new_n731), .A3(new_n337), .A4(new_n632), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n644), .B(new_n794), .C1(new_n558), .C2(new_n577), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n690), .A2(new_n708), .A3(new_n659), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n797), .A2(new_n615), .B1(new_n716), .B2(new_n634), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n714), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n485), .A2(new_n599), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n581), .A2(new_n327), .A3(new_n582), .A4(new_n800), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n578), .A2(new_n681), .A3(new_n691), .A4(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n666), .B(new_n671), .C1(new_n607), .C2(new_n601), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n581), .A2(new_n327), .A3(new_n582), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n483), .A2(new_n605), .A3(new_n484), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n616), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n616), .B(KEYINPUT113), .C1(new_n804), .C2(new_n805), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n802), .A2(new_n803), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n799), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n697), .B1(new_n658), .B2(new_n662), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n590), .A2(new_n683), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n615), .A2(new_n670), .A3(new_n633), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n651), .A2(new_n813), .A3(new_n706), .A4(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n630), .A2(KEYINPUT106), .A3(new_n637), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT106), .B1(new_n630), .B2(new_n637), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n812), .B(new_n815), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n642), .A2(KEYINPUT52), .A3(new_n812), .A4(new_n815), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n811), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT53), .B1(new_n811), .B2(new_n822), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT54), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n820), .A2(new_n821), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n802), .A2(new_n803), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n808), .A2(new_n809), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n714), .A3(new_n829), .A4(new_n798), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n826), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n811), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n759), .B1(new_n793), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n669), .A2(KEYINPUT49), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n722), .A2(new_n670), .A3(new_n654), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n719), .A2(new_n837), .A3(new_n229), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n669), .A2(KEYINPUT49), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n651), .A2(new_n653), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n836), .A2(new_n841), .ZN(G75));
  XOR2_X1   g656(.A(new_n455), .B(new_n459), .Z(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT55), .ZN(new_n844));
  OAI21_X1  g658(.A(G902), .B1(new_n823), .B2(new_n824), .ZN(new_n845));
  INV_X1    g659(.A(G210), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n845), .A2(KEYINPUT119), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(KEYINPUT56), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n845), .B2(new_n846), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n212), .A2(G952), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n845), .A2(KEYINPUT120), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n831), .A2(new_n833), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n855), .A3(G902), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n482), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  XOR2_X1   g671(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n858));
  NAND2_X1  g672(.A1(new_n844), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n852), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n850), .A2(new_n860), .ZN(G51));
  NAND2_X1  g675(.A1(new_n853), .A2(new_n856), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n735), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n825), .A2(new_n834), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n427), .B(KEYINPUT57), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n863), .A2(KEYINPUT122), .B1(new_n418), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n862), .A2(new_n868), .A3(new_n735), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n851), .B1(new_n867), .B2(new_n869), .ZN(G54));
  NOR2_X1   g684(.A1(new_n270), .A2(new_n271), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(KEYINPUT58), .A2(G475), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n855), .B1(new_n854), .B2(G902), .ZN(new_n875));
  AOI211_X1 g689(.A(KEYINPUT120), .B(new_n220), .C1(new_n831), .C2(new_n833), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n852), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n872), .B1(new_n862), .B2(new_n873), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT123), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n871), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n851), .B1(new_n862), .B2(new_n874), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n885), .ZN(G60));
  NAND2_X1  g700(.A1(G478), .A2(G902), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT59), .Z(new_n888));
  NOR2_X1   g702(.A1(new_n835), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n852), .B1(new_n889), .B2(new_n592), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n592), .B2(new_n889), .ZN(G63));
  NOR2_X1   g705(.A1(new_n823), .A2(new_n824), .ZN(new_n892));
  XNOR2_X1  g706(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n893));
  NAND2_X1  g707(.A1(G217), .A2(G902), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n612), .ZN(new_n897));
  INV_X1    g711(.A(new_n225), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n897), .B(new_n852), .C1(new_n898), .C2(new_n896), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(G66));
  NAND3_X1  g715(.A1(new_n323), .A2(G224), .A3(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n810), .B2(G953), .ZN(new_n903));
  INV_X1    g717(.A(G898), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n455), .B1(new_n904), .B2(G953), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n903), .B(new_n905), .ZN(G69));
  AOI21_X1  g720(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n760), .A2(new_n228), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n740), .A2(new_n908), .A3(new_n813), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n741), .A2(new_n717), .A3(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n757), .A2(new_n910), .A3(new_n714), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n642), .A2(new_n812), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT125), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n212), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n264), .A2(new_n265), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n559), .B(new_n915), .Z(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(G900), .B2(G953), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT126), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n916), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n913), .A2(new_n656), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n731), .B1(new_n600), .B2(new_n605), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n924), .A2(new_n646), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n666), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n757), .A2(new_n741), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n922), .A2(new_n923), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n920), .B1(new_n928), .B2(new_n212), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n907), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n907), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n928), .A2(new_n212), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n931), .B(new_n918), .C1(new_n932), .C2(new_n920), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n933), .ZN(G72));
  INV_X1    g748(.A(new_n810), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n922), .A2(new_n935), .A3(new_n923), .A4(new_n927), .ZN(new_n936));
  NAND2_X1  g750(.A1(G472), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT63), .Z(new_n938));
  AOI211_X1 g752(.A(new_n520), .B(new_n510), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n911), .A2(new_n935), .A3(new_n913), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n521), .B(new_n509), .C1(new_n940), .C2(new_n938), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n938), .B1(new_n522), .B2(new_n648), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT127), .Z(new_n943));
  OAI21_X1  g757(.A(new_n852), .B1(new_n892), .B2(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n939), .A2(new_n941), .A3(new_n944), .ZN(G57));
endmodule


