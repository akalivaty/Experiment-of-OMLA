

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739;

  NOR2_X1 U369 ( .A1(n545), .A2(n402), .ZN(n629) );
  XNOR2_X1 U370 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n516) );
  INV_X2 U371 ( .A(KEYINPUT64), .ZN(n409) );
  BUF_X2 U372 ( .A(G119), .Z(n407) );
  NAND2_X2 U373 ( .A1(G214), .A2(n523), .ZN(n660) );
  NOR2_X2 U374 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X2 U375 ( .A(n461), .B(n460), .ZN(n704) );
  XNOR2_X2 U376 ( .A(n492), .B(n416), .ZN(n708) );
  XNOR2_X2 U377 ( .A(G902), .B(KEYINPUT15), .ZN(n608) );
  INV_X1 U378 ( .A(G146), .ZN(n437) );
  NOR2_X1 U379 ( .A1(n398), .A2(n592), .ZN(n657) );
  NOR2_X1 U380 ( .A1(n689), .A2(G902), .ZN(n483) );
  XNOR2_X1 U381 ( .A(n586), .B(KEYINPUT35), .ZN(n735) );
  AND2_X1 U382 ( .A1(n536), .A2(n629), .ZN(n537) );
  XNOR2_X1 U383 ( .A(n581), .B(n447), .ZN(n675) );
  NAND2_X1 U384 ( .A1(n645), .A2(n644), .ZN(n398) );
  XNOR2_X1 U385 ( .A(G101), .B(G119), .ZN(n503) );
  INV_X1 U386 ( .A(KEYINPUT47), .ZN(n414) );
  AND2_X1 U387 ( .A1(n729), .A2(n393), .ZN(n392) );
  NAND2_X1 U388 ( .A1(n538), .A2(n366), .ZN(n365) );
  NOR2_X1 U389 ( .A1(n565), .A2(n537), .ZN(n366) );
  XNOR2_X1 U390 ( .A(n415), .B(n414), .ZN(n538) );
  XNOR2_X1 U391 ( .A(n540), .B(KEYINPUT40), .ZN(n738) );
  NOR2_X1 U392 ( .A1(n531), .A2(n554), .ZN(n627) );
  XNOR2_X1 U393 ( .A(n583), .B(n582), .ZN(n585) );
  XNOR2_X1 U394 ( .A(n364), .B(n363), .ZN(n529) );
  XNOR2_X1 U395 ( .A(n514), .B(n436), .ZN(n386) );
  XNOR2_X1 U396 ( .A(n556), .B(n419), .ZN(n631) );
  XNOR2_X1 U397 ( .A(n655), .B(KEYINPUT104), .ZN(n578) );
  NOR2_X1 U398 ( .A1(n594), .A2(n528), .ZN(n435) );
  BUF_X1 U399 ( .A(n645), .Z(n395) );
  OR2_X2 U400 ( .A1(n380), .A2(n379), .ZN(n655) );
  XNOR2_X1 U401 ( .A(n555), .B(KEYINPUT1), .ZN(n645) );
  XNOR2_X1 U402 ( .A(n497), .B(n496), .ZN(n649) );
  XNOR2_X1 U403 ( .A(n698), .B(n697), .ZN(n700) );
  XNOR2_X1 U404 ( .A(n425), .B(n423), .ZN(n698) );
  XNOR2_X1 U405 ( .A(n512), .B(n352), .ZN(n689) );
  XNOR2_X1 U406 ( .A(n723), .B(n417), .ZN(n416) );
  XNOR2_X1 U407 ( .A(n489), .B(n418), .ZN(n417) );
  INV_X1 U408 ( .A(n503), .ZN(n505) );
  XOR2_X1 U409 ( .A(G137), .B(G140), .Z(n486) );
  XNOR2_X1 U410 ( .A(KEYINPUT16), .B(G110), .ZN(n449) );
  BUF_X1 U411 ( .A(n438), .Z(n347) );
  XNOR2_X1 U412 ( .A(G128), .B(n407), .ZN(n490) );
  XNOR2_X1 U413 ( .A(n490), .B(G110), .ZN(n418) );
  BUF_X1 U414 ( .A(n475), .Z(n348) );
  XNOR2_X1 U415 ( .A(n426), .B(n477), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n426), .B(n477), .ZN(n724) );
  AND2_X1 U417 ( .A1(n737), .A2(n597), .ZN(n596) );
  NOR2_X2 U418 ( .A1(n641), .A2(n611), .ZN(n350) );
  BUF_X1 U419 ( .A(n374), .Z(n351) );
  NOR2_X2 U420 ( .A1(n641), .A2(n611), .ZN(n706) );
  XNOR2_X2 U421 ( .A(n401), .B(n353), .ZN(n532) );
  NOR2_X2 U422 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U423 ( .A(n389), .B(n388), .ZN(n648) );
  INV_X1 U424 ( .A(KEYINPUT21), .ZN(n388) );
  NAND2_X1 U425 ( .A1(n493), .A2(G221), .ZN(n389) );
  NAND2_X1 U426 ( .A1(n381), .A2(n384), .ZN(n380) );
  NAND2_X1 U427 ( .A1(G472), .A2(G902), .ZN(n384) );
  XNOR2_X1 U428 ( .A(n370), .B(KEYINPUT73), .ZN(n508) );
  NAND2_X1 U429 ( .A1(n716), .A2(n371), .ZN(n370) );
  INV_X1 U430 ( .A(G237), .ZN(n371) );
  NAND2_X1 U431 ( .A1(n413), .A2(n648), .ZN(n412) );
  INV_X1 U432 ( .A(n528), .ZN(n413) );
  NAND2_X1 U433 ( .A1(n578), .A2(n557), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n462), .B(G478), .ZN(n551) );
  AND2_X1 U435 ( .A1(n649), .A2(n355), .ZN(n644) );
  NOR2_X1 U436 ( .A1(n649), .A2(n587), .ZN(n588) );
  XNOR2_X1 U437 ( .A(n474), .B(n473), .ZN(n542) );
  NOR2_X1 U438 ( .A1(n698), .A2(G902), .ZN(n474) );
  XOR2_X1 U439 ( .A(KEYINPUT5), .B(G137), .Z(n507) );
  INV_X1 U440 ( .A(n618), .ZN(n431) );
  INV_X1 U441 ( .A(KEYINPUT44), .ZN(n428) );
  XOR2_X1 U442 ( .A(G107), .B(G104), .Z(n450) );
  XNOR2_X1 U443 ( .A(G101), .B(G110), .ZN(n478) );
  NOR2_X1 U444 ( .A1(n365), .A2(n564), .ZN(n378) );
  OR2_X1 U445 ( .A1(G902), .A2(G237), .ZN(n523) );
  XNOR2_X1 U446 ( .A(n434), .B(KEYINPUT6), .ZN(n433) );
  INV_X1 U447 ( .A(KEYINPUT103), .ZN(n434) );
  XNOR2_X1 U448 ( .A(n469), .B(n476), .ZN(n424) );
  XNOR2_X1 U449 ( .A(n520), .B(n394), .ZN(n470) );
  XNOR2_X1 U450 ( .A(G143), .B(G140), .ZN(n394) );
  AND2_X2 U451 ( .A1(n375), .A2(n439), .ZN(n729) );
  NOR2_X1 U452 ( .A1(n734), .A2(n440), .ZN(n439) );
  XNOR2_X1 U453 ( .A(n376), .B(n566), .ZN(n375) );
  INV_X1 U454 ( .A(n638), .ZN(n440) );
  XNOR2_X1 U455 ( .A(n526), .B(n525), .ZN(n539) );
  XNOR2_X1 U456 ( .A(n524), .B(KEYINPUT85), .ZN(n525) );
  NAND2_X1 U457 ( .A1(n386), .A2(n385), .ZN(n526) );
  AND2_X1 U458 ( .A1(n662), .A2(n355), .ZN(n443) );
  INV_X1 U459 ( .A(KEYINPUT102), .ZN(n420) );
  NOR2_X1 U460 ( .A1(n708), .A2(G902), .ZN(n497) );
  BUF_X1 U461 ( .A(n730), .Z(n408) );
  NOR2_X1 U462 ( .A1(n408), .A2(G952), .ZN(n709) );
  XOR2_X1 U463 ( .A(KEYINPUT38), .B(n362), .Z(n661) );
  NAND2_X1 U464 ( .A1(n513), .A2(n383), .ZN(n382) );
  INV_X1 U465 ( .A(G902), .ZN(n383) );
  XNOR2_X1 U466 ( .A(n484), .B(KEYINPUT20), .ZN(n493) );
  NAND2_X1 U467 ( .A1(G237), .A2(G234), .ZN(n498) );
  AND2_X1 U468 ( .A1(n435), .A2(n661), .ZN(n385) );
  INV_X1 U469 ( .A(KEYINPUT94), .ZN(n387) );
  XNOR2_X1 U470 ( .A(n360), .B(n511), .ZN(n612) );
  XOR2_X1 U471 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n459) );
  XOR2_X1 U472 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n455) );
  XNOR2_X1 U473 ( .A(KEYINPUT9), .B(KEYINPUT100), .ZN(n454) );
  AND2_X1 U474 ( .A1(n729), .A2(KEYINPUT2), .ZN(n391) );
  INV_X1 U475 ( .A(KEYINPUT30), .ZN(n436) );
  XNOR2_X1 U476 ( .A(n552), .B(KEYINPUT106), .ZN(n584) );
  XNOR2_X1 U477 ( .A(n530), .B(KEYINPUT108), .ZN(n545) );
  INV_X1 U478 ( .A(KEYINPUT28), .ZN(n363) );
  XNOR2_X1 U479 ( .A(n470), .B(n467), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n424), .B(n468), .ZN(n423) );
  NAND2_X1 U481 ( .A1(n556), .A2(n539), .ZN(n540) );
  XNOR2_X1 U482 ( .A(n372), .B(n356), .ZN(n562) );
  INV_X1 U483 ( .A(KEYINPUT32), .ZN(n368) );
  INV_X1 U484 ( .A(KEYINPUT107), .ZN(n419) );
  INV_X1 U485 ( .A(n649), .ZN(n603) );
  INV_X1 U486 ( .A(KEYINPUT86), .ZN(n410) );
  INV_X1 U487 ( .A(KEYINPUT121), .ZN(n404) );
  XOR2_X1 U488 ( .A(n481), .B(n480), .Z(n352) );
  AND2_X1 U489 ( .A1(n523), .A2(G210), .ZN(n353) );
  AND2_X1 U490 ( .A1(n737), .A2(n428), .ZN(n354) );
  XOR2_X1 U491 ( .A(n648), .B(n387), .Z(n355) );
  XNOR2_X1 U492 ( .A(KEYINPUT110), .B(KEYINPUT36), .ZN(n356) );
  XNOR2_X1 U493 ( .A(KEYINPUT65), .B(n548), .ZN(n357) );
  INV_X1 U494 ( .A(n608), .ZN(n393) );
  XOR2_X1 U495 ( .A(n687), .B(n686), .Z(n358) );
  XOR2_X1 U496 ( .A(n604), .B(KEYINPUT66), .Z(n359) );
  INV_X1 U497 ( .A(G953), .ZN(n716) );
  XNOR2_X1 U498 ( .A(n724), .B(n437), .ZN(n512) );
  XNOR2_X1 U499 ( .A(n349), .B(n437), .ZN(n360) );
  BUF_X1 U500 ( .A(n390), .Z(n361) );
  AND2_X1 U501 ( .A1(n374), .A2(n392), .ZN(n609) );
  BUF_X1 U502 ( .A(n532), .Z(n362) );
  AND2_X2 U503 ( .A1(n374), .A2(n391), .ZN(n606) );
  XNOR2_X2 U504 ( .A(n441), .B(n359), .ZN(n374) );
  XNOR2_X1 U505 ( .A(n369), .B(n368), .ZN(n737) );
  NAND2_X1 U506 ( .A1(n438), .A2(n596), .ZN(n367) );
  NOR2_X2 U507 ( .A1(n624), .A2(n735), .ZN(n438) );
  NAND2_X1 U508 ( .A1(n367), .A2(n599), .ZN(n432) );
  XNOR2_X1 U509 ( .A(n400), .B(KEYINPUT95), .ZN(n399) );
  NOR2_X2 U510 ( .A1(n590), .A2(n395), .ZN(n600) );
  NOR2_X1 U511 ( .A1(n590), .A2(n589), .ZN(n369) );
  NAND2_X1 U512 ( .A1(n559), .A2(n631), .ZN(n567) );
  NAND2_X1 U513 ( .A1(n560), .A2(n561), .ZN(n372) );
  BUF_X1 U514 ( .A(n624), .Z(n373) );
  INV_X1 U515 ( .A(n351), .ZN(n396) );
  NAND2_X1 U516 ( .A1(n374), .A2(n716), .ZN(n717) );
  NAND2_X1 U517 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U518 ( .A(n549), .B(n357), .ZN(n377) );
  NOR2_X1 U519 ( .A1(n612), .A2(n382), .ZN(n379) );
  NAND2_X1 U520 ( .A1(n612), .A2(G472), .ZN(n381) );
  AND2_X1 U521 ( .A1(n386), .A2(n435), .ZN(n553) );
  NAND2_X1 U522 ( .A1(n390), .A2(n443), .ZN(n442) );
  XNOR2_X2 U523 ( .A(n577), .B(KEYINPUT0), .ZN(n390) );
  NAND2_X1 U524 ( .A1(n390), .A2(n657), .ZN(n591) );
  NAND2_X1 U525 ( .A1(n390), .A2(n592), .ZN(n593) );
  NAND2_X1 U526 ( .A1(n675), .A2(n361), .ZN(n583) );
  XNOR2_X1 U527 ( .A(n636), .B(KEYINPUT84), .ZN(n564) );
  NOR2_X2 U528 ( .A1(n562), .A2(n563), .ZN(n636) );
  XNOR2_X1 U529 ( .A(n518), .B(n517), .ZN(n445) );
  NAND2_X1 U530 ( .A1(n683), .A2(n608), .ZN(n401) );
  NOR2_X2 U531 ( .A1(n398), .A2(n601), .ZN(n581) );
  AND2_X1 U532 ( .A1(n396), .A2(n605), .ZN(n640) );
  NAND2_X1 U533 ( .A1(n397), .A2(n712), .ZN(n722) );
  XNOR2_X2 U534 ( .A(n397), .B(n444), .ZN(n683) );
  XNOR2_X2 U535 ( .A(n446), .B(n522), .ZN(n397) );
  NAND2_X1 U536 ( .A1(n399), .A2(n664), .ZN(n597) );
  NOR2_X2 U537 ( .A1(n634), .A2(n620), .ZN(n400) );
  NOR2_X2 U538 ( .A1(n593), .A2(n594), .ZN(n620) );
  XNOR2_X2 U539 ( .A(n591), .B(KEYINPUT31), .ZN(n634) );
  INV_X1 U540 ( .A(n362), .ZN(n531) );
  BUF_X1 U541 ( .A(n576), .Z(n402) );
  NOR2_X2 U542 ( .A1(n705), .A2(n709), .ZN(n405) );
  NAND2_X1 U543 ( .A1(n706), .A2(G478), .ZN(n703) );
  NOR2_X2 U544 ( .A1(n701), .A2(n709), .ZN(n702) );
  NAND2_X1 U545 ( .A1(n350), .A2(G475), .ZN(n699) );
  NOR2_X2 U546 ( .A1(n615), .A2(n709), .ZN(n617) );
  NAND2_X1 U547 ( .A1(n350), .A2(G217), .ZN(n707) );
  NOR2_X2 U548 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U549 ( .A(n403), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U550 ( .A1(n688), .A2(n709), .ZN(n403) );
  XNOR2_X1 U551 ( .A(n405), .B(n404), .ZN(G63) );
  XNOR2_X1 U552 ( .A(n406), .B(n358), .ZN(n688) );
  NAND2_X1 U553 ( .A1(n706), .A2(G210), .ZN(n406) );
  XNOR2_X2 U554 ( .A(n409), .B(G953), .ZN(n730) );
  XNOR2_X2 U555 ( .A(G116), .B(KEYINPUT3), .ZN(n504) );
  XNOR2_X2 U556 ( .A(n442), .B(KEYINPUT22), .ZN(n590) );
  XNOR2_X2 U557 ( .A(n483), .B(n482), .ZN(n555) );
  OR2_X2 U558 ( .A1(n598), .A2(KEYINPUT44), .ZN(n599) );
  NOR2_X1 U559 ( .A1(n580), .A2(n579), .ZN(n624) );
  XNOR2_X2 U560 ( .A(n505), .B(n504), .ZN(n519) );
  XNOR2_X2 U561 ( .A(n519), .B(n449), .ZN(n446) );
  XNOR2_X1 U562 ( .A(n411), .B(n410), .ZN(n602) );
  AND2_X1 U563 ( .A1(n600), .A2(n601), .ZN(n411) );
  NOR2_X1 U564 ( .A1(n649), .A2(n412), .ZN(n557) );
  NAND2_X1 U565 ( .A1(n629), .A2(n535), .ZN(n415) );
  XNOR2_X2 U566 ( .A(G146), .B(G125), .ZN(n515) );
  INV_X1 U567 ( .A(n542), .ZN(n550) );
  XNOR2_X2 U568 ( .A(n421), .B(n420), .ZN(n556) );
  NAND2_X1 U569 ( .A1(n542), .A2(n551), .ZN(n421) );
  INV_X1 U570 ( .A(n543), .ZN(n422) );
  XNOR2_X1 U571 ( .A(n426), .B(n445), .ZN(n444) );
  XNOR2_X2 U572 ( .A(n475), .B(KEYINPUT4), .ZN(n426) );
  NAND2_X1 U573 ( .A1(n429), .A2(n427), .ZN(n441) );
  NAND2_X1 U574 ( .A1(n347), .A2(n354), .ZN(n427) );
  XNOR2_X1 U575 ( .A(n430), .B(KEYINPUT87), .ZN(n429) );
  NAND2_X1 U576 ( .A1(n432), .A2(n431), .ZN(n430) );
  XNOR2_X2 U577 ( .A(n655), .B(n433), .ZN(n601) );
  NOR2_X2 U578 ( .A1(n603), .A2(n602), .ZN(n618) );
  XOR2_X1 U579 ( .A(KEYINPUT90), .B(KEYINPUT33), .Z(n447) );
  XNOR2_X1 U580 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n448) );
  INV_X1 U581 ( .A(KEYINPUT45), .ZN(n604) );
  XNOR2_X1 U582 ( .A(n479), .B(n450), .ZN(n481) );
  XNOR2_X1 U583 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U584 ( .A(KEYINPUT88), .ZN(n533) );
  INV_X1 U585 ( .A(G472), .ZN(n513) );
  XNOR2_X1 U586 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U587 ( .A(n612), .B(n448), .ZN(n613) );
  XNOR2_X1 U588 ( .A(n614), .B(n613), .ZN(n615) );
  XOR2_X1 U589 ( .A(G107), .B(G122), .Z(n521) );
  XOR2_X1 U590 ( .A(n521), .B(G116), .Z(n453) );
  XNOR2_X2 U591 ( .A(G128), .B(KEYINPUT78), .ZN(n451) );
  XNOR2_X2 U592 ( .A(n451), .B(G143), .ZN(n475) );
  XNOR2_X1 U593 ( .A(n348), .B(G134), .ZN(n452) );
  XNOR2_X1 U594 ( .A(n453), .B(n452), .ZN(n457) );
  XNOR2_X1 U595 ( .A(n455), .B(n454), .ZN(n456) );
  NAND2_X1 U596 ( .A1(G234), .A2(n730), .ZN(n458) );
  XNOR2_X1 U597 ( .A(n459), .B(n458), .ZN(n491) );
  NAND2_X1 U598 ( .A1(G217), .A2(n491), .ZN(n460) );
  NOR2_X1 U599 ( .A1(n704), .A2(G902), .ZN(n462) );
  XOR2_X1 U600 ( .A(G113), .B(G104), .Z(n520) );
  NAND2_X1 U601 ( .A1(G214), .A2(n508), .ZN(n469) );
  XOR2_X1 U602 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n464) );
  XNOR2_X1 U603 ( .A(G122), .B(KEYINPUT12), .ZN(n463) );
  XNOR2_X1 U604 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U605 ( .A(KEYINPUT97), .B(n465), .Z(n468) );
  XOR2_X1 U606 ( .A(KEYINPUT70), .B(G131), .Z(n476) );
  XNOR2_X1 U607 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n466) );
  XNOR2_X1 U608 ( .A(n466), .B(n515), .ZN(n485) );
  INV_X1 U609 ( .A(n485), .ZN(n467) );
  XOR2_X1 U610 ( .A(KEYINPUT13), .B(KEYINPUT99), .Z(n472) );
  XNOR2_X1 U611 ( .A(KEYINPUT98), .B(G475), .ZN(n471) );
  XNOR2_X1 U612 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U613 ( .A1(n422), .A2(n542), .ZN(n633) );
  XNOR2_X1 U614 ( .A(G134), .B(n476), .ZN(n477) );
  XNOR2_X1 U615 ( .A(n478), .B(n486), .ZN(n479) );
  NAND2_X1 U616 ( .A1(G227), .A2(n730), .ZN(n480) );
  INV_X1 U617 ( .A(G469), .ZN(n482) );
  NAND2_X1 U618 ( .A1(n608), .A2(G234), .ZN(n484) );
  XNOR2_X1 U619 ( .A(n486), .B(n485), .ZN(n723) );
  XOR2_X1 U620 ( .A(KEYINPUT93), .B(KEYINPUT76), .Z(n488) );
  XNOR2_X1 U621 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n487) );
  XNOR2_X1 U622 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U623 ( .A1(G221), .A2(n491), .ZN(n492) );
  XOR2_X1 U624 ( .A(KEYINPUT75), .B(KEYINPUT25), .Z(n495) );
  NAND2_X1 U625 ( .A1(n493), .A2(G217), .ZN(n494) );
  XNOR2_X1 U626 ( .A(n495), .B(n494), .ZN(n496) );
  NAND2_X1 U627 ( .A1(n555), .A2(n644), .ZN(n594) );
  XNOR2_X1 U628 ( .A(n498), .B(KEYINPUT14), .ZN(n499) );
  XNOR2_X1 U629 ( .A(KEYINPUT72), .B(n499), .ZN(n500) );
  NAND2_X1 U630 ( .A1(G952), .A2(n500), .ZN(n673) );
  NOR2_X1 U631 ( .A1(G953), .A2(n673), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n500), .A2(G902), .ZN(n572) );
  OR2_X1 U633 ( .A1(n572), .A2(n408), .ZN(n501) );
  NOR2_X1 U634 ( .A1(G900), .A2(n501), .ZN(n502) );
  NOR2_X1 U635 ( .A1(n574), .A2(n502), .ZN(n528) );
  XNOR2_X1 U636 ( .A(n519), .B(G113), .ZN(n506) );
  XNOR2_X1 U637 ( .A(n507), .B(n506), .ZN(n510) );
  NAND2_X1 U638 ( .A1(G210), .A2(n508), .ZN(n509) );
  NAND2_X1 U639 ( .A1(n578), .A2(n660), .ZN(n514) );
  NAND2_X1 U640 ( .A1(G224), .A2(n730), .ZN(n518) );
  XNOR2_X1 U641 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U642 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U643 ( .A(KEYINPUT39), .ZN(n524) );
  NAND2_X1 U644 ( .A1(n633), .A2(n539), .ZN(n527) );
  XNOR2_X1 U645 ( .A(n527), .B(KEYINPUT111), .ZN(n734) );
  INV_X1 U646 ( .A(n551), .ZN(n543) );
  NOR2_X1 U647 ( .A1(n633), .A2(n556), .ZN(n595) );
  NOR2_X1 U648 ( .A1(KEYINPUT71), .A2(n595), .ZN(n535) );
  NAND2_X1 U649 ( .A1(n529), .A2(n555), .ZN(n530) );
  NAND2_X1 U650 ( .A1(n532), .A2(n660), .ZN(n534) );
  XNOR2_X2 U651 ( .A(n534), .B(n533), .ZN(n560) );
  XNOR2_X2 U652 ( .A(n560), .B(KEYINPUT19), .ZN(n576) );
  AND2_X1 U653 ( .A1(KEYINPUT71), .A2(n595), .ZN(n536) );
  NAND2_X1 U654 ( .A1(n661), .A2(n660), .ZN(n541) );
  XNOR2_X1 U655 ( .A(n541), .B(KEYINPUT109), .ZN(n665) );
  NOR2_X1 U656 ( .A1(n543), .A2(n542), .ZN(n662) );
  NAND2_X1 U657 ( .A1(n665), .A2(n662), .ZN(n544) );
  XNOR2_X1 U658 ( .A(n544), .B(KEYINPUT41), .ZN(n674) );
  INV_X1 U659 ( .A(n545), .ZN(n546) );
  NAND2_X1 U660 ( .A1(n674), .A2(n546), .ZN(n547) );
  XNOR2_X1 U661 ( .A(n547), .B(KEYINPUT42), .ZN(n739) );
  NAND2_X1 U662 ( .A1(n738), .A2(n739), .ZN(n549) );
  XOR2_X1 U663 ( .A(KEYINPUT46), .B(KEYINPUT83), .Z(n548) );
  NOR2_X1 U664 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U665 ( .A1(n553), .A2(n584), .ZN(n554) );
  XNOR2_X1 U666 ( .A(KEYINPUT80), .B(n627), .ZN(n565) );
  INV_X1 U667 ( .A(n395), .ZN(n563) );
  INV_X1 U668 ( .A(n557), .ZN(n558) );
  NOR2_X1 U669 ( .A1(n558), .A2(n601), .ZN(n559) );
  INV_X1 U670 ( .A(n567), .ZN(n561) );
  XOR2_X1 U671 ( .A(KEYINPUT48), .B(KEYINPUT82), .Z(n566) );
  NOR2_X1 U672 ( .A1(n395), .A2(n567), .ZN(n568) );
  NAND2_X1 U673 ( .A1(n568), .A2(n660), .ZN(n569) );
  XNOR2_X1 U674 ( .A(n569), .B(KEYINPUT43), .ZN(n570) );
  NAND2_X1 U675 ( .A1(n570), .A2(n531), .ZN(n638) );
  NOR2_X1 U676 ( .A1(G898), .A2(n716), .ZN(n571) );
  XOR2_X1 U677 ( .A(KEYINPUT92), .B(n571), .Z(n712) );
  NOR2_X1 U678 ( .A1(n572), .A2(n712), .ZN(n573) );
  NOR2_X2 U679 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U680 ( .A(n600), .B(KEYINPUT105), .ZN(n580) );
  OR2_X1 U681 ( .A1(n649), .A2(n578), .ZN(n579) );
  INV_X1 U682 ( .A(KEYINPUT34), .ZN(n582) );
  NAND2_X1 U683 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U684 ( .A1(n645), .A2(n601), .ZN(n587) );
  XNOR2_X1 U685 ( .A(KEYINPUT77), .B(n588), .ZN(n589) );
  INV_X1 U686 ( .A(n655), .ZN(n592) );
  INV_X1 U687 ( .A(n595), .ZN(n664) );
  INV_X1 U688 ( .A(n597), .ZN(n598) );
  INV_X1 U689 ( .A(KEYINPUT2), .ZN(n605) );
  XNOR2_X2 U690 ( .A(n606), .B(KEYINPUT74), .ZN(n641) );
  NAND2_X1 U691 ( .A1(n393), .A2(KEYINPUT2), .ZN(n607) );
  XNOR2_X1 U692 ( .A(n607), .B(KEYINPUT67), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n706), .A2(G472), .ZN(n614) );
  INV_X1 U694 ( .A(KEYINPUT63), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n617), .B(n616), .ZN(G57) );
  XOR2_X1 U696 ( .A(G101), .B(n618), .Z(G3) );
  NAND2_X1 U697 ( .A1(n631), .A2(n620), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(G104), .ZN(G6) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n622) );
  NAND2_X1 U700 ( .A1(n620), .A2(n633), .ZN(n621) );
  XNOR2_X1 U701 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U702 ( .A(G107), .B(n623), .ZN(G9) );
  XOR2_X1 U703 ( .A(n373), .B(G110), .Z(G12) );
  XOR2_X1 U704 ( .A(G128), .B(KEYINPUT29), .Z(n626) );
  NAND2_X1 U705 ( .A1(n629), .A2(n633), .ZN(n625) );
  XNOR2_X1 U706 ( .A(n626), .B(n625), .ZN(G30) );
  XNOR2_X1 U707 ( .A(G143), .B(n627), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n628), .B(KEYINPUT113), .ZN(G45) );
  NAND2_X1 U709 ( .A1(n631), .A2(n629), .ZN(n630) );
  XNOR2_X1 U710 ( .A(n630), .B(G146), .ZN(G48) );
  NAND2_X1 U711 ( .A1(n631), .A2(n634), .ZN(n632) );
  XNOR2_X1 U712 ( .A(n632), .B(G113), .ZN(G15) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U714 ( .A(n635), .B(G116), .ZN(G18) );
  XNOR2_X1 U715 ( .A(G125), .B(n636), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n637), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U717 ( .A(G140), .B(n638), .ZN(G42) );
  NOR2_X1 U718 ( .A1(n729), .A2(KEYINPUT2), .ZN(n639) );
  XNOR2_X1 U719 ( .A(n639), .B(KEYINPUT81), .ZN(n643) );
  NOR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n679) );
  XOR2_X1 U722 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n647) );
  OR2_X1 U723 ( .A1(n395), .A2(n644), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n647), .B(n646), .ZN(n653) );
  NOR2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n651) );
  XNOR2_X1 U726 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n658), .B(KEYINPUT51), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n659), .A2(n674), .ZN(n670) );
  OR2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U737 ( .A1(n675), .A2(n668), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U739 ( .A(KEYINPUT52), .B(n671), .Z(n672) );
  NOR2_X1 U740 ( .A1(n673), .A2(n672), .ZN(n677) );
  AND2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U744 ( .A1(G953), .A2(n680), .ZN(n682) );
  XNOR2_X1 U745 ( .A(KEYINPUT53), .B(KEYINPUT116), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n682), .B(n681), .ZN(G75) );
  XOR2_X1 U747 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n685) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT79), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n685), .B(n684), .ZN(n687) );
  XOR2_X1 U750 ( .A(KEYINPUT89), .B(KEYINPUT54), .Z(n686) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  XNOR2_X1 U752 ( .A(n689), .B(KEYINPUT118), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U754 ( .A1(n350), .A2(G469), .ZN(n692) );
  XNOR2_X1 U755 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U756 ( .A1(n709), .A2(n694), .ZN(G54) );
  XOR2_X1 U757 ( .A(KEYINPUT120), .B(KEYINPUT91), .Z(n696) );
  XNOR2_X1 U758 ( .A(KEYINPUT59), .B(KEYINPUT119), .ZN(n695) );
  XNOR2_X1 U759 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U760 ( .A(n699), .B(n700), .ZN(n701) );
  XNOR2_X1 U761 ( .A(n702), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U762 ( .A(n703), .B(n704), .ZN(n705) );
  XNOR2_X1 U763 ( .A(n707), .B(n708), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n711), .B(KEYINPUT122), .ZN(G66) );
  NAND2_X1 U765 ( .A1(G953), .A2(G224), .ZN(n713) );
  XNOR2_X1 U766 ( .A(KEYINPUT61), .B(n713), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n714), .A2(G898), .ZN(n715) );
  XNOR2_X1 U768 ( .A(KEYINPUT123), .B(n715), .ZN(n719) );
  XOR2_X1 U769 ( .A(n717), .B(KEYINPUT124), .Z(n718) );
  NOR2_X1 U770 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U771 ( .A(KEYINPUT125), .B(n720), .Z(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(G69) );
  XOR2_X1 U773 ( .A(n349), .B(n723), .Z(n728) );
  XOR2_X1 U774 ( .A(G227), .B(n728), .Z(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U776 ( .A1(n726), .A2(G953), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n727), .B(KEYINPUT126), .ZN(n733) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(n408), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(G72) );
  XOR2_X1 U781 ( .A(G134), .B(n734), .Z(G36) );
  XNOR2_X1 U782 ( .A(n735), .B(G122), .ZN(n736) );
  XNOR2_X1 U783 ( .A(n736), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U784 ( .A(n407), .B(n737), .ZN(G21) );
  XNOR2_X1 U785 ( .A(n738), .B(G131), .ZN(G33) );
  XNOR2_X1 U786 ( .A(G137), .B(n739), .ZN(G39) );
endmodule

