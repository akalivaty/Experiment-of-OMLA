//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n606, new_n608, new_n609, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  XOR2_X1   g035(.A(KEYINPUT3), .B(G2104), .Z(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n468));
  XNOR2_X1  g043(.A(new_n467), .B(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  OAI211_X1 g046(.A(KEYINPUT70), .B(G2104), .C1(new_n471), .C2(KEYINPUT69), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT3), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT69), .B1(new_n471), .B2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n472), .A2(new_n475), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n470), .A2(new_n480), .ZN(G160));
  XNOR2_X1  g056(.A(new_n478), .B(KEYINPUT72), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n472), .A2(new_n475), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n484), .A2(G2105), .A3(new_n476), .ZN(new_n485));
  MUX2_X1   g060(.A(G100), .B(G112), .S(G2105), .Z(new_n486));
  AOI22_X1  g061(.A1(new_n485), .A2(G124), .B1(G2104), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n472), .A2(new_n475), .A3(new_n476), .A4(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n491), .A2(KEYINPUT73), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G102), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n491), .B2(KEYINPUT73), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT74), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n484), .A2(new_n499), .A3(new_n476), .A4(new_n490), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT74), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n491), .A2(KEYINPUT73), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n496), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n477), .A2(G138), .ZN(new_n505));
  NOR3_X1   g080(.A1(new_n461), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n478), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n498), .A2(new_n503), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT76), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT77), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(new_n519), .A3(G543), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n516), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n513), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n522), .A2(new_n527), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n520), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT78), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT79), .ZN(new_n537));
  XOR2_X1   g112(.A(new_n537), .B(KEYINPUT7), .Z(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(G89), .B2(new_n526), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n534), .A2(KEYINPUT78), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(new_n539), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(new_n521), .A2(G52), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT80), .B(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n526), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n513), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  XOR2_X1   g124(.A(KEYINPUT81), .B(G43), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n521), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n526), .A2(G81), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n513), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT82), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n520), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n520), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n513), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n526), .B2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G299));
  XNOR2_X1  g146(.A(new_n548), .B(KEYINPUT83), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G301));
  NAND2_X1  g148(.A1(new_n521), .A2(G49), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n526), .A2(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND4_X1  g152(.A1(new_n516), .A2(new_n519), .A3(G48), .A4(G543), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n516), .A2(new_n519), .A3(G86), .A4(new_n525), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n513), .C2(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(new_n526), .A2(G85), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  XNOR2_X1  g158(.A(KEYINPUT84), .B(G47), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n582), .B1(new_n513), .B2(new_n583), .C1(new_n520), .C2(new_n584), .ZN(G290));
  NAND3_X1  g160(.A1(G301), .A2(KEYINPUT85), .A3(G868), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n587));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n572), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n521), .A2(G54), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n513), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n526), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n586), .B(new_n589), .C1(new_n601), .C2(G868), .ZN(G284));
  XOR2_X1   g177(.A(G284), .B(KEYINPUT87), .Z(G321));
  MUX2_X1   g178(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g179(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n601), .B1(new_n606), .B2(G860), .ZN(G148));
  NOR2_X1   g182(.A1(new_n555), .A2(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n600), .A2(G559), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G323));
  XNOR2_X1  g185(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n611));
  XNOR2_X1  g186(.A(G323), .B(new_n611), .ZN(G282));
  NAND2_X1  g187(.A1(new_n485), .A2(G123), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT90), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n482), .A2(G135), .ZN(new_n615));
  AND2_X1   g190(.A1(G111), .A2(G2105), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G99), .B2(new_n477), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n465), .C2(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(G2096), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n477), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n622), .A2(KEYINPUT13), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(KEYINPUT13), .B2(new_n622), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n623), .A2(new_n624), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n619), .A2(new_n620), .A3(new_n628), .ZN(G156));
  XOR2_X1   g204(.A(G2443), .B(G2446), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT92), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT91), .B(KEYINPUT16), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G1341), .B(G1348), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT93), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n641), .B2(new_n642), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n637), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n648), .A3(G14), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(KEYINPUT17), .A3(new_n653), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n653), .B1(new_n652), .B2(KEYINPUT17), .ZN(new_n659));
  INV_X1    g234(.A(new_n654), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n653), .A2(new_n654), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n652), .B1(new_n662), .B2(KEYINPUT17), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n657), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(G2096), .Z(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(G2100), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(G2100), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n670), .C2(new_n674), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT33), .B(G1976), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  MUX2_X1   g266(.A(G6), .B(G305), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G22), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G166), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1971), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n691), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n686), .A2(G24), .ZN(new_n702));
  XOR2_X1   g277(.A(G290), .B(KEYINPUT97), .Z(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n686), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(G1986), .Z(new_n705));
  NOR2_X1   g280(.A1(G25), .A2(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(KEYINPUT95), .B1(G95), .B2(G2105), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g283(.A1(KEYINPUT95), .A2(G95), .A3(G2105), .ZN(new_n709));
  OAI221_X1 g284(.A(G2104), .B1(G107), .B2(new_n477), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT96), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n485), .A2(G119), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n711), .B(new_n712), .C1(G131), .C2(new_n482), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n706), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n700), .A2(new_n701), .A3(new_n705), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT36), .ZN(new_n718));
  NOR2_X1   g293(.A1(G4), .A2(G16), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n601), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1348), .ZN(new_n721));
  NOR2_X1   g296(.A1(G29), .A2(G35), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G162), .B2(G29), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT29), .Z(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT100), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G27), .A2(G29), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G164), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT99), .B(G2078), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G32), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n482), .A2(G141), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT98), .Z(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT26), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n466), .A2(G105), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n738), .B(new_n739), .C1(new_n485), .C2(G129), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n734), .B1(new_n742), .B2(new_n733), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR4_X1   g320(.A1(new_n721), .A2(new_n728), .A3(new_n732), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n733), .A2(G26), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n482), .A2(G140), .ZN(new_n749));
  MUX2_X1   g324(.A(G104), .B(G116), .S(G2105), .Z(new_n750));
  AOI22_X1  g325(.A1(new_n485), .A2(G128), .B1(G2104), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n748), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n686), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n686), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n754), .B1(new_n756), .B2(G1966), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n686), .A2(G5), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G171), .B2(new_n686), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n618), .A2(new_n733), .B1(new_n759), .B2(G1961), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G1961), .B2(new_n759), .ZN(new_n761));
  NOR2_X1   g336(.A1(G16), .A2(G19), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n556), .B2(G16), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1341), .Z(new_n764));
  NAND2_X1  g339(.A1(G160), .A2(G29), .ZN(new_n765));
  AND2_X1   g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  NOR2_X1   g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n733), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(G2084), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT30), .B(G28), .Z(new_n771));
  OAI211_X1 g346(.A(new_n769), .B(new_n770), .C1(G29), .C2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(G2084), .B1(new_n765), .B2(new_n768), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n761), .A2(new_n764), .A3(new_n774), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n757), .B(new_n775), .C1(new_n725), .C2(new_n724), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n482), .A2(G139), .ZN(new_n777));
  INV_X1    g352(.A(G127), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n461), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G115), .B2(G2104), .ZN(new_n780));
  AOI21_X1  g355(.A(KEYINPUT25), .B1(new_n466), .B2(G103), .ZN(new_n781));
  AND3_X1   g356(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n777), .B1(new_n477), .B2(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G33), .B(new_n783), .S(G29), .Z(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G2072), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n756), .A2(G1966), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n686), .A2(G20), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT23), .Z(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G299), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n785), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n727), .B2(new_n726), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n718), .A2(new_n746), .A3(new_n776), .A4(new_n792), .ZN(G150));
  INV_X1    g368(.A(G150), .ZN(G311));
  NOR2_X1   g369(.A1(new_n600), .A2(new_n606), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT38), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n555), .A2(KEYINPUT101), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT102), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n521), .A2(G55), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n526), .A2(G93), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n799), .B(new_n800), .C1(new_n513), .C2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n797), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n798), .B1(new_n797), .B2(new_n802), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n804), .A2(new_n805), .B1(KEYINPUT101), .B2(new_n555), .ZN(new_n806));
  INV_X1    g381(.A(new_n805), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n555), .A2(KEYINPUT101), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n807), .A2(new_n808), .A3(new_n803), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n796), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n813));
  AOI21_X1  g388(.A(G860), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n802), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT37), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(G145));
  XNOR2_X1  g393(.A(new_n488), .B(G160), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(new_n618), .Z(new_n820));
  OR2_X1    g395(.A1(new_n741), .A2(new_n752), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n741), .A2(new_n752), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n492), .A2(new_n497), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n510), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n783), .B(new_n825), .Z(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n482), .A2(G142), .ZN(new_n829));
  INV_X1    g404(.A(G118), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n830), .A2(KEYINPUT103), .A3(G2105), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT103), .B1(new_n830), .B2(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n485), .A2(G130), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n622), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n713), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n821), .A2(new_n822), .A3(new_n826), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n828), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n828), .A2(new_n839), .ZN(new_n843));
  INV_X1    g418(.A(new_n838), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n840), .A2(new_n841), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n820), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n820), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n840), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(G37), .B1(new_n850), .B2(new_n845), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g428(.A1(new_n802), .A2(G868), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n811), .B(new_n609), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n597), .A2(G299), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n597), .A2(G299), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT105), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT105), .B1(new_n597), .B2(G299), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT106), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n858), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT106), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n856), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n855), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n863), .A2(new_n867), .A3(new_n856), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(KEYINPUT41), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n855), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(G290), .B(G288), .ZN(new_n872));
  XNOR2_X1  g447(.A(G303), .B(G305), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT42), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n871), .B(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n854), .B1(new_n877), .B2(G868), .ZN(G295));
  AOI21_X1  g453(.A(new_n854), .B1(new_n877), .B2(G868), .ZN(G331));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n880));
  NAND2_X1  g455(.A1(G286), .A2(G171), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n572), .B2(G286), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n806), .A2(new_n809), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n806), .B2(new_n809), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n868), .B(new_n869), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n865), .A2(new_n862), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n885), .A2(KEYINPUT107), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n870), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n874), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n861), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n885), .B(new_n874), .C1(new_n889), .C2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT43), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n885), .B1(new_n889), .B2(new_n893), .ZN(new_n898));
  INV_X1    g473(.A(new_n874), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n895), .A4(new_n894), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n880), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n892), .B2(new_n896), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n900), .A2(KEYINPUT43), .A3(new_n895), .A4(new_n894), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n903), .A2(new_n906), .ZN(G397));
  AOI21_X1  g482(.A(G1384), .B1(new_n824), .B2(new_n510), .ZN(new_n908));
  XOR2_X1   g483(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n480), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n911), .A2(new_n464), .A3(G40), .A4(new_n469), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n908), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G1996), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n742), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n752), .B(G2067), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n913), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(G1996), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n742), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n920), .A2(KEYINPUT110), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(KEYINPUT110), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n713), .A2(new_n715), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n713), .A2(new_n715), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n913), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(G290), .A2(G1986), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT109), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(G1986), .B2(G290), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(new_n918), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n484), .A2(G138), .A3(new_n477), .A4(new_n476), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n506), .B1(new_n939), .B2(KEYINPUT4), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n500), .A2(new_n502), .A3(new_n496), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n937), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n908), .A2(KEYINPUT112), .A3(KEYINPUT45), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n912), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n511), .A2(new_n938), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n909), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1971), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT50), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n912), .B1(new_n908), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n948), .B2(KEYINPUT50), .ZN(new_n956));
  AOI211_X1 g531(.A(KEYINPUT113), .B(new_n953), .C1(new_n511), .C2(new_n938), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n952), .B1(G2090), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G303), .A2(G8), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT55), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(G8), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n908), .A2(new_n947), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G8), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n688), .A2(G1976), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT52), .ZN(new_n970));
  INV_X1    g545(.A(G1976), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  OR2_X1    g548(.A1(G305), .A2(G1981), .ZN(new_n974));
  NAND2_X1  g549(.A1(G305), .A2(G1981), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n974), .A2(KEYINPUT49), .A3(new_n975), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n967), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n970), .A2(new_n973), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n963), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n511), .A2(new_n938), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n910), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n947), .B1(new_n908), .B2(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n947), .B(KEYINPUT116), .C1(new_n908), .C2(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1966), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G2084), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(new_n954), .C1(new_n956), .C2(new_n957), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n966), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G168), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT63), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n959), .A2(G8), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n982), .B(new_n997), .C1(new_n962), .C2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n912), .B1(new_n942), .B2(KEYINPUT50), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n511), .A2(new_n953), .A3(new_n938), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(G2090), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n951), .B2(new_n950), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n961), .B1(new_n1004), .B2(new_n966), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n963), .A2(new_n1005), .A3(new_n981), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n996), .B1(new_n1006), .B2(new_n995), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n981), .A2(G8), .A3(new_n959), .A4(new_n962), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n688), .A2(new_n971), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT114), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(KEYINPUT114), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n980), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n974), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n967), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1008), .A2(new_n1014), .A3(KEYINPUT115), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n999), .A2(new_n1007), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1956), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n511), .A2(new_n953), .A3(new_n938), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n947), .B1(new_n908), .B2(new_n953), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n946), .A2(new_n947), .A3(new_n949), .A4(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1002), .A2(KEYINPUT117), .A3(new_n1020), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n570), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n566), .B2(new_n565), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT57), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n570), .A2(KEYINPUT119), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n570), .A2(KEYINPUT119), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1033), .A2(new_n1034), .B1(new_n566), .B2(new_n565), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1032), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1029), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n1041));
  INV_X1    g616(.A(G1348), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n958), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n964), .A2(G2067), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  AOI211_X1 g621(.A(KEYINPUT120), .B(new_n1044), .C1(new_n958), .C2(new_n1042), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT117), .B1(new_n1002), .B2(new_n1020), .ZN(new_n1049));
  AOI211_X1 g624(.A(new_n1024), .B(G1956), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n1038), .A3(new_n1027), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n601), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1040), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT61), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1038), .B1(new_n1051), .B2(new_n1027), .ZN(new_n1056));
  AND4_X1   g631(.A1(new_n1038), .A2(new_n1025), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT122), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1059));
  NOR2_X1   g634(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n946), .A2(new_n914), .A3(new_n947), .A4(new_n949), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n964), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1065), .B2(new_n556), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n555), .B(new_n1060), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1059), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1058), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1040), .A2(new_n1052), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1055), .B1(new_n1070), .B2(KEYINPUT122), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT60), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n600), .ZN(new_n1074));
  OR3_X1    g649(.A1(new_n1046), .A2(new_n1047), .A3(KEYINPUT60), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT60), .B(new_n601), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1054), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n989), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(G2078), .ZN(new_n1081));
  INV_X1    g656(.A(G2078), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n946), .A2(new_n1082), .A3(new_n947), .A4(new_n949), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1079), .A2(new_n1081), .B1(new_n1083), .B2(new_n1080), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT124), .B(G1961), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n958), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(G301), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1084), .A2(KEYINPUT125), .A3(G301), .A4(new_n1086), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1083), .A2(new_n1080), .ZN(new_n1093));
  INV_X1    g668(.A(new_n946), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n947), .B(new_n1081), .C1(new_n908), .C2(new_n910), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1086), .B(new_n1093), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1096), .B2(G171), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1091), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G286), .A2(G8), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT123), .ZN(new_n1100));
  INV_X1    g675(.A(new_n954), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT113), .B1(new_n983), .B2(new_n953), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n948), .A2(new_n955), .A3(KEYINPUT50), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1104), .A2(new_n992), .B1(new_n990), .B2(new_n989), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT51), .B(new_n1100), .C1(new_n1105), .C2(new_n966), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1099), .B(KEYINPUT123), .Z(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n994), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n991), .A2(new_n993), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1106), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n963), .A2(new_n1005), .A3(new_n981), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1096), .A2(new_n572), .ZN(new_n1114));
  AOI21_X1  g689(.A(G301), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1092), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1098), .A2(new_n1112), .A3(new_n1113), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1019), .B1(new_n1078), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1112), .A2(KEYINPUT62), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1113), .B(new_n1115), .C1(new_n1112), .C2(KEYINPUT62), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AND4_X1   g697(.A1(new_n1005), .A2(new_n1115), .A3(new_n963), .A4(new_n981), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(KEYINPUT126), .C1(KEYINPUT62), .C2(new_n1112), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1119), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n936), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n919), .A2(KEYINPUT46), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n919), .A2(KEYINPUT46), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n913), .B1(new_n741), .B2(new_n916), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT47), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n933), .A2(new_n913), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT48), .Z(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n931), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(G2067), .B2(new_n752), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1136), .B2(new_n913), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1126), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n1140));
  NAND3_X1  g714(.A1(new_n666), .A2(G319), .A3(new_n667), .ZN(new_n1141));
  OAI211_X1 g715(.A(new_n684), .B(new_n649), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g716(.A(new_n1142), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1143));
  NAND4_X1  g717(.A1(new_n1143), .A2(new_n852), .A3(new_n904), .A4(new_n905), .ZN(G225));
  INV_X1    g718(.A(G225), .ZN(G308));
endmodule


