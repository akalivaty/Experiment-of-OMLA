//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1310, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(new_n206), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n209), .B(new_n214), .C1(new_n215), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n215), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT64), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT2), .B(G226), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G68), .B(G77), .Z(new_n235));
  XOR2_X1   g0035(.A(G50), .B(G58), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  NAND2_X1  g0041(.A1(G33), .A2(G41), .ZN(new_n242));
  NAND3_X1  g0042(.A1(new_n242), .A2(G1), .A3(G13), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G1698), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  AND2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n247), .A2(G223), .B1(G77), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n245), .A2(G222), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT66), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n244), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT65), .B(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI211_X1 g0059(.A(G1), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n243), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n260), .B1(G226), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n256), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G200), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n256), .A2(G190), .A3(new_n264), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n212), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n203), .A2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G50), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n273), .A2(new_n276), .B1(new_n277), .B2(new_n270), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR3_X1   g0081(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n282));
  OAI22_X1  g0082(.A1(new_n279), .A2(new_n281), .B1(new_n282), .B2(new_n204), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n204), .A2(G33), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT67), .ZN(new_n285));
  INV_X1    g0085(.A(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT8), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT8), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G58), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n283), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n272), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n278), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n293), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n268), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT10), .B1(new_n267), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n297), .A2(new_n295), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n252), .A2(new_n255), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n264), .B1(new_n301), .B2(new_n243), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n300), .A2(new_n303), .A3(new_n304), .A4(new_n268), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n296), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G179), .B2(new_n302), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n292), .A2(G77), .A3(new_n269), .A4(new_n274), .ZN(new_n310));
  INV_X1    g0110(.A(G77), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n270), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G20), .A2(G77), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  INV_X1    g0115(.A(new_n290), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n314), .B1(new_n284), .B2(new_n315), .C1(new_n316), .C2(new_n281), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n313), .B1(new_n317), .B2(new_n272), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n245), .A2(G232), .A3(new_n253), .ZN(new_n319));
  INV_X1    g0119(.A(G107), .ZN(new_n320));
  INV_X1    g0120(.A(G238), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n319), .B1(new_n320), .B2(new_n245), .C1(new_n246), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n244), .ZN(new_n323));
  INV_X1    g0123(.A(G41), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT65), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT65), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G41), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n203), .B(G274), .C1(new_n328), .C2(G45), .ZN(new_n329));
  INV_X1    g0129(.A(G244), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n262), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n318), .B1(new_n333), .B2(new_n307), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n322), .B2(new_n244), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n323), .A2(G190), .A3(new_n332), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(new_n318), .C1(new_n266), .C2(new_n335), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n306), .A2(new_n309), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT68), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT68), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n306), .A2(new_n341), .A3(new_n344), .A4(new_n309), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT69), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n253), .A2(G226), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n250), .B2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n245), .A2(KEYINPUT69), .A3(G226), .A4(new_n253), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(G232), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n243), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n263), .A2(G238), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n329), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT13), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n356), .A2(new_n329), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT13), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n353), .B1(new_n348), .B2(new_n349), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(new_n243), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G200), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n285), .A2(G77), .ZN(new_n365));
  INV_X1    g0165(.A(G68), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT11), .A3(new_n272), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT12), .B1(new_n269), .B2(G68), .ZN(new_n370));
  OR3_X1    g0170(.A1(new_n269), .A2(KEYINPUT12), .A3(G68), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n203), .B2(G20), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n370), .A2(new_n371), .B1(new_n273), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT11), .B1(new_n368), .B2(new_n272), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n358), .A2(new_n362), .A3(KEYINPUT70), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT70), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(KEYINPUT13), .C1(new_n355), .C2(new_n357), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n336), .B1(new_n379), .B2(new_n381), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT71), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n363), .B2(G169), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n363), .A2(G169), .A3(new_n387), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n376), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n343), .A2(new_n345), .A3(new_n383), .A4(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n329), .B1(new_n227), .B2(new_n262), .ZN(new_n395));
  INV_X1    g0195(.A(G226), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G1698), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n245), .B(new_n397), .C1(G223), .C2(G1698), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n243), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G179), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n395), .B2(new_n400), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n245), .B2(G20), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n366), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  NOR2_X1   g0211(.A1(G58), .A2(G68), .ZN(new_n412));
  OAI21_X1  g0212(.A(G20), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G159), .ZN(new_n414));
  NOR4_X1   g0214(.A1(new_n414), .A2(KEYINPUT72), .A3(G20), .A4(G33), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT72), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n280), .B2(G159), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n413), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n406), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n272), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT73), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(KEYINPUT73), .B(new_n413), .C1(new_n415), .C2(new_n417), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT7), .B1(new_n250), .B2(new_n204), .ZN(new_n426));
  NOR4_X1   g0226(.A1(new_n248), .A2(new_n249), .A3(new_n407), .A4(G20), .ZN(new_n427));
  OAI21_X1  g0227(.A(G68), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(KEYINPUT74), .A3(KEYINPUT16), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n408), .A2(new_n409), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n423), .A2(new_n424), .B1(new_n431), .B2(G68), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT74), .B1(new_n432), .B2(KEYINPUT16), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n421), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n273), .A2(new_n290), .A3(new_n274), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n269), .B2(new_n290), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT75), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n405), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT18), .ZN(new_n440));
  INV_X1    g0240(.A(new_n424), .ZN(new_n441));
  INV_X1    g0241(.A(G33), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n204), .A2(new_n442), .A3(G159), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT72), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n280), .A2(new_n416), .A3(G159), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT73), .B1(new_n446), .B2(new_n413), .ZN(new_n447));
  OAI211_X1 g0247(.A(KEYINPUT16), .B(new_n428), .C1(new_n441), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT74), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n420), .B1(new_n450), .B2(new_n429), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n404), .B1(new_n451), .B2(new_n437), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT76), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n452), .B2(new_n454), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n440), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n401), .A2(G190), .ZN(new_n458));
  OAI21_X1  g0258(.A(G200), .B1(new_n395), .B2(new_n400), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n434), .A2(new_n438), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n451), .A2(new_n437), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(KEYINPUT17), .A3(new_n460), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n457), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT77), .B1(new_n394), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n393), .A2(new_n383), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(KEYINPUT68), .B2(new_n342), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT77), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT76), .B1(new_n439), .B2(KEYINPUT18), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n466), .B1(new_n475), .B2(new_n440), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n471), .A2(new_n472), .A3(new_n476), .A4(new_n345), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n320), .B1(KEYINPUT83), .B2(KEYINPUT25), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n269), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n270), .A2(KEYINPUT83), .A3(KEYINPUT25), .A4(new_n320), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n203), .A2(G33), .ZN(new_n483));
  AND4_X1   g0283(.A1(new_n212), .A2(new_n269), .A3(new_n271), .A4(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n481), .A2(new_n482), .B1(new_n484), .B2(G107), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n204), .B(G87), .C1(new_n248), .C2(new_n249), .ZN(new_n487));
  NAND2_X1  g0287(.A1(KEYINPUT80), .A2(KEYINPUT22), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n245), .A2(new_n204), .A3(G87), .A4(new_n488), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT23), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n204), .B2(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n320), .A2(KEYINPUT23), .A3(G20), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT81), .B1(new_n498), .B2(G20), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT81), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(new_n204), .A3(G33), .A4(G116), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n492), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n292), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n492), .B(new_n503), .C1(KEYINPUT82), .C2(KEYINPUT24), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n486), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n509));
  OAI211_X1 g0309(.A(G250), .B(new_n253), .C1(new_n248), .C2(new_n249), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n244), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT5), .B1(new_n325), .B2(new_n327), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT5), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n203), .B(G45), .C1(new_n515), .C2(G41), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n244), .A2(new_n257), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G264), .B(new_n243), .C1(new_n514), .C2(new_n516), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n513), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n307), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n513), .A2(new_n519), .A3(new_n336), .A4(new_n520), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n508), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n504), .A2(new_n505), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(new_n272), .A3(new_n507), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n521), .A2(new_n266), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n521), .A2(G190), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(new_n485), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n531), .A2(new_n204), .ZN(new_n532));
  INV_X1    g0332(.A(G87), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n320), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT79), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G87), .A2(G97), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(KEYINPUT79), .A3(new_n320), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n532), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n204), .B(G68), .C1(new_n248), .C2(new_n249), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n284), .B2(new_n534), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n272), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n315), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(new_n269), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n484), .A2(new_n546), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n321), .A2(new_n253), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n330), .A2(G1698), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(new_n248), .C2(new_n249), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n243), .B1(new_n553), .B2(new_n498), .ZN(new_n554));
  INV_X1    g0354(.A(G250), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n259), .B2(G1), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n203), .A2(new_n257), .A3(G45), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n243), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n336), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n550), .B(new_n561), .C1(G169), .C2(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n531), .A2(new_n204), .ZN(new_n563));
  NOR4_X1   g0363(.A1(new_n536), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT79), .B1(new_n538), .B2(new_n320), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n541), .A3(new_n543), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n547), .B1(new_n567), .B2(new_n272), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n560), .A2(G190), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n484), .A2(G87), .ZN(new_n570));
  OAI21_X1  g0370(.A(G200), .B1(new_n554), .B2(new_n559), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n525), .A2(new_n530), .A3(new_n562), .A4(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G270), .B(new_n243), .C1(new_n514), .C2(new_n516), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n519), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n484), .A2(G116), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n269), .A2(G116), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n271), .A2(new_n212), .B1(G20), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(G33), .A2(G283), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n204), .C1(G33), .C2(new_n534), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(KEYINPUT20), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT20), .B1(new_n580), .B2(new_n582), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n576), .B(new_n578), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(new_n253), .C1(new_n248), .C2(new_n249), .ZN(new_n587));
  OAI211_X1 g0387(.A(G264), .B(G1698), .C1(new_n248), .C2(new_n249), .ZN(new_n588));
  OR2_X1    g0388(.A1(KEYINPUT3), .A2(G33), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT3), .A2(G33), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(G303), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n244), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n575), .A2(new_n586), .A3(G179), .A4(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n519), .A3(new_n574), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n595), .A2(new_n596), .A3(G169), .A4(new_n586), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n580), .A2(new_n582), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n583), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n577), .B1(new_n484), .B2(G116), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n307), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n595), .B1(new_n603), .B2(new_n596), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n594), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n586), .B1(new_n596), .B2(G200), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n378), .B2(new_n596), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT4), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(G1698), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(G244), .C1(new_n249), .C2(new_n248), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n330), .B1(new_n589), .B2(new_n590), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n581), .C1(new_n613), .C2(KEYINPUT4), .ZN(new_n614));
  OAI21_X1  g0414(.A(G250), .B1(new_n248), .B2(new_n249), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n253), .B1(new_n615), .B2(KEYINPUT4), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT78), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n555), .B1(new_n589), .B2(new_n590), .ZN(new_n618));
  OAI21_X1  g0418(.A(G1698), .B1(new_n618), .B2(new_n610), .ZN(new_n619));
  OAI21_X1  g0419(.A(G244), .B1(new_n248), .B2(new_n249), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(new_n610), .B1(G33), .B2(G283), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT78), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n619), .A2(new_n621), .A3(new_n622), .A4(new_n612), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n617), .A2(new_n244), .A3(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(G257), .B(new_n243), .C1(new_n514), .C2(new_n516), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n519), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n336), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT6), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n629), .A2(new_n534), .A3(G107), .ZN(new_n630));
  XNOR2_X1  g0430(.A(G97), .B(G107), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n632), .A2(new_n204), .B1(new_n311), .B2(new_n281), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n320), .B1(new_n408), .B2(new_n409), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n272), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n269), .A2(G97), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n484), .B2(G97), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n619), .A2(new_n621), .A3(new_n612), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n243), .B1(new_n639), .B2(KEYINPUT78), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n626), .B1(new_n640), .B2(new_n623), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n628), .B(new_n638), .C1(new_n641), .C2(G169), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n624), .A2(G190), .A3(new_n627), .ZN(new_n643));
  INV_X1    g0443(.A(new_n637), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n631), .A2(new_n629), .ZN(new_n645));
  INV_X1    g0445(.A(new_n630), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n431), .A2(G107), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n644), .B1(new_n650), .B2(new_n272), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n643), .B(new_n651), .C1(new_n641), .C2(new_n266), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n573), .A2(new_n609), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n478), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT84), .ZN(G372));
  NAND2_X1  g0456(.A1(new_n624), .A2(new_n627), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n657), .B2(new_n307), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n638), .B1(new_n657), .B2(G200), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n628), .A2(new_n658), .B1(new_n659), .B2(new_n643), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT87), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n553), .A2(new_n498), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n662), .A2(new_n244), .B1(KEYINPUT85), .B2(new_n558), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT85), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n243), .A2(new_n556), .A3(new_n557), .A4(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n266), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n545), .A2(new_n548), .A3(new_n570), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT86), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n558), .A2(KEYINPUT85), .ZN(new_n669));
  NOR2_X1   g0469(.A1(G238), .A2(G1698), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n330), .B2(G1698), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n671), .A2(new_n245), .B1(G33), .B2(G116), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n665), .B(new_n669), .C1(new_n672), .C2(new_n243), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G200), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT86), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(new_n568), .A3(new_n675), .A4(new_n570), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n668), .A2(new_n569), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n307), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n550), .A3(new_n561), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n677), .A2(new_n530), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n660), .A2(new_n661), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n508), .A2(new_n524), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n605), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n677), .A2(new_n530), .A3(new_n679), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT87), .B1(new_n653), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n562), .A2(new_n572), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT26), .B1(new_n642), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n679), .B(KEYINPUT88), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n677), .A2(new_n679), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n692), .A2(KEYINPUT26), .A3(new_n642), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n478), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n452), .A2(new_n454), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n440), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n334), .A2(new_n337), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n699), .A2(new_n383), .B1(new_n391), .B2(new_n392), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n698), .B1(new_n700), .B2(new_n466), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n306), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n702), .A2(new_n309), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n696), .A2(new_n703), .ZN(G369));
  NAND3_X1  g0504(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n586), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n605), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n713), .B(new_n714), .C1(new_n609), .C2(new_n711), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n525), .A2(new_n710), .ZN(new_n718));
  INV_X1    g0518(.A(new_n710), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n530), .B1(new_n508), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n718), .B1(new_n525), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n605), .A2(new_n719), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT90), .Z(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(new_n721), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n718), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n207), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n328), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n203), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n537), .A2(new_n579), .A3(new_n539), .ZN(new_n732));
  INV_X1    g0532(.A(new_n729), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n731), .A2(new_n732), .B1(new_n210), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n710), .B1(new_n687), .B2(new_n694), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n683), .A2(new_n685), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n653), .A2(KEYINPUT94), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT94), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n642), .A2(new_n652), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT95), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT26), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n642), .B2(new_n688), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT93), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(KEYINPUT93), .B(new_n746), .C1(new_n642), .C2(new_n688), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n692), .A2(new_n642), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n746), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT95), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n740), .A2(new_n741), .A3(new_n753), .A4(new_n743), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n745), .A2(new_n690), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n739), .B1(new_n755), .B2(new_n719), .ZN(new_n756));
  INV_X1    g0556(.A(G330), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n513), .A2(new_n520), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n554), .A2(new_n336), .A3(new_n559), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n759), .A2(new_n575), .A3(new_n760), .A4(new_n593), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n758), .B1(new_n657), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n560), .A2(G179), .A3(new_n520), .A4(new_n513), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n596), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n641), .A2(new_n764), .A3(KEYINPUT30), .ZN(new_n765));
  AND3_X1   g0565(.A1(new_n596), .A2(new_n336), .A3(new_n673), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n657), .A2(new_n766), .A3(new_n521), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n762), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT92), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n762), .A2(new_n765), .A3(new_n767), .A4(KEYINPUT92), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n710), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT31), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n654), .A2(new_n719), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n762), .A2(new_n767), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT91), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n765), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(KEYINPUT91), .ZN(new_n778));
  OAI211_X1 g0578(.A(KEYINPUT31), .B(new_n710), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n757), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n738), .A2(new_n756), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n735), .B1(new_n781), .B2(G1), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT96), .ZN(G364));
  NAND2_X1  g0583(.A1(new_n204), .A2(G13), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G45), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n730), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n717), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(G330), .B2(new_n715), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n728), .A2(new_n250), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G355), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G116), .B2(new_n207), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n728), .A2(new_n245), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n259), .B2(new_n211), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n237), .A2(G45), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n212), .B1(G20), .B2(new_n307), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n788), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G179), .A2(G200), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n806), .A2(G20), .A3(new_n378), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n245), .B1(new_n808), .B2(G329), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n806), .A2(G190), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G20), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n809), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(G20), .A2(G179), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT98), .Z(new_n816));
  NOR2_X1   g0616(.A1(new_n266), .A2(G190), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g0618(.A(KEYINPUT33), .B(G317), .Z(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G190), .A2(G200), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n814), .B(new_n820), .C1(G311), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n336), .A2(G200), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT99), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G20), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G190), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n816), .A2(G190), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(G200), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G283), .A2(new_n828), .B1(new_n830), .B2(G322), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n827), .A2(new_n378), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n829), .A2(new_n266), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G303), .A2(new_n832), .B1(new_n833), .B2(G326), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n824), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n808), .A2(G159), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT32), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n250), .B(new_n837), .C1(G77), .C2(new_n823), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n828), .A2(G107), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n830), .A2(G58), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G87), .A2(new_n832), .B1(new_n833), .B2(G50), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n818), .A2(new_n366), .B1(new_n813), .B2(new_n534), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT100), .Z(new_n844));
  OAI21_X1  g0644(.A(new_n835), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n805), .B1(new_n845), .B2(new_n802), .ZN(new_n846));
  INV_X1    g0646(.A(new_n801), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n715), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n790), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  INV_X1    g0650(.A(KEYINPUT102), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n334), .A2(new_n337), .A3(new_n719), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n318), .A2(new_n719), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n340), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n851), .B(new_n852), .C1(new_n854), .C2(new_n699), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n340), .A2(new_n853), .B1(new_n334), .B2(new_n337), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n334), .A2(new_n337), .A3(new_n719), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT102), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n737), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n859), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n695), .A2(new_n719), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n780), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n788), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n802), .A2(new_n799), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n787), .B1(new_n311), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n245), .B1(new_n808), .B2(G311), .ZN(new_n869));
  XOR2_X1   g0669(.A(KEYINPUT101), .B(G283), .Z(new_n870));
  OAI221_X1 g0670(.A(new_n869), .B1(new_n813), .B2(new_n534), .C1(new_n818), .C2(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(G294), .A2(new_n830), .B1(new_n833), .B2(G303), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n828), .A2(G87), .ZN(new_n873));
  INV_X1    g0673(.A(new_n832), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n872), .B(new_n873), .C1(new_n320), .C2(new_n874), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n871), .B(new_n875), .C1(G116), .C2(new_n823), .ZN(new_n876));
  INV_X1    g0676(.A(new_n818), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G150), .A2(new_n877), .B1(new_n823), .B2(G159), .ZN(new_n878));
  INV_X1    g0678(.A(new_n830), .ZN(new_n879));
  INV_X1    g0679(.A(G143), .ZN(new_n880));
  INV_X1    g0680(.A(G137), .ZN(new_n881));
  INV_X1    g0681(.A(new_n833), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n878), .B1(new_n879), .B2(new_n880), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT34), .ZN(new_n884));
  INV_X1    g0684(.A(G132), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n245), .B1(new_n885), .B2(new_n807), .C1(new_n813), .C2(new_n286), .ZN(new_n886));
  INV_X1    g0686(.A(new_n828), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(new_n366), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n886), .B(new_n888), .C1(G50), .C2(new_n832), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n876), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n802), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n868), .B1(new_n890), .B2(new_n891), .C1(new_n861), .C2(new_n800), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n866), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(G384));
  OR2_X1    g0694(.A1(new_n647), .A2(KEYINPUT35), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n647), .A2(KEYINPUT35), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n895), .A2(G116), .A3(new_n213), .A4(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT36), .Z(new_n898));
  OAI211_X1 g0698(.A(new_n211), .B(G77), .C1(new_n286), .C2(new_n366), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n277), .A2(G68), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n203), .B(G13), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n772), .A2(new_n773), .ZN(new_n903));
  INV_X1    g0703(.A(new_n573), .ZN(new_n904));
  INV_X1    g0704(.A(new_n609), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n660), .A4(new_n719), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n770), .A2(KEYINPUT31), .A3(new_n710), .A4(new_n771), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n903), .A2(new_n906), .A3(new_n910), .A4(new_n907), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n478), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT105), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n392), .A2(new_n710), .ZN(new_n915));
  INV_X1    g0715(.A(new_n390), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n916), .A2(new_n384), .A3(new_n388), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n383), .B(new_n915), .C1(new_n917), .C2(new_n376), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n377), .A2(new_n382), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n392), .B(new_n710), .C1(new_n391), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n861), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n910), .B1(new_n774), .B2(new_n907), .ZN(new_n924));
  INV_X1    g0724(.A(new_n911), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n708), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n451), .B2(new_n437), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n452), .B(KEYINPUT18), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n930), .B2(new_n466), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n461), .A2(new_n452), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT37), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT37), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n461), .A2(new_n452), .A3(new_n928), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  AND4_X1   g0737(.A1(new_n934), .A2(new_n461), .A3(new_n452), .A4(new_n928), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n272), .B1(new_n432), .B2(KEYINPUT16), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n450), .B2(new_n429), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n927), .B1(new_n940), .B2(new_n436), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n404), .B1(new_n940), .B2(new_n436), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n942), .A3(new_n461), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n938), .B1(KEYINPUT37), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n941), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n944), .B1(new_n468), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n937), .B1(new_n946), .B2(KEYINPUT38), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT40), .B1(new_n926), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT38), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n941), .B1(new_n457), .B2(new_n467), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(new_n944), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n943), .A2(KEYINPUT37), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n935), .ZN(new_n953));
  OAI211_X1 g0753(.A(KEYINPUT38), .B(new_n953), .C1(new_n476), .C2(new_n941), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT40), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n922), .B1(new_n909), .B2(new_n911), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n948), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n757), .B1(new_n914), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n914), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n478), .B1(new_n756), .B2(new_n738), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n703), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n951), .A2(new_n954), .A3(KEYINPUT39), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n393), .A2(new_n710), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n947), .C2(KEYINPUT39), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n951), .A2(new_n954), .ZN(new_n966));
  AOI211_X1 g0766(.A(KEYINPUT103), .B(new_n857), .C1(new_n736), .C2(new_n861), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT103), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n862), .B2(new_n852), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n966), .B(new_n921), .C1(new_n967), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n930), .A2(new_n708), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n962), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n960), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n203), .B2(new_n785), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n960), .A2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n902), .B1(new_n975), .B2(new_n976), .ZN(G367));
  INV_X1    g0777(.A(KEYINPUT106), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n741), .A2(new_n743), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n638), .A2(new_n710), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n682), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n710), .B1(new_n981), .B2(new_n642), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n642), .A2(new_n719), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n725), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n982), .B1(new_n986), .B2(KEYINPUT42), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(KEYINPUT42), .B2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n667), .A2(new_n710), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n677), .A2(new_n679), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n690), .B2(new_n989), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n978), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n988), .A2(new_n978), .A3(new_n992), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n995), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n722), .A2(new_n984), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n997), .B2(new_n998), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n729), .B(KEYINPUT41), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n984), .B1(new_n725), .B2(new_n718), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT44), .Z(new_n1005));
  NOR3_X1   g0805(.A1(new_n725), .A2(new_n984), .A3(new_n718), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT45), .ZN(new_n1007));
  AND3_X1   g0807(.A1(new_n1005), .A2(new_n722), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n722), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n724), .B(new_n721), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(KEYINPUT107), .B2(new_n716), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n716), .B(KEYINPUT107), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n781), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT108), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(KEYINPUT108), .A3(new_n781), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1010), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1003), .B1(new_n1019), .B2(new_n781), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n786), .A2(G1), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1001), .B(new_n1002), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n832), .A2(G116), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT46), .Z(new_n1024));
  AOI22_X1  g0824(.A1(G303), .A2(new_n830), .B1(new_n833), .B2(G311), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n534), .B2(new_n887), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n822), .A2(new_n870), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n245), .B1(new_n808), .B2(G317), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n813), .B2(new_n320), .C1(new_n818), .C2(new_n810), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT110), .Z(new_n1031));
  NAND2_X1  g0831(.A1(new_n812), .A2(G68), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n879), .B2(new_n279), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT111), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n245), .B1(new_n881), .B2(new_n807), .C1(new_n822), .C2(new_n277), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G159), .B2(new_n877), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n286), .A2(new_n874), .B1(new_n887), .B2(new_n311), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G143), .B2(new_n833), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT47), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT47), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n802), .A3(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n803), .B1(new_n207), .B2(new_n315), .C1(new_n795), .C2(new_n233), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n788), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT109), .Z(new_n1046));
  OAI211_X1 g0846(.A(new_n1043), .B(new_n1046), .C1(new_n847), .C2(new_n991), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1022), .A2(new_n1047), .ZN(G387));
  NOR2_X1   g0848(.A1(new_n721), .A2(new_n847), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n230), .A2(new_n259), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1050), .A2(new_n794), .B1(new_n732), .B2(new_n791), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n290), .A2(new_n277), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n259), .B1(new_n366), .B2(new_n311), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(new_n732), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n320), .B2(new_n728), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n788), .B1(new_n1058), .B2(new_n804), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G77), .A2(new_n832), .B1(new_n828), .B2(G97), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G50), .A2(new_n830), .B1(new_n833), .B2(G159), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n877), .A2(new_n290), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n245), .B1(new_n279), .B2(new_n807), .C1(new_n813), .C2(new_n315), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n823), .B2(G68), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n245), .B1(new_n808), .B2(G326), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n874), .A2(new_n810), .B1(new_n813), .B2(new_n870), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G303), .A2(new_n823), .B1(new_n877), .B2(G311), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n830), .A2(G317), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n833), .A2(G322), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1067), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1066), .B1(new_n579), .B2(new_n887), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1065), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1049), .B(new_n1059), .C1(new_n802), .C2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1015), .A2(new_n729), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1014), .A2(new_n781), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(G393));
  NAND2_X1  g0883(.A1(new_n794), .A2(new_n240), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n804), .B1(G97), .B2(new_n728), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n787), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n245), .B1(new_n808), .B2(G322), .ZN(new_n1087));
  INV_X1    g0887(.A(G303), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1087), .B1(new_n813), .B2(new_n579), .C1(new_n818), .C2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n839), .B1(new_n874), .B2(new_n870), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G294), .C2(new_n823), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G311), .A2(new_n830), .B1(new_n833), .B2(G317), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT52), .Z(new_n1093));
  AOI22_X1  g0893(.A1(G150), .A2(new_n833), .B1(new_n830), .B2(G159), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT51), .Z(new_n1095));
  OAI22_X1  g0895(.A1(new_n277), .A2(new_n818), .B1(new_n822), .B2(new_n316), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT113), .Z(new_n1097));
  OAI21_X1  g0897(.A(new_n245), .B1(new_n807), .B2(new_n880), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G77), .B2(new_n812), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n873), .B(new_n1099), .C1(new_n874), .C2(new_n366), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1091), .A2(new_n1093), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1086), .B1(new_n891), .B2(new_n1102), .C1(new_n985), .C2(new_n847), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1010), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1021), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n733), .B1(new_n1104), .B2(new_n1015), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1019), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(G390));
  NAND3_X1  g0909(.A1(new_n478), .A2(G330), .A3(new_n912), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n961), .A2(new_n1110), .A3(new_n703), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n755), .A2(new_n719), .A3(new_n861), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n852), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT114), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(KEYINPUT114), .A3(new_n852), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n757), .B(new_n859), .C1(new_n909), .C2(new_n911), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT115), .B1(new_n1118), .B2(new_n921), .ZN(new_n1119));
  OAI211_X1 g0919(.A(G330), .B(new_n861), .C1(new_n924), .C2(new_n925), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT115), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n918), .A2(new_n920), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n780), .A2(new_n861), .A3(new_n921), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1117), .A2(new_n1119), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1122), .B1(new_n864), .B2(new_n859), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n912), .A2(G330), .A3(new_n923), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n862), .A2(new_n968), .A3(new_n852), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n710), .B(new_n859), .C1(new_n687), .C2(new_n694), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT103), .B1(new_n1129), .B2(new_n857), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1126), .A2(new_n1127), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1111), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n963), .B1(new_n947), .B2(KEYINPUT39), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1122), .B1(new_n1130), .B2(new_n1128), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n964), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1112), .A2(KEYINPUT114), .A3(new_n852), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT114), .B1(new_n1112), .B2(new_n852), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n1122), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n947), .A2(new_n964), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1127), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1136), .B(new_n1124), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1133), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT116), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1146), .A2(new_n1147), .A3(new_n729), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n1146), .B2(new_n729), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1133), .B1(new_n1145), .B2(new_n1144), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT118), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1144), .A2(new_n1021), .A3(new_n1145), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1134), .A2(new_n799), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n787), .B1(new_n316), .B2(new_n867), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n888), .B1(G87), .B2(new_n832), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n245), .B1(new_n808), .B2(G294), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n813), .B2(new_n311), .C1(new_n822), .C2(new_n534), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G107), .B2(new_n877), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G116), .A2(new_n830), .B1(new_n833), .B2(G283), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1156), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1161), .A2(KEYINPUT117), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1163), .A2(new_n882), .B1(new_n879), .B2(new_n885), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G50), .B2(new_n828), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n832), .A2(G150), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT53), .Z(new_n1167));
  AOI21_X1  g0967(.A(new_n250), .B1(new_n808), .B2(G125), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n813), .B2(new_n414), .C1(new_n818), .C2(new_n881), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT54), .B(G143), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n823), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1165), .A2(new_n1167), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1162), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(KEYINPUT117), .B2(new_n1161), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1154), .B(new_n1155), .C1(new_n891), .C2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1152), .B1(new_n1153), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1153), .A2(new_n1152), .A3(new_n1176), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT119), .B1(new_n1151), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n921), .B1(new_n967), .B2(new_n969), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n964), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1115), .A2(new_n921), .A3(new_n1116), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1134), .A2(new_n1184), .B1(new_n1185), .B2(new_n1140), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1145), .B1(new_n1186), .B2(new_n1127), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1111), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1124), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1121), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1188), .B1(new_n1192), .B2(new_n1131), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n729), .B1(new_n1187), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT116), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1146), .A2(new_n1147), .A3(new_n729), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1150), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT119), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1153), .A2(new_n1152), .A3(new_n1176), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(new_n1177), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1181), .A2(new_n1202), .ZN(G378));
  INV_X1    g1003(.A(KEYINPUT122), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n306), .A2(new_n309), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n293), .A2(new_n927), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1207), .B(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n928), .B1(new_n467), .B2(new_n698), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n936), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n949), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n954), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n956), .A2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1215), .A2(KEYINPUT40), .B1(new_n955), .B2(new_n956), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1210), .B1(new_n1216), .B2(new_n757), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n965), .A2(new_n970), .A3(new_n971), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1210), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n955), .A2(new_n956), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT40), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n956), .B2(new_n1214), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G330), .B(new_n1219), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1217), .A2(new_n1218), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1218), .B1(new_n1217), .B2(new_n1223), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1204), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1219), .B1(new_n958), .B2(G330), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n757), .B(new_n1210), .C1(new_n948), .C2(new_n957), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n972), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1217), .A2(new_n1218), .A3(new_n1223), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(KEYINPUT122), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1226), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1210), .A2(new_n799), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n277), .B1(G33), .B2(G41), .C1(new_n328), .C2(new_n245), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n245), .B(new_n328), .C1(new_n808), .C2(G283), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1235), .A2(new_n1032), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n534), .B2(new_n818), .C1(new_n315), .C2(new_n822), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n828), .A2(G58), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n874), .B2(new_n311), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n320), .A2(new_n879), .B1(new_n882), .B2(new_n579), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1237), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1234), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT121), .Z(new_n1245));
  OAI22_X1  g1045(.A1(new_n818), .A2(new_n885), .B1(new_n813), .B2(new_n279), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G137), .B2(new_n823), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G125), .A2(new_n833), .B1(new_n830), .B2(G128), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n874), .C2(new_n1170), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(KEYINPUT59), .ZN(new_n1250));
  AOI211_X1 g1050(.A(G33), .B(G41), .C1(new_n808), .C2(G124), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n887), .B2(new_n414), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1249), .B2(KEYINPUT59), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1250), .A2(new_n1253), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n891), .B1(new_n1245), .B2(new_n1254), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n787), .B(new_n1255), .C1(new_n277), .C2(new_n867), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1232), .A2(new_n1021), .B1(new_n1233), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1188), .B1(new_n1187), .B2(new_n1193), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1225), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1229), .A2(KEYINPUT123), .A3(new_n1230), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1258), .A2(KEYINPUT57), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n729), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT57), .B1(new_n1232), .B2(new_n1258), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1257), .B1(new_n1263), .B2(new_n1264), .ZN(G375));
  OAI21_X1  g1065(.A(new_n1021), .B1(new_n1192), .B2(new_n1131), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G77), .A2(new_n828), .B1(new_n832), .B2(G97), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G283), .A2(new_n830), .B1(new_n833), .B2(G294), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n877), .A2(G116), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n250), .B1(new_n1088), .B2(new_n807), .C1(new_n813), .C2(new_n315), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n823), .B2(G107), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n245), .B1(new_n1163), .B2(new_n807), .C1(new_n813), .C2(new_n277), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n823), .B2(G150), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1274), .A2(new_n1238), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n833), .A2(G132), .B1(new_n877), .B2(new_n1171), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n881), .B2(new_n879), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1275), .B1(new_n414), .B2(new_n874), .C1(new_n1277), .C2(KEYINPUT124), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1277), .A2(KEYINPUT124), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1272), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n802), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n787), .B1(new_n366), .B2(new_n867), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1281), .B(new_n1282), .C1(new_n921), .C2(new_n800), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1266), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1003), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1125), .A2(new_n1132), .A3(new_n1111), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1193), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(G381));
  NOR3_X1   g1089(.A1(new_n1224), .A2(new_n1225), .A3(new_n1204), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT122), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1021), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1233), .A2(new_n1256), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1232), .A2(new_n1258), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT57), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1261), .A2(new_n1260), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1296), .B1(new_n1146), .B2(new_n1188), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n733), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1294), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1022), .A2(new_n1047), .A3(new_n1108), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1153), .A2(new_n1176), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1150), .B1(new_n1194), .B2(KEYINPUT116), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(new_n1196), .ZN(new_n1306));
  OR2_X1    g1106(.A1(G393), .A2(G396), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(G381), .A2(G384), .A3(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1301), .A2(new_n1303), .A3(new_n1306), .A4(new_n1308), .ZN(G407));
  INV_X1    g1109(.A(G213), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(G343), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1301), .A2(new_n1306), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(G407), .A2(G213), .A3(new_n1312), .ZN(G409));
  INV_X1    g1113(.A(new_n1311), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1287), .A2(KEYINPUT60), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT60), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1125), .A2(new_n1316), .A3(new_n1111), .A4(new_n1132), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1133), .A2(new_n733), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n893), .B(new_n1284), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1321));
  AOI21_X1  g1121(.A(G384), .B1(new_n1321), .B2(new_n1285), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G375), .B1(new_n1181), .B2(new_n1202), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1232), .A2(new_n1286), .A3(new_n1258), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1261), .A2(new_n1021), .A3(new_n1260), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1325), .A2(new_n1293), .A3(new_n1326), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1327), .A2(new_n1306), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1314), .B(new_n1323), .C1(new_n1324), .C2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT62), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1321), .A2(new_n1285), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n893), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1321), .A2(G384), .A3(new_n1285), .ZN(new_n1334));
  INV_X1    g1134(.A(G2897), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1314), .A2(new_n1335), .ZN(new_n1336));
  AND4_X1   g1136(.A1(KEYINPUT125), .A2(new_n1333), .A3(new_n1334), .A4(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1333), .A2(KEYINPUT125), .A3(new_n1334), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT125), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1340), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1339), .B(new_n1341), .C1(new_n1335), .C2(new_n1314), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1338), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1328), .B1(G378), .B2(new_n1301), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1343), .B1(new_n1344), .B2(new_n1311), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1199), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1301), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1327), .A2(new_n1306), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT62), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1350), .A2(new_n1351), .A3(new_n1314), .A4(new_n1323), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1330), .A2(new_n1331), .A3(new_n1345), .A4(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT127), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G393), .A2(G396), .ZN(new_n1355));
  AND3_X1   g1155(.A1(new_n1307), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1354), .B1(new_n1307), .B2(new_n1355), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1108), .B1(new_n1022), .B2(new_n1047), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1358), .B1(new_n1360), .B2(new_n1302), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1358), .ZN(new_n1362));
  NOR3_X1   g1162(.A1(new_n1303), .A2(new_n1359), .A3(new_n1362), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1361), .A2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1353), .A2(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1311), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1336), .B1(new_n1323), .B2(KEYINPUT125), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1337), .B1(new_n1367), .B2(new_n1341), .ZN(new_n1368));
  OAI21_X1  g1168(.A(KEYINPUT126), .B1(new_n1366), .B2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(KEYINPUT126), .ZN(new_n1370));
  OAI211_X1 g1170(.A(new_n1370), .B(new_n1343), .C1(new_n1344), .C2(new_n1311), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1369), .A2(new_n1371), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1331), .B1(new_n1361), .B2(new_n1363), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1323), .ZN(new_n1374));
  AOI211_X1 g1174(.A(new_n1311), .B(new_n1374), .C1(new_n1348), .C2(new_n1349), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1373), .B1(new_n1375), .B2(KEYINPUT63), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT63), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1329), .A2(new_n1377), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1372), .A2(new_n1376), .A3(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1365), .A2(new_n1379), .ZN(G405));
  INV_X1    g1180(.A(new_n1306), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1348), .B1(new_n1301), .B2(new_n1381), .ZN(new_n1382));
  OR2_X1    g1182(.A1(new_n1382), .A2(new_n1323), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1382), .A2(new_n1323), .ZN(new_n1384));
  AND3_X1   g1184(.A1(new_n1383), .A2(new_n1364), .A3(new_n1384), .ZN(new_n1385));
  AOI21_X1  g1185(.A(new_n1364), .B1(new_n1383), .B2(new_n1384), .ZN(new_n1386));
  NOR2_X1   g1186(.A1(new_n1385), .A2(new_n1386), .ZN(G402));
endmodule


