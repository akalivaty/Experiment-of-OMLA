//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  AOI22_X1  g0005(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G97), .A2(G257), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G58), .A2(G232), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G50), .A2(G226), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR3_X1   g0016(.A1(new_n210), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G77), .A2(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  OAI21_X1  g0020(.A(KEYINPUT64), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR3_X1    g0021(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT64), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n217), .A2(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n221), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n220), .ZN(new_n230));
  INV_X1    g0030(.A(G58), .ZN(new_n231));
  INV_X1    g0031(.A(G68), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n224), .B(new_n228), .C1(new_n230), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n212), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT66), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT67), .B(G107), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  OR2_X1    g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G222), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G223), .A2(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n261), .B(new_n265), .C1(G77), .C2(new_n257), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n264), .A2(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G226), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n266), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G200), .ZN(new_n274));
  INV_X1    g0074(.A(G190), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n229), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR3_X1   g0080(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n278), .A2(new_n280), .B1(new_n281), .B2(new_n220), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n220), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n277), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT68), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n219), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n277), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n290), .B(G50), .C1(G1), .C2(new_n220), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G50), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT9), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n274), .B1(new_n275), .B2(new_n273), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n296), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n295), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n273), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G179), .B2(new_n273), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  OAI211_X1 g0113(.A(G226), .B(new_n258), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(G232), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G97), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT74), .A4(new_n316), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n265), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n269), .B1(new_n271), .B2(G238), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT13), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT76), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT75), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n323), .B2(KEYINPUT13), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT13), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n321), .A2(KEYINPUT75), .A3(new_n329), .A4(new_n322), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n321), .B2(new_n322), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT76), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n326), .A2(new_n328), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n333), .A2(new_n334), .A3(G169), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(new_n333), .B2(G169), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n321), .A2(new_n329), .A3(new_n322), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n331), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G179), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n335), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G13), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(G1), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT71), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(G20), .ZN(new_n345));
  INV_X1    g0145(.A(new_n277), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n288), .A2(KEYINPUT71), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(KEYINPUT73), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(new_n219), .B2(G20), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT12), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n345), .A2(new_n347), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n232), .A2(G20), .ZN(new_n357));
  INV_X1    g0157(.A(G77), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n357), .B1(new_n284), .B2(new_n358), .C1(new_n280), .C2(new_n293), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n277), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT11), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n288), .A2(new_n353), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n354), .A2(new_n356), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n333), .B2(G200), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT77), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n338), .B2(G190), .ZN(new_n367));
  NOR4_X1   g0167(.A1(new_n337), .A2(new_n331), .A3(KEYINPUT77), .A4(new_n275), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n365), .A2(KEYINPUT78), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT78), .B1(new_n365), .B2(new_n369), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n341), .A2(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT69), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n257), .A2(G238), .A3(G1698), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(new_n203), .C2(new_n257), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n265), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n271), .A2(G244), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n270), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G200), .ZN(new_n380));
  INV_X1    g0180(.A(new_n283), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n279), .B1(G20), .B2(G77), .ZN(new_n382));
  OR2_X1    g0182(.A1(KEYINPUT15), .A2(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT15), .A2(G87), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT70), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(KEYINPUT70), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n382), .B1(new_n389), .B2(new_n284), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n352), .A2(G77), .B1(new_n277), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n355), .A2(new_n358), .ZN(new_n392));
  XOR2_X1   g0192(.A(new_n392), .B(KEYINPUT72), .Z(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n380), .B(new_n395), .C1(new_n275), .C2(new_n379), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n379), .A2(new_n306), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n377), .A2(new_n398), .A3(new_n270), .A4(new_n378), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n394), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT17), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n257), .B2(G20), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n312), .A2(new_n313), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n232), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G58), .A2(G68), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n233), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G20), .ZN(new_n411));
  INV_X1    g0211(.A(G159), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n280), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n403), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n406), .B2(new_n220), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n312), .A2(new_n313), .A3(new_n404), .A4(G20), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n411), .B(KEYINPUT79), .C1(new_n412), .C2(new_n280), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT79), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n280), .A2(new_n412), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n220), .B1(new_n233), .B2(new_n409), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n418), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n414), .A2(new_n423), .A3(new_n277), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT80), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(G223), .B(new_n258), .C1(new_n312), .C2(new_n313), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT81), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n257), .A2(KEYINPUT81), .A3(G223), .A4(new_n258), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n257), .A2(G226), .A3(G1698), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n429), .A2(new_n430), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n269), .B1(new_n433), .B2(new_n265), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n271), .A2(G232), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(G190), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n283), .B1(new_n219), .B2(G20), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n290), .B1(new_n289), .B2(new_n283), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n414), .A2(new_n423), .A3(KEYINPUT80), .A4(new_n277), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n426), .A2(new_n436), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n433), .A2(new_n265), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n270), .A3(new_n435), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G200), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n402), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n426), .A2(new_n438), .A3(new_n439), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(KEYINPUT17), .A3(new_n443), .A4(new_n436), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(G169), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n434), .A2(G179), .A3(new_n435), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(KEYINPUT82), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT82), .B1(new_n449), .B2(new_n450), .ZN(new_n453));
  OAI211_X1 g0253(.A(KEYINPUT18), .B(new_n446), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT82), .ZN(new_n456));
  INV_X1    g0256(.A(new_n450), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n306), .B1(new_n434), .B2(new_n435), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n451), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT18), .B1(new_n460), .B2(new_n446), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n445), .B(new_n448), .C1(new_n455), .C2(new_n461), .ZN(new_n462));
  NOR4_X1   g0262(.A1(new_n311), .A2(new_n372), .A3(new_n401), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n264), .A2(G274), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n219), .B(G45), .C1(new_n263), .C2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT88), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n464), .ZN(new_n471));
  OAI211_X1 g0271(.A(G270), .B(new_n264), .C1(new_n471), .C2(new_n466), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n258), .A2(G257), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G264), .A2(G1698), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n476), .C1(new_n312), .C2(new_n313), .ZN(new_n477));
  INV_X1    g0277(.A(G303), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n255), .A2(new_n478), .A3(new_n256), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT90), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n477), .A2(KEYINPUT90), .A3(new_n479), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n265), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G200), .ZN(new_n486));
  AOI21_X1  g0286(.A(G20), .B1(new_n262), .B2(G97), .ZN(new_n487));
  AND3_X1   g0287(.A1(KEYINPUT86), .A2(G33), .A3(G283), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT86), .B1(G33), .B2(G283), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n276), .A2(new_n229), .B1(G20), .B2(new_n211), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT20), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n493), .A2(new_n494), .B1(new_n211), .B2(new_n355), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n350), .A2(new_n351), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n219), .A2(G33), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(G116), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n486), .A2(KEYINPUT91), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT91), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n495), .ZN(new_n501));
  INV_X1    g0301(.A(G200), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n474), .B2(new_n484), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n500), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n474), .A2(G190), .A3(new_n484), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n499), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n497), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n211), .B(new_n507), .C1(new_n350), .C2(new_n351), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n355), .A2(new_n211), .ZN(new_n509));
  INV_X1    g0309(.A(new_n494), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n492), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n485), .B(G169), .C1(new_n508), .C2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n485), .A2(new_n398), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n501), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n501), .A2(KEYINPUT21), .A3(G169), .A4(new_n485), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n506), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n220), .A2(G107), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n343), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n521), .A2(KEYINPUT25), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(KEYINPUT25), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n346), .A2(new_n288), .A3(new_n497), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n203), .C2(new_n524), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n525), .B(KEYINPUT93), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n220), .A2(G33), .A3(G116), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n520), .B(KEYINPUT23), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT22), .ZN(new_n529));
  AOI21_X1  g0329(.A(G20), .B1(new_n255), .B2(new_n256), .ZN(new_n530));
  OR2_X1    g0330(.A1(new_n214), .A2(KEYINPUT92), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n220), .B1(new_n312), .B2(new_n313), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n534), .A2(KEYINPUT22), .A3(new_n531), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n527), .B(new_n528), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n530), .A2(new_n532), .A3(new_n529), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT22), .B1(new_n534), .B2(new_n531), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n541), .A2(KEYINPUT24), .A3(new_n527), .A4(new_n528), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n277), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n468), .A2(new_n469), .ZN(new_n544));
  INV_X1    g0344(.A(new_n465), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n215), .A2(new_n258), .ZN(new_n547));
  OAI221_X1 g0347(.A(new_n547), .B1(G257), .B2(new_n258), .C1(new_n312), .C2(new_n313), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n265), .ZN(new_n551));
  OAI211_X1 g0351(.A(G264), .B(new_n264), .C1(new_n471), .C2(new_n466), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n264), .B1(new_n548), .B2(new_n549), .ZN(new_n555));
  INV_X1    g0355(.A(new_n552), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n470), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G190), .ZN(new_n558));
  AND4_X1   g0358(.A1(new_n526), .A2(new_n543), .A3(new_n554), .A4(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n546), .A2(new_n551), .A3(new_n398), .A4(new_n552), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n557), .B2(G169), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n526), .B2(new_n543), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT94), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT94), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n543), .A2(new_n526), .A3(new_n554), .A4(new_n558), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n543), .A2(new_n526), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n561), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n488), .A2(new_n489), .ZN(new_n569));
  OAI211_X1 g0369(.A(G250), .B(G1698), .C1(new_n312), .C2(new_n313), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n570), .A2(KEYINPUT87), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(KEYINPUT87), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n257), .A2(G244), .A3(new_n258), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT4), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n265), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n471), .A2(new_n466), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n265), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G257), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n546), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n306), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n289), .A2(new_n202), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n524), .B2(new_n202), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT84), .ZN(new_n588));
  NAND2_X1  g0388(.A1(KEYINPUT6), .A2(G97), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(G107), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n203), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(G97), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G97), .A2(G107), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT6), .B1(new_n204), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(G20), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n279), .A2(G77), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT83), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n595), .A2(new_n598), .A3(KEYINPUT85), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT85), .B1(new_n595), .B2(new_n598), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n203), .B1(new_n405), .B2(new_n407), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n587), .B1(new_n602), .B2(new_n346), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n579), .A2(new_n398), .A3(new_n546), .A4(new_n582), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n584), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n219), .A2(G45), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n268), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n257), .A2(G244), .A3(G1698), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G116), .ZN(new_n609));
  OAI211_X1 g0409(.A(G238), .B(new_n258), .C1(new_n312), .C2(new_n313), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n607), .B1(new_n611), .B2(new_n265), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n264), .A2(G250), .A3(new_n606), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT89), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT89), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n264), .A2(new_n615), .A3(G250), .A4(new_n606), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n612), .A2(G190), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n502), .B1(new_n612), .B2(new_n617), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n214), .A2(new_n202), .A3(new_n203), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n316), .A2(new_n220), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n622), .A3(KEYINPUT19), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT19), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n316), .B2(G20), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n623), .B(new_n625), .C1(new_n232), .C2(new_n534), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n277), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n389), .A2(new_n355), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n290), .A2(G87), .A3(new_n497), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n611), .A2(new_n265), .ZN(new_n631));
  INV_X1    g0431(.A(new_n607), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n631), .A2(new_n398), .A3(new_n632), .A4(new_n617), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n627), .B(new_n628), .C1(new_n389), .C2(new_n524), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n612), .A2(new_n617), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n306), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n620), .A2(new_n630), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n583), .A2(G200), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n595), .A2(new_n598), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT85), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n601), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n595), .A2(new_n598), .A3(KEYINPUT85), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n586), .B1(new_n645), .B2(new_n277), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n579), .A2(G190), .A3(new_n546), .A4(new_n582), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n639), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n605), .A2(new_n638), .A3(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n463), .A2(new_n519), .A3(new_n568), .A4(new_n649), .ZN(G372));
  NAND2_X1  g0450(.A1(new_n365), .A2(new_n369), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT78), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n365), .A2(new_n369), .A3(KEYINPUT78), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n400), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n336), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n333), .A2(new_n334), .A3(G169), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n339), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n363), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n445), .A3(new_n448), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n449), .A2(new_n450), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n446), .A2(KEYINPUT18), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT18), .B1(new_n446), .B2(new_n664), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n309), .B1(new_n668), .B2(new_n304), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n649), .A2(KEYINPUT95), .A3(new_n565), .ZN(new_n670));
  INV_X1    g0470(.A(new_n518), .ZN(new_n671));
  INV_X1    g0471(.A(new_n562), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT95), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n605), .A2(new_n638), .A3(new_n648), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n559), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n645), .A2(new_n277), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n678), .A2(new_n587), .B1(new_n583), .B2(new_n306), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n638), .A2(new_n679), .A3(KEYINPUT26), .A4(new_n604), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT96), .ZN(new_n681));
  INV_X1    g0481(.A(new_n605), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT96), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT26), .A4(new_n638), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  INV_X1    g0485(.A(new_n638), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(new_n605), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n635), .A2(new_n637), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n677), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n463), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n669), .A2(new_n692), .ZN(G369));
  NAND2_X1  g0493(.A1(new_n343), .A2(new_n220), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n695), .A2(new_n696), .A3(G213), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G343), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT97), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n501), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n519), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n671), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT98), .B(G330), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n566), .A2(new_n699), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n563), .B2(new_n567), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n562), .B2(new_n700), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n673), .B(new_n699), .C1(new_n568), .C2(new_n562), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n226), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n621), .A2(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n234), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n687), .A2(new_n680), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n689), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n673), .A2(new_n565), .A3(new_n649), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n699), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n691), .A2(new_n699), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(KEYINPUT29), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n636), .A2(new_n553), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n570), .B(KEYINPUT87), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n569), .A3(new_n576), .A4(new_n577), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n728), .A2(new_n265), .B1(G257), .B2(new_n581), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n515), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(G179), .B1(new_n612), .B2(new_n617), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n583), .A2(new_n485), .A3(new_n553), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT99), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n735), .A2(new_n736), .B1(new_n731), .B2(new_n730), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT99), .B1(new_n732), .B2(new_n734), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT31), .B(new_n700), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n730), .A2(new_n731), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n700), .B1(new_n735), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n568), .A2(new_n519), .A3(new_n649), .A4(new_n699), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n704), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n725), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n718), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n703), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(G355), .B(KEYINPUT100), .ZN(new_n755));
  INV_X1    g0555(.A(G45), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n249), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n406), .B1(new_n234), .B2(G45), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n226), .B1(new_n406), .B2(new_n755), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n220), .B1(KEYINPUT101), .B2(new_n306), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(KEYINPUT101), .B2(new_n306), .ZN(new_n761));
  INV_X1    g0561(.A(new_n229), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n752), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n759), .B(new_n765), .C1(new_n211), .C2(new_n226), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n398), .A2(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n220), .A2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n398), .A2(new_n502), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n769), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G317), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G179), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n769), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G329), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n502), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n769), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n781), .B(new_n785), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n220), .B1(new_n782), .B2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n774), .B(new_n789), .C1(G294), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n220), .A2(new_n275), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n768), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G322), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n793), .A2(new_n787), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G303), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n793), .A2(new_n775), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n257), .B1(new_n801), .B2(G326), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n792), .A2(new_n796), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n790), .A2(KEYINPUT102), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n790), .A2(KEYINPUT102), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n202), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n798), .A2(G87), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n777), .A2(G68), .ZN(new_n810));
  INV_X1    g0610(.A(new_n788), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G107), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT32), .B1(new_n783), .B2(new_n412), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n809), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n783), .A2(KEYINPUT32), .A3(new_n412), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n808), .A2(new_n814), .A3(new_n406), .A4(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n795), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n293), .B2(new_n800), .C1(new_n231), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n772), .A2(new_n358), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n803), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n764), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n342), .A2(G20), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n219), .B1(new_n822), .B2(G45), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n713), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n754), .A2(new_n766), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n703), .A2(new_n704), .ZN(new_n827));
  INV_X1    g0627(.A(new_n825), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n705), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT103), .Z(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n397), .A2(new_n399), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT105), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n700), .A2(new_n394), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n396), .A2(new_n400), .A3(new_n835), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n834), .B1(new_n833), .B2(new_n835), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n724), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n699), .B(new_n839), .C1(new_n677), .C2(new_n690), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(new_n747), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n828), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n788), .A2(new_n232), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n771), .A2(G159), .B1(new_n795), .B2(G143), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n848), .B2(new_n800), .C1(new_n278), .C2(new_n776), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT104), .B(KEYINPUT34), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n850), .B1(new_n293), .B2(new_n797), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n846), .B(new_n851), .C1(G58), .C2(new_n791), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n849), .A2(new_n850), .B1(G132), .B2(new_n784), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(new_n257), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n797), .A2(new_n203), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n855), .B(new_n808), .C1(G294), .C2(new_n795), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n811), .A2(G87), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n772), .A2(new_n211), .B1(new_n783), .B2(new_n773), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G283), .B2(new_n777), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n257), .B1(new_n801), .B2(G303), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n856), .A2(new_n857), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n763), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n764), .A2(new_n750), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n828), .B(new_n862), .C1(new_n358), .C2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n839), .B2(new_n751), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n845), .A2(new_n865), .ZN(G384));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n460), .A2(new_n446), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n440), .A2(new_n444), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n446), .A2(new_n697), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n418), .A2(new_n422), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n403), .B1(new_n874), .B2(new_n408), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n277), .A3(new_n423), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n438), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n664), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n440), .B2(new_n444), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT108), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT108), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n878), .B(new_n881), .C1(new_n440), .C2(new_n444), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n697), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n873), .B1(KEYINPUT37), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n883), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n462), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n867), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n889), .A2(new_n872), .B1(new_n462), .B2(new_n886), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(KEYINPUT31), .B(new_n700), .C1(new_n735), .C2(new_n740), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n744), .A2(new_n743), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n839), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n364), .A2(new_n699), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n372), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n661), .A2(new_n655), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT40), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT111), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT110), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT40), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n894), .A2(new_n839), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n372), .A2(new_n896), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n898), .B1(new_n661), .B2(new_n655), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n905), .B(new_n903), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n871), .B1(new_n444), .B2(new_n440), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n446), .A2(new_n664), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n872), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n448), .B(new_n445), .C1(new_n665), .C2(new_n666), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n914), .B2(new_n871), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n867), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n891), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n902), .B1(new_n904), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(KEYINPUT110), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n900), .A2(new_n903), .B1(new_n891), .B2(new_n916), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT111), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n901), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n463), .A2(new_n894), .ZN(new_n926));
  XNOR2_X1  g0726(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n925), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n704), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n897), .A2(new_n899), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n656), .A2(new_n699), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n842), .A2(KEYINPUT107), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT107), .B1(new_n842), .B2(new_n932), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n931), .B(new_n892), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n917), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n661), .A2(new_n700), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n888), .A2(new_n891), .A3(KEYINPUT39), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n667), .A2(new_n697), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n935), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT109), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n935), .A2(new_n940), .A3(new_n944), .A4(new_n941), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n930), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n725), .A2(new_n463), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n669), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n947), .B(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n219), .B2(new_n822), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n592), .A2(new_n594), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n211), .B1(new_n953), .B2(KEYINPUT35), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n954), .B(new_n230), .C1(KEYINPUT35), .C2(new_n953), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT36), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n232), .A2(KEYINPUT106), .A3(G50), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT106), .B1(new_n232), .B2(G50), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n409), .A2(G77), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n957), .B(new_n958), .C1(new_n234), .C2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n342), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n951), .A2(new_n956), .A3(new_n961), .ZN(G367));
  NAND2_X1  g0762(.A1(new_n226), .A2(new_n406), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n765), .B1(new_n226), .B2(new_n389), .C1(new_n244), .C2(new_n963), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n788), .A2(new_n202), .B1(new_n783), .B2(new_n778), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n406), .B1(new_n203), .B2(new_n790), .C1(new_n817), .C2(new_n478), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(G283), .C2(new_n771), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n798), .A2(G116), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT46), .ZN(new_n969));
  INV_X1    g0769(.A(G294), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n967), .B(new_n969), .C1(new_n970), .C2(new_n776), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G311), .B2(new_n801), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n795), .A2(G150), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n797), .A2(new_n231), .ZN(new_n974));
  INV_X1    g0774(.A(new_n807), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(G68), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n771), .A2(G50), .B1(new_n784), .B2(G137), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G159), .A2(new_n777), .B1(new_n811), .B2(G77), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n976), .A2(new_n257), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n974), .B(new_n979), .C1(G143), .C2(new_n801), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n972), .B1(new_n973), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT47), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n825), .B(new_n964), .C1(new_n982), .C2(new_n763), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n699), .A2(new_n630), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n638), .B(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n983), .B1(new_n752), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n648), .B1(new_n646), .B2(new_n699), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(new_n682), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n671), .A2(new_n700), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n707), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n605), .B1(new_n988), .B2(new_n672), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n991), .A2(KEYINPUT42), .B1(new_n699), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT114), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(KEYINPUT42), .B2(new_n991), .ZN(new_n995));
  INV_X1    g0795(.A(new_n985), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n709), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n682), .A2(new_n700), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n682), .B2(new_n988), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n998), .A2(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1007), .B(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n705), .B(new_n708), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(new_n990), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n748), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n710), .A2(new_n989), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(KEYINPUT116), .B(KEYINPUT44), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n710), .A2(new_n1001), .ZN(new_n1017));
  XOR2_X1   g0817(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  OR3_X1    g0820(.A1(new_n1020), .A2(KEYINPUT117), .A3(new_n709), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1020), .B1(KEYINPUT117), .B2(new_n709), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1013), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n748), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n713), .B(KEYINPUT41), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n824), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n987), .B1(new_n1010), .B2(new_n1026), .ZN(G387));
  NOR2_X1   g0827(.A1(new_n748), .A2(new_n1012), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1013), .B1(KEYINPUT118), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n713), .C1(KEYINPUT118), .C2(new_n1028), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1012), .A2(new_n824), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G322), .A2(new_n801), .B1(new_n777), .B2(G311), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n478), .B2(new_n772), .C1(new_n778), .C2(new_n817), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT48), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n786), .B2(new_n790), .C1(new_n970), .C2(new_n797), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n784), .A2(G326), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n257), .B1(new_n811), .B2(G116), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n807), .A2(new_n389), .B1(new_n278), .B2(new_n783), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n817), .A2(new_n293), .B1(new_n788), .B2(new_n202), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n257), .B1(new_n776), .B2(new_n283), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n797), .A2(new_n358), .ZN(new_n1043));
  NOR4_X1   g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n232), .B2(new_n772), .C1(new_n412), .C2(new_n800), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n763), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n241), .A2(new_n756), .A3(new_n257), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT50), .B1(new_n283), .B2(G50), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(G68), .A2(G77), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n756), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n406), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1047), .B1(new_n715), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n765), .B1(new_n1053), .B2(new_n712), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G107), .B2(new_n712), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1046), .A2(new_n828), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n708), .A2(new_n752), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1030), .A2(new_n1031), .A3(new_n1058), .ZN(G393));
  XNOR2_X1  g0859(.A(new_n1020), .B(new_n999), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1023), .B(new_n713), .C1(new_n1013), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n824), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n795), .A2(G159), .B1(new_n801), .B2(G150), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G143), .B2(new_n784), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n975), .A2(G77), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n771), .A2(new_n381), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n857), .B1(new_n293), .B2(new_n776), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n406), .B(new_n1068), .C1(G68), .C2(new_n798), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n776), .A2(new_n478), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n817), .A2(new_n773), .B1(new_n778), .B2(new_n800), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n798), .A2(G283), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n812), .B1(new_n772), .B2(new_n970), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G116), .B2(new_n791), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n257), .B1(new_n784), .B2(G322), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1070), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n828), .B1(new_n1079), .B2(new_n764), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n765), .B1(new_n202), .B2(new_n226), .C1(new_n253), .C2(new_n963), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n1001), .C2(new_n753), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1062), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1061), .A2(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(KEYINPUT119), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n931), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n842), .A2(new_n932), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT107), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n842), .A2(KEYINPUT107), .A3(new_n932), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1085), .B1(new_n1091), .B2(new_n938), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n937), .A2(new_n939), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n938), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(KEYINPUT119), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1092), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n722), .A2(new_n840), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n656), .B2(new_n699), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1095), .B(new_n917), .C1(new_n1099), .C2(new_n1086), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n747), .A2(new_n931), .A3(new_n839), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1097), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n931), .A2(G330), .A3(new_n905), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n824), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1093), .A2(new_n750), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1066), .B1(new_n211), .B2(new_n817), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT121), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n777), .A2(G107), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n809), .B1(new_n783), .B2(new_n970), .C1(new_n786), .C2(new_n800), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n846), .B(new_n1112), .C1(G97), .C2(new_n771), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1110), .A2(new_n406), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(G132), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n817), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n797), .A2(new_n278), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1118));
  XNOR2_X1  g0918(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G137), .A2(new_n777), .B1(new_n784), .B2(G125), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(new_n412), .C2(new_n807), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n801), .A2(G128), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT54), .B(G143), .Z(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n257), .B1(new_n293), .B2(new_n788), .C1(new_n772), .C2(new_n1124), .ZN(new_n1125));
  OR4_X1    g0925(.A1(new_n1116), .A2(new_n1121), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n763), .B1(new_n1114), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n828), .B(new_n1127), .C1(new_n283), .C2(new_n863), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1108), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1107), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1104), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1131), .B2(new_n1101), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n463), .A2(G330), .A3(new_n894), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n948), .A2(new_n669), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n931), .B1(new_n747), .B2(new_n839), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1105), .A2(new_n1137), .B1(new_n934), .B2(new_n933), .ZN(new_n1138));
  INV_X1    g0938(.A(G330), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1086), .B1(new_n1139), .B2(new_n895), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1133), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n714), .B1(new_n1133), .B2(new_n1144), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1130), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(G378));
  INV_X1    g0948(.A(KEYINPUT123), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n943), .A2(new_n945), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n919), .A2(new_n924), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n901), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n311), .A2(KEYINPUT55), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT55), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n304), .A2(new_n1154), .A3(new_n310), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n697), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n305), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1153), .A2(new_n1155), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1154), .B1(new_n304), .B2(new_n310), .ZN(new_n1160));
  AOI211_X1 g0960(.A(KEYINPUT55), .B(new_n309), .C1(new_n301), .C2(new_n303), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AND4_X1   g0966(.A1(G330), .A2(new_n1151), .A3(new_n1152), .A4(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n925), .B2(G330), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1150), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1151), .A2(G330), .A3(new_n1152), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1166), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n925), .A2(G330), .A3(new_n1166), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n946), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1149), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT123), .B1(new_n1176), .B2(new_n1150), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n824), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n293), .B1(new_n312), .B2(G41), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n975), .A2(G150), .B1(G137), .B2(new_n771), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G125), .A2(new_n801), .B1(new_n777), .B2(G132), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n797), .C2(new_n1124), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G128), .B2(new_n795), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT59), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G33), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G41), .B1(new_n784), .B2(G124), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n412), .C2(new_n788), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1179), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n976), .B1(new_n203), .B2(new_n817), .C1(new_n389), .C2(new_n772), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G97), .B2(new_n777), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n800), .A2(new_n211), .B1(new_n788), .B2(new_n231), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n406), .B1(new_n783), .B2(new_n786), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1192), .A2(new_n1043), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n263), .A3(new_n1194), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT58), .Z(new_n1196));
  OAI21_X1  g0996(.A(new_n764), .B1(new_n1189), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n828), .B1(new_n293), .B2(new_n863), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n1166), .C2(new_n751), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1178), .A2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1172), .A2(new_n946), .A3(new_n1173), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n946), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1202));
  OAI21_X1  g1002(.A(KEYINPUT123), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1177), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1144), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1136), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT57), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(KEYINPUT57), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n713), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1200), .B1(new_n1208), .B2(new_n1211), .ZN(G375));
  AOI21_X1  g1012(.A(new_n406), .B1(new_n795), .B2(G137), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n1115), .B2(new_n800), .C1(new_n412), .C2(new_n797), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G50), .B2(new_n975), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G58), .A2(new_n811), .B1(new_n784), .B2(G128), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n776), .C2(new_n1124), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G150), .B2(new_n771), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n389), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n975), .A2(new_n1219), .B1(G283), .B2(new_n795), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n257), .B1(new_n777), .B2(G116), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n478), .C2(new_n783), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n772), .A2(new_n203), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n797), .A2(new_n202), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n800), .A2(new_n970), .B1(new_n788), .B2(new_n358), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n764), .B1(new_n1218), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n863), .A2(new_n232), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n825), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1086), .B2(new_n750), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1142), .B2(new_n824), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1135), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1025), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1231), .B1(new_n1144), .B2(new_n1233), .ZN(G381));
  NAND2_X1  g1034(.A1(new_n1178), .A2(new_n1199), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1207), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT57), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1206), .A2(new_n1136), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n714), .B1(new_n1239), .B2(KEYINPUT57), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1235), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1147), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1030), .A2(new_n831), .A3(new_n1031), .A4(new_n1058), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1242), .A2(G390), .A3(new_n1243), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(G387), .A2(G381), .A3(G384), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(G407));
  INV_X1    g1046(.A(G343), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(G213), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT124), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(new_n1242), .C2(new_n1250), .ZN(G409));
  NAND3_X1  g1051(.A1(new_n1205), .A2(new_n1025), .A3(new_n1207), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1209), .A2(new_n824), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n1147), .A3(new_n1199), .A4(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1250), .B(new_n1254), .C1(new_n1241), .C2(new_n1147), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1232), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1232), .A2(new_n1256), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(new_n713), .A3(new_n1143), .A4(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(G384), .A3(new_n1231), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G384), .B1(new_n1259), .B2(new_n1231), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT62), .B1(new_n1255), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1249), .A2(G2897), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(G2897), .A3(new_n1249), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1255), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1249), .B1(G375), .B2(G378), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1263), .A4(new_n1254), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1265), .A2(new_n1270), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(G390), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G387), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1243), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(KEYINPUT126), .A3(new_n1243), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n987), .B(G390), .C1(new_n1010), .C2(new_n1026), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G387), .A2(new_n1275), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1284), .A2(KEYINPUT127), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1285), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1274), .A2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1293), .A2(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1255), .B2(new_n1264), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1271), .A2(KEYINPUT63), .A3(new_n1263), .A4(new_n1254), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1269), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n1268), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1255), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1294), .A2(new_n1296), .A3(new_n1297), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1292), .A2(new_n1302), .ZN(G405));
  NAND2_X1  g1103(.A1(G375), .A2(G378), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1242), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1263), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1242), .A3(new_n1264), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1306), .A2(new_n1293), .A3(new_n1307), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


