

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U324 ( .A(n432), .B(KEYINPUT55), .ZN(n433) );
  XNOR2_X1 U325 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U326 ( .A(n356), .B(n399), .Z(n291) );
  XNOR2_X1 U327 ( .A(n387), .B(KEYINPUT45), .ZN(n388) );
  XNOR2_X1 U328 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U329 ( .A(KEYINPUT107), .B(KEYINPUT47), .ZN(n384) );
  XNOR2_X1 U330 ( .A(n385), .B(n384), .ZN(n393) );
  INV_X1 U331 ( .A(KEYINPUT32), .ZN(n343) );
  XNOR2_X1 U332 ( .A(n344), .B(n343), .ZN(n345) );
  NOR2_X1 U333 ( .A1(n507), .A2(n411), .ZN(n564) );
  XNOR2_X1 U334 ( .A(n395), .B(n394), .ZN(n538) );
  XNOR2_X1 U335 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U336 ( .A(n434), .B(n433), .ZN(n449) );
  XNOR2_X1 U337 ( .A(KEYINPUT122), .B(n565), .ZN(n577) );
  XNOR2_X1 U338 ( .A(n448), .B(n447), .ZN(n522) );
  XNOR2_X1 U339 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n450) );
  XNOR2_X1 U340 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(G57GAT), .B(G155GAT), .Z(n293) );
  XNOR2_X1 U342 ( .A(G148GAT), .B(G162GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n295) );
  XOR2_X1 U344 ( .A(G29GAT), .B(G85GAT), .Z(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n312) );
  XOR2_X1 U346 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n297) );
  XNOR2_X1 U347 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U349 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n299) );
  XNOR2_X1 U350 ( .A(KEYINPUT86), .B(KEYINPUT1), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(n301), .B(n300), .Z(n310) );
  XNOR2_X1 U353 ( .A(G127GAT), .B(G134GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n302), .B(KEYINPUT76), .ZN(n303) );
  XOR2_X1 U355 ( .A(n303), .B(KEYINPUT0), .Z(n305) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(G120GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n448) );
  XOR2_X1 U358 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n307) );
  XNOR2_X1 U359 ( .A(KEYINPUT3), .B(KEYINPUT83), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U361 ( .A(G141GAT), .B(n308), .Z(n431) );
  XNOR2_X1 U362 ( .A(n448), .B(n431), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n314) );
  NAND2_X1 U365 ( .A1(G225GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n507) );
  XOR2_X1 U367 ( .A(G29GAT), .B(G43GAT), .Z(n316) );
  XNOR2_X1 U368 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n360) );
  XOR2_X1 U370 ( .A(G15GAT), .B(G1GAT), .Z(n377) );
  XOR2_X1 U371 ( .A(n360), .B(n377), .Z(n318) );
  NAND2_X1 U372 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U374 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n320) );
  XNOR2_X1 U375 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U377 ( .A(n322), .B(n321), .Z(n330) );
  XOR2_X1 U378 ( .A(G113GAT), .B(G50GAT), .Z(n324) );
  XNOR2_X1 U379 ( .A(G169GAT), .B(G36GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U381 ( .A(G8GAT), .B(G141GAT), .Z(n326) );
  XNOR2_X1 U382 ( .A(G22GAT), .B(G197GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n566) );
  XOR2_X1 U386 ( .A(KEYINPUT13), .B(KEYINPUT68), .Z(n332) );
  XNOR2_X1 U387 ( .A(G71GAT), .B(G78GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U389 ( .A(G57GAT), .B(n333), .ZN(n380) );
  INV_X1 U390 ( .A(n380), .ZN(n337) );
  XOR2_X1 U391 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n335) );
  XNOR2_X1 U392 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n337), .B(n336), .ZN(n348) );
  XOR2_X1 U395 ( .A(G64GAT), .B(G92GAT), .Z(n339) );
  XNOR2_X1 U396 ( .A(G176GAT), .B(G204GAT), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n400) );
  XOR2_X1 U398 ( .A(G99GAT), .B(G85GAT), .Z(n356) );
  XNOR2_X1 U399 ( .A(n400), .B(n356), .ZN(n341) );
  AND2_X1 U400 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n346) );
  XNOR2_X1 U402 ( .A(G106GAT), .B(KEYINPUT69), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n342), .B(G148GAT), .ZN(n423) );
  XNOR2_X1 U404 ( .A(n423), .B(KEYINPUT31), .ZN(n344) );
  XOR2_X1 U405 ( .A(n348), .B(n347), .Z(n571) );
  INV_X1 U406 ( .A(KEYINPUT65), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n571), .B(n349), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n350), .B(KEYINPUT41), .ZN(n552) );
  NOR2_X1 U409 ( .A1(n566), .A2(n552), .ZN(n352) );
  INV_X1 U410 ( .A(KEYINPUT46), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n383) );
  XOR2_X1 U412 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n354) );
  XNOR2_X1 U413 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n368) );
  XNOR2_X1 U415 ( .A(G36GAT), .B(G190GAT), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n355), .B(G218GAT), .ZN(n399) );
  NAND2_X1 U417 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n291), .B(n357), .ZN(n359) );
  INV_X1 U419 ( .A(G92GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n360), .B(G134GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U423 ( .A(G50GAT), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U424 ( .A(G106GAT), .B(n413), .ZN(n364) );
  INV_X1 U425 ( .A(KEYINPUT9), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n386) );
  XOR2_X1 U427 ( .A(G22GAT), .B(G155GAT), .Z(n412) );
  XOR2_X1 U428 ( .A(n412), .B(KEYINPUT15), .Z(n370) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U431 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n372) );
  XNOR2_X1 U432 ( .A(G64GAT), .B(KEYINPUT74), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U434 ( .A(n374), .B(n373), .Z(n379) );
  XNOR2_X1 U435 ( .A(G127GAT), .B(G211GAT), .ZN(n375) );
  XOR2_X1 U436 ( .A(G8GAT), .B(G183GAT), .Z(n396) );
  XNOR2_X1 U437 ( .A(n375), .B(n396), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U440 ( .A(n381), .B(n380), .Z(n576) );
  INV_X1 U441 ( .A(n576), .ZN(n480) );
  XNOR2_X1 U442 ( .A(KEYINPUT106), .B(n480), .ZN(n559) );
  NOR2_X1 U443 ( .A1(n386), .A2(n559), .ZN(n382) );
  NAND2_X1 U444 ( .A1(n383), .A2(n382), .ZN(n385) );
  XNOR2_X1 U445 ( .A(KEYINPUT36), .B(n386), .ZN(n580) );
  AND2_X1 U446 ( .A1(n580), .A2(n480), .ZN(n389) );
  INV_X1 U447 ( .A(KEYINPUT108), .ZN(n387) );
  NOR2_X1 U448 ( .A1(n571), .A2(n390), .ZN(n391) );
  NAND2_X1 U449 ( .A1(n391), .A2(n566), .ZN(n392) );
  NAND2_X1 U450 ( .A1(n393), .A2(n392), .ZN(n395) );
  XOR2_X1 U451 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n394) );
  XOR2_X1 U452 ( .A(KEYINPUT89), .B(n396), .Z(n398) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n408) );
  XOR2_X1 U455 ( .A(n400), .B(n399), .Z(n406) );
  XOR2_X1 U456 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n402) );
  XNOR2_X1 U457 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n437) );
  XOR2_X1 U459 ( .A(G211GAT), .B(KEYINPUT21), .Z(n404) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(KEYINPUT81), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n422) );
  XNOR2_X1 U462 ( .A(n437), .B(n422), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n511) );
  XOR2_X1 U465 ( .A(n511), .B(KEYINPUT116), .Z(n409) );
  NOR2_X1 U466 ( .A1(n538), .A2(n409), .ZN(n410) );
  XOR2_X1 U467 ( .A(KEYINPUT54), .B(n410), .Z(n411) );
  XOR2_X1 U468 ( .A(G78GAT), .B(G218GAT), .Z(n415) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n427) );
  XOR2_X1 U471 ( .A(G204GAT), .B(KEYINPUT79), .Z(n417) );
  XNOR2_X1 U472 ( .A(KEYINPUT85), .B(KEYINPUT22), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U474 ( .A(KEYINPUT24), .B(KEYINPUT80), .Z(n419) );
  XNOR2_X1 U475 ( .A(KEYINPUT84), .B(KEYINPUT23), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U477 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U480 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n431), .B(n430), .ZN(n460) );
  NAND2_X1 U484 ( .A1(n564), .A2(n460), .ZN(n434) );
  XOR2_X1 U485 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n432) );
  XOR2_X1 U486 ( .A(G190GAT), .B(G43GAT), .Z(n436) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U489 ( .A(n438), .B(n437), .Z(n446) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT77), .Z(n440) );
  XNOR2_X1 U491 ( .A(G99GAT), .B(KEYINPUT78), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U493 ( .A(G183GAT), .B(G71GAT), .Z(n442) );
  XNOR2_X1 U494 ( .A(G15GAT), .B(G176GAT), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U498 ( .A1(n449), .A2(n522), .ZN(n553) );
  INV_X1 U499 ( .A(n553), .ZN(n560) );
  NAND2_X1 U500 ( .A1(n560), .A2(n386), .ZN(n451) );
  XOR2_X1 U501 ( .A(KEYINPUT34), .B(KEYINPUT94), .Z(n470) );
  NOR2_X1 U502 ( .A1(n566), .A2(n571), .ZN(n483) );
  AND2_X1 U503 ( .A1(n522), .A2(n511), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n452), .B(KEYINPUT91), .ZN(n453) );
  NAND2_X1 U505 ( .A1(n453), .A2(n460), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT25), .B(n454), .Z(n457) );
  XNOR2_X1 U507 ( .A(n511), .B(KEYINPUT27), .ZN(n461) );
  NOR2_X1 U508 ( .A1(n460), .A2(n522), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n455), .B(KEYINPUT26), .ZN(n563) );
  NAND2_X1 U510 ( .A1(n461), .A2(n563), .ZN(n456) );
  NAND2_X1 U511 ( .A1(n457), .A2(n456), .ZN(n458) );
  XOR2_X1 U512 ( .A(KEYINPUT92), .B(n458), .Z(n459) );
  NOR2_X1 U513 ( .A1(n507), .A2(n459), .ZN(n464) );
  XOR2_X1 U514 ( .A(KEYINPUT28), .B(n460), .Z(n515) );
  NAND2_X1 U515 ( .A1(n461), .A2(n507), .ZN(n462) );
  XNOR2_X1 U516 ( .A(KEYINPUT90), .B(n462), .ZN(n537) );
  OR2_X1 U517 ( .A1(n515), .A2(n537), .ZN(n521) );
  NOR2_X1 U518 ( .A1(n521), .A2(n522), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n479) );
  NOR2_X1 U520 ( .A1(n386), .A2(n576), .ZN(n466) );
  XNOR2_X1 U521 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n467) );
  NOR2_X1 U523 ( .A1(n479), .A2(n467), .ZN(n468) );
  XOR2_X1 U524 ( .A(KEYINPUT93), .B(n468), .Z(n495) );
  AND2_X1 U525 ( .A1(n483), .A2(n495), .ZN(n476) );
  NAND2_X1 U526 ( .A1(n476), .A2(n507), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U528 ( .A(G1GAT), .B(n471), .Z(G1324GAT) );
  NAND2_X1 U529 ( .A1(n511), .A2(n476), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT35), .B(KEYINPUT95), .Z(n474) );
  NAND2_X1 U532 ( .A1(n476), .A2(n522), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U534 ( .A(G15GAT), .B(n475), .Z(G1326GAT) );
  NAND2_X1 U535 ( .A1(n515), .A2(n476), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT96), .ZN(n478) );
  XNOR2_X1 U537 ( .A(G22GAT), .B(n478), .ZN(G1327GAT) );
  XOR2_X1 U538 ( .A(G29GAT), .B(KEYINPUT39), .Z(n487) );
  NOR2_X1 U539 ( .A1(n480), .A2(n479), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n580), .A2(n481), .ZN(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT37), .B(n482), .ZN(n506) );
  NAND2_X1 U542 ( .A1(n483), .A2(n506), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(KEYINPUT97), .ZN(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT38), .B(n485), .ZN(n491) );
  NAND2_X1 U545 ( .A1(n507), .A2(n491), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  NAND2_X1 U547 ( .A1(n491), .A2(n511), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U549 ( .A1(n491), .A2(n522), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  XNOR2_X1 U552 ( .A(G50GAT), .B(KEYINPUT98), .ZN(n493) );
  NAND2_X1 U553 ( .A1(n515), .A2(n491), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1331GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT99), .B(KEYINPUT42), .Z(n497) );
  INV_X1 U556 ( .A(n566), .ZN(n494) );
  NOR2_X1 U557 ( .A1(n552), .A2(n494), .ZN(n505) );
  AND2_X1 U558 ( .A1(n495), .A2(n505), .ZN(n502) );
  NAND2_X1 U559 ( .A1(n502), .A2(n507), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n498), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n511), .A2(n502), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT100), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(n500), .ZN(G1333GAT) );
  NAND2_X1 U565 ( .A1(n522), .A2(n502), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U567 ( .A(G78GAT), .B(KEYINPUT43), .Z(n504) );
  NAND2_X1 U568 ( .A1(n502), .A2(n515), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n509) );
  AND2_X1 U571 ( .A1(n506), .A2(n505), .ZN(n516) );
  NAND2_X1 U572 ( .A1(n516), .A2(n507), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  XOR2_X1 U575 ( .A(G92GAT), .B(KEYINPUT103), .Z(n513) );
  NAND2_X1 U576 ( .A1(n516), .A2(n511), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n522), .A2(n516), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U580 ( .A(G106GAT), .B(KEYINPUT104), .ZN(n520) );
  XOR2_X1 U581 ( .A(KEYINPUT105), .B(KEYINPUT44), .Z(n518) );
  NAND2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1339GAT) );
  NOR2_X1 U585 ( .A1(n538), .A2(n521), .ZN(n523) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n566), .A2(n529), .ZN(n525) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(KEYINPUT109), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(G1340GAT) );
  NOR2_X1 U590 ( .A1(n552), .A2(n529), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT49), .B(KEYINPUT110), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(n528), .ZN(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT111), .B(KEYINPUT50), .Z(n531) );
  INV_X1 U595 ( .A(n529), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n533), .A2(n559), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n535) );
  NAND2_X1 U600 ( .A1(n533), .A2(n386), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G134GAT), .B(n536), .ZN(G1343GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n539), .A2(n563), .ZN(n547) );
  NOR2_X1 U605 ( .A1(n566), .A2(n547), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT113), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n543) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n552), .A2(n547), .ZN(n544) );
  XOR2_X1 U612 ( .A(n545), .B(n544), .Z(G1345GAT) );
  NOR2_X1 U613 ( .A1(n576), .A2(n547), .ZN(n546) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n546), .Z(G1346GAT) );
  INV_X1 U615 ( .A(n386), .ZN(n548) );
  NOR2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G162GAT), .B(KEYINPUT115), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1347GAT) );
  NOR2_X1 U619 ( .A1(n566), .A2(n553), .ZN(n551) );
  XOR2_X1 U620 ( .A(G169GAT), .B(n551), .Z(G1348GAT) );
  NOR2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n555) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U625 ( .A(KEYINPUT56), .B(n556), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U631 ( .A1(n577), .A2(n566), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  INV_X1 U636 ( .A(n577), .ZN(n579) );
  AND2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n573) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(G218GAT), .B(n583), .Z(G1355GAT) );
endmodule

