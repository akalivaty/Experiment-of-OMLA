//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT65), .B(G68), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n207), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n203), .A2(G50), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT0), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n207), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n223), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n227), .B1(new_n224), .B2(new_n226), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n218), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT67), .B(G107), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G200), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G97), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G226), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n252), .B(new_n253), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT72), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT72), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n263), .B2(new_n219), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT68), .A2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT68), .A2(G41), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT69), .B(G45), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n267), .B(G274), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT70), .A2(G1), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT70), .A2(G1), .ZN(new_n275));
  OAI22_X1  g0075(.A1(new_n274), .A2(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT71), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT71), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n278), .B1(G41), .B2(G45), .C1(new_n274), .C2(new_n275), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n220), .B1(new_n261), .B2(new_n262), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n277), .A2(new_n279), .A3(G238), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n266), .A2(new_n273), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n283), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n266), .A2(new_n273), .A3(new_n285), .A4(new_n281), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n250), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n219), .ZN(new_n289));
  INV_X1    g0089(.A(G20), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n208), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G77), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n293), .A2(new_n243), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n289), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT11), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT70), .A2(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT70), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G13), .A3(G20), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G68), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT12), .ZN(new_n304));
  INV_X1    g0104(.A(new_n302), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT12), .A3(new_n209), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n290), .B1(new_n299), .B2(new_n300), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n289), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G68), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n298), .A2(new_n304), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n287), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n282), .A2(KEYINPUT13), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(G190), .A3(new_n286), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n284), .B2(new_n286), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n312), .A2(G179), .A3(new_n286), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n316), .B2(new_n317), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n310), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n251), .A2(G222), .A3(new_n254), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n251), .A2(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G223), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(new_n295), .B2(new_n251), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n265), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n277), .A2(new_n280), .A3(new_n279), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G226), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n328), .A3(new_n273), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  OR3_X1    g0130(.A1(new_n329), .A2(new_n330), .A3(G179), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n329), .B2(G179), .ZN(new_n332));
  OAI21_X1  g0132(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n333));
  INV_X1    g0133(.A(G150), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n333), .B1(new_n334), .B2(new_n293), .C1(new_n335), .C2(new_n294), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n289), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n301), .A2(G20), .ZN(new_n338));
  INV_X1    g0138(.A(new_n289), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(G50), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n307), .A2(G13), .A3(new_n243), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n329), .A2(new_n315), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n331), .A2(new_n332), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n337), .A3(KEYINPUT76), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT76), .ZN(new_n348));
  XOR2_X1   g0148(.A(KEYINPUT8), .B(G58), .Z(new_n349));
  INV_X1    g0149(.A(new_n294), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n349), .A2(new_n350), .B1(G150), .B2(new_n292), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n339), .B1(new_n351), .B2(new_n333), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n348), .B1(new_n352), .B2(new_n342), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n329), .A2(G200), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT9), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n347), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n326), .A2(new_n328), .A3(G190), .A4(new_n273), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n355), .A2(new_n356), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT10), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n358), .A2(new_n359), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT10), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(new_n356), .A4(new_n355), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n346), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n273), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n251), .A2(G232), .A3(new_n254), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n367), .B1(new_n368), .B2(new_n251), .C1(new_n323), .C2(new_n210), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n366), .B1(new_n369), .B2(new_n265), .ZN(new_n370));
  INV_X1    g0170(.A(G179), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n327), .A2(G244), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(G169), .B1(new_n370), .B2(new_n372), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n335), .B1(KEYINPUT74), .B2(new_n293), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(KEYINPUT74), .B2(new_n293), .ZN(new_n377));
  XOR2_X1   g0177(.A(KEYINPUT15), .B(G87), .Z(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(new_n350), .B1(G20), .B2(G77), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n339), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n308), .A2(G77), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G77), .B2(new_n302), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n374), .A2(new_n375), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n369), .A2(new_n265), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n386), .A2(new_n372), .A3(G190), .A4(new_n273), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n383), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n250), .B1(new_n370), .B2(new_n372), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(KEYINPUT75), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n388), .A2(new_n389), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n365), .A2(new_n395), .A3(KEYINPUT77), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT77), .B1(new_n365), .B2(new_n395), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n314), .B(new_n321), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n277), .A2(new_n279), .A3(G232), .A4(new_n280), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n273), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT82), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(KEYINPUT82), .A3(new_n273), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n251), .A2(G223), .A3(new_n254), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT81), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n407), .C1(new_n323), .C2(new_n256), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n265), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n403), .A2(new_n371), .A3(new_n404), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT83), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n401), .A2(new_n402), .B1(new_n265), .B2(new_n408), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT83), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n371), .A4(new_n404), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n403), .A2(new_n404), .A3(new_n409), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n315), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n302), .A2(new_n335), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n308), .B2(new_n335), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G159), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n293), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT65), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G68), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n425), .A3(G58), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n203), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G20), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT80), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n422), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(KEYINPUT80), .A3(G20), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT7), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n251), .A2(new_n432), .A3(G20), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT3), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G33), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT7), .B1(new_n437), .B2(new_n290), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n208), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n430), .A2(new_n431), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT16), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n339), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n432), .B1(new_n251), .B2(G20), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n435), .A2(G33), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT7), .B(new_n290), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(KEYINPUT79), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(new_n432), .C1(new_n251), .C2(G20), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(G68), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n450), .A2(new_n430), .A3(KEYINPUT16), .A4(new_n431), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n420), .B1(new_n442), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n399), .B1(new_n417), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(KEYINPUT83), .A2(new_n410), .B1(new_n415), .B2(new_n315), .ZN(new_n454));
  INV_X1    g0254(.A(new_n203), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n208), .B2(G58), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n429), .B1(new_n456), .B2(new_n290), .ZN(new_n457));
  INV_X1    g0257(.A(new_n422), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n431), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n439), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n441), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(new_n289), .A3(new_n451), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n419), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n454), .A2(new_n463), .A3(KEYINPUT18), .A4(new_n414), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n453), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n415), .A2(G200), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n412), .A2(G190), .A3(new_n404), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(new_n462), .A3(new_n419), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT17), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT17), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n452), .A2(new_n470), .A3(new_n466), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT84), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n398), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n251), .A2(G257), .A3(new_n254), .ZN(new_n476));
  INV_X1    g0276(.A(G303), .ZN(new_n477));
  INV_X1    g0277(.A(G264), .ZN(new_n478));
  OAI221_X1 g0278(.A(new_n476), .B1(new_n477), .B2(new_n251), .C1(new_n323), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n265), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT87), .B1(new_n482), .B2(G41), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT87), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n262), .A3(KEYINPUT5), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n280), .A3(G274), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT68), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n262), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(new_n482), .A3(new_n268), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(G45), .B1(new_n274), .B2(new_n275), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT86), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G45), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n299), .B2(new_n300), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT86), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n490), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n487), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n490), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(G270), .A3(new_n280), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT91), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n487), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n495), .A2(new_n496), .A3(new_n490), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n496), .B1(new_n495), .B2(new_n490), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT91), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n508), .A3(new_n501), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n481), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n301), .A2(G33), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n302), .A2(new_n511), .A3(G116), .A4(new_n339), .ZN(new_n512));
  INV_X1    g0312(.A(G116), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n307), .A2(G13), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(G20), .B1(G33), .B2(G283), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n261), .A2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT92), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n288), .A2(new_n219), .B1(G20), .B2(new_n513), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT20), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n518), .A2(KEYINPUT92), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT92), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n516), .B2(new_n517), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n520), .B(KEYINPUT20), .C1(new_n522), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n515), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G169), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n510), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT93), .B1(new_n529), .B2(KEYINPUT21), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT21), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n510), .B2(new_n528), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n510), .A2(G179), .A3(new_n527), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT93), .ZN(new_n535));
  NOR4_X1   g0335(.A1(new_n510), .A2(new_n528), .A3(new_n535), .A4(new_n531), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n530), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n509), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n508), .B1(new_n507), .B2(new_n501), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n480), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n527), .B1(new_n540), .B2(G200), .ZN(new_n541));
  INV_X1    g0341(.A(G190), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n540), .ZN(new_n543));
  XNOR2_X1  g0343(.A(KEYINPUT89), .B(G87), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT90), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT90), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n548), .A3(new_n545), .ZN(new_n549));
  NAND3_X1  g0349(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n547), .A2(new_n549), .B1(new_n290), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n251), .A2(new_n290), .A3(G68), .ZN(new_n552));
  INV_X1    g0352(.A(G97), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n294), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(KEYINPUT19), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n289), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n302), .A2(new_n339), .A3(new_n511), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G87), .ZN(new_n559));
  INV_X1    g0359(.A(new_n378), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n305), .A2(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n556), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G274), .ZN(new_n563));
  OAI211_X1 g0363(.A(G45), .B(new_n563), .C1(new_n274), .C2(new_n275), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n280), .B(new_n564), .C1(new_n495), .C2(G250), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT88), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G250), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n258), .B1(new_n492), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(KEYINPUT88), .A3(new_n564), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n251), .A2(G244), .A3(G1698), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n255), .C2(new_n210), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n265), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n567), .A2(new_n570), .B1(new_n574), .B2(new_n265), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n562), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n434), .A2(new_n436), .A3(G244), .A4(new_n254), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT4), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n254), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G283), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n265), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n500), .A2(G257), .A3(new_n280), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n507), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G200), .ZN(new_n591));
  OAI21_X1  g0391(.A(G107), .B1(new_n433), .B2(new_n438), .ZN(new_n592));
  XNOR2_X1  g0392(.A(G97), .B(G107), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT6), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT85), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n553), .A2(KEYINPUT6), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(new_n595), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n596), .A2(G20), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n292), .A2(G77), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n592), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n289), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n302), .A2(G97), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n558), .B2(G97), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n588), .A2(new_n507), .A3(G190), .A4(new_n589), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n591), .A2(new_n602), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n604), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n588), .A2(new_n507), .A3(new_n371), .A4(new_n589), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n590), .A2(new_n315), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n558), .A2(new_n378), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n556), .A2(new_n561), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n576), .A2(new_n315), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n578), .A2(new_n371), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n580), .A2(new_n606), .A3(new_n610), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n500), .A2(G264), .A3(new_n280), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n434), .A2(new_n436), .A3(G250), .A4(new_n254), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n434), .A2(new_n436), .A3(G257), .A4(G1698), .ZN(new_n619));
  INV_X1    g0419(.A(G294), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n619), .C1(new_n261), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n265), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n507), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n315), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n507), .A2(new_n371), .A3(new_n617), .A4(new_n622), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT25), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n302), .B2(G107), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n307), .A2(KEYINPUT25), .A3(G13), .A4(new_n368), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n368), .B2(new_n557), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n434), .A2(new_n436), .A3(new_n290), .A4(G87), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT22), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT22), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n251), .A2(new_n634), .A3(new_n290), .A4(G87), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n573), .A2(G20), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT94), .B1(new_n290), .B2(G107), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT23), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT23), .ZN(new_n640));
  OAI211_X1 g0440(.A(KEYINPUT94), .B(new_n640), .C1(new_n290), .C2(G107), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n637), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n636), .A2(KEYINPUT24), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n642), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT24), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n339), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n631), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n626), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n645), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n289), .A3(new_n643), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n622), .A2(new_n617), .ZN(new_n651));
  OAI21_X1  g0451(.A(G200), .B1(new_n651), .B2(new_n498), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n558), .A2(G107), .B1(new_n628), .B2(new_n629), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n507), .A2(G190), .A3(new_n617), .A4(new_n622), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n650), .A2(new_n652), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT95), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n647), .A2(new_n654), .A3(new_n652), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n650), .A2(new_n653), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n624), .A3(new_n625), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT95), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n616), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n475), .A2(new_n537), .A3(new_n543), .A4(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n615), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n532), .A2(new_n533), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n527), .A2(G169), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n540), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n535), .B1(new_n667), .B2(new_n531), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n529), .A2(KEYINPUT93), .A3(KEYINPUT21), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n665), .A2(new_n668), .A3(new_n669), .A4(new_n659), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n606), .A2(new_n610), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n577), .A2(KEYINPUT96), .ZN(new_n672));
  OR3_X1    g0472(.A1(new_n578), .A2(KEYINPUT96), .A3(new_n250), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n579), .A4(new_n562), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n671), .A2(new_n657), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n664), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n580), .A2(new_n615), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT26), .B1(new_n677), .B2(new_n610), .ZN(new_n678));
  INV_X1    g0478(.A(new_n610), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n674), .A2(new_n679), .A3(new_n680), .A4(new_n615), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n475), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n321), .A2(new_n385), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(new_n472), .A3(new_n314), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n465), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n361), .A2(new_n364), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n346), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n684), .A2(new_n690), .ZN(G369));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n290), .A2(G13), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n301), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n527), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n537), .A2(new_n543), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n665), .A2(new_n669), .A3(new_n668), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n527), .A3(new_n699), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n692), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n699), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n659), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT98), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n656), .A2(new_n661), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n658), .A2(new_n699), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n537), .A2(new_n699), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n712), .A2(new_n716), .B1(new_n648), .B2(new_n706), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(G399));
  NAND3_X1  g0518(.A1(new_n547), .A2(new_n513), .A3(new_n549), .ZN(new_n719));
  INV_X1    g0519(.A(new_n225), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n271), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n719), .A2(new_n267), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n222), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(KEYINPUT99), .B(KEYINPUT28), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n699), .B1(new_n676), .B2(new_n682), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n537), .A2(new_n662), .A3(new_n543), .A4(new_n706), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  INV_X1    g0531(.A(new_n623), .ZN(new_n732));
  AND4_X1   g0532(.A1(new_n732), .A2(new_n589), .A3(new_n588), .A4(new_n578), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(G179), .A3(new_n510), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n733), .A2(KEYINPUT30), .A3(G179), .A4(new_n510), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n732), .A2(G179), .A3(new_n578), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n540), .A3(new_n590), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n731), .B1(new_n740), .B2(new_n699), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n730), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n731), .A3(new_n699), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(G330), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n677), .A2(KEYINPUT26), .A3(new_n610), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n674), .A2(new_n615), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n679), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(new_n748), .B2(KEYINPUT26), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n699), .B1(new_n676), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n728), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n729), .A2(new_n745), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n726), .B1(new_n752), .B2(G1), .ZN(G364));
  AOI21_X1  g0553(.A(new_n267), .B1(new_n693), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n721), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n219), .B1(G20), .B2(new_n315), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n290), .A2(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n421), .ZN(new_n763));
  XNOR2_X1  g0563(.A(KEYINPUT102), .B(KEYINPUT32), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n765), .B1(new_n553), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(G20), .A2(G179), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT101), .Z(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n542), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n250), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n250), .A2(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n760), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n775), .A2(G20), .A3(G190), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n251), .B1(new_n776), .B2(new_n368), .C1(new_n544), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n774), .A2(new_n202), .B1(KEYINPUT103), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n771), .A2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n250), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n769), .B(new_n780), .C1(G50), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(G200), .ZN(new_n784));
  AOI22_X1  g0584(.A1(KEYINPUT103), .A2(new_n779), .B1(new_n784), .B2(G58), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n772), .A2(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n783), .B(new_n785), .C1(new_n295), .C2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n777), .ZN(new_n789));
  INV_X1    g0589(.A(new_n762), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n789), .A2(G303), .B1(new_n790), .B2(G329), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n437), .C1(new_n792), .C2(new_n776), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G294), .B2(new_n767), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n782), .A2(G326), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n773), .A2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G311), .A2(new_n786), .B1(new_n784), .B2(G322), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n794), .A2(new_n795), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n759), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n759), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT100), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n720), .A2(new_n437), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G355), .A2(new_n807), .B1(new_n513), .B2(new_n720), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n248), .A2(new_n494), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n720), .A2(new_n251), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n222), .B2(new_n272), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n808), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n757), .B(new_n800), .C1(new_n806), .C2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT104), .Z(new_n814));
  NAND3_X1  g0614(.A1(new_n701), .A2(new_n703), .A3(new_n803), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n701), .A2(new_n703), .A3(new_n692), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n705), .A2(new_n757), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  OAI21_X1  g0620(.A(new_n390), .B1(new_n383), .B2(new_n706), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n385), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n384), .A2(new_n706), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n727), .B(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n756), .B1(new_n826), .B2(new_n744), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n744), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n758), .A2(new_n801), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n757), .B1(new_n295), .B2(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G150), .A2(new_n773), .B1(new_n786), .B2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  INV_X1    g0632(.A(new_n782), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  INV_X1    g0634(.A(new_n784), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n831), .B1(new_n832), .B2(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n251), .B1(new_n762), .B2(new_n839), .C1(new_n768), .C2(new_n201), .ZN(new_n840));
  INV_X1    g0640(.A(new_n776), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G68), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n243), .B2(new_n777), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n840), .B1(KEYINPUT106), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(KEYINPUT106), .B2(new_n843), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n836), .B2(new_n837), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G283), .A2(new_n773), .B1(new_n782), .B2(G303), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n513), .B2(new_n787), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT105), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n768), .A2(new_n553), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n789), .A2(G107), .B1(new_n841), .B2(G87), .ZN(new_n851));
  INV_X1    g0651(.A(G311), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n851), .B(new_n437), .C1(new_n852), .C2(new_n762), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n850), .B(new_n853), .C1(G294), .C2(new_n784), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n838), .A2(new_n846), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n830), .B1(new_n855), .B2(new_n759), .C1(new_n825), .C2(new_n802), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n828), .A2(new_n856), .ZN(G384));
  NAND3_X1  g0657(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT35), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n513), .B(new_n221), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n860), .A2(KEYINPUT107), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(KEYINPUT107), .B2(new_n860), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT36), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n723), .A2(G77), .A3(new_n426), .ZN(new_n864));
  AOI211_X1 g0664(.A(G13), .B(new_n301), .C1(new_n864), .C2(new_n244), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n451), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n450), .A2(new_n430), .A3(new_n431), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n339), .B1(new_n868), .B2(new_n441), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n867), .B1(new_n869), .B2(KEYINPUT108), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT108), .ZN(new_n871));
  INV_X1    g0671(.A(new_n459), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n872), .B2(new_n450), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n873), .B2(new_n339), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n420), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n468), .B1(new_n875), .B2(new_n697), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n417), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n697), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n463), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(new_n468), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n454), .A2(new_n463), .A3(new_n414), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n875), .A2(new_n697), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT109), .B1(new_n473), .B2(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n453), .A2(new_n464), .B1(new_n469), .B2(new_n471), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT109), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n870), .A2(new_n874), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n879), .B1(new_n890), .B2(new_n420), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(KEYINPUT38), .B(new_n885), .C1(new_n887), .C2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n882), .B1(new_n881), .B2(new_n883), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n888), .A2(new_n880), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n310), .A2(new_n699), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n321), .A2(new_n314), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n310), .B(new_n699), .C1(new_n318), .C2(new_n320), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n824), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n742), .A2(new_n743), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n742), .A2(new_n743), .A3(new_n904), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n885), .B1(new_n887), .B2(new_n892), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n894), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n909), .B2(new_n893), .ZN(new_n910));
  OAI211_X1 g0710(.A(G330), .B(new_n906), .C1(new_n910), .C2(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n475), .A2(new_n745), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n742), .A2(KEYINPUT40), .A3(new_n904), .A4(new_n743), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n893), .B2(new_n899), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n473), .A2(KEYINPUT109), .A3(new_n886), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n889), .B1(new_n888), .B2(new_n891), .ZN(new_n917));
  AOI221_X4 g0717(.A(new_n894), .B1(new_n878), .B2(new_n884), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n919), .B2(new_n885), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n905), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n475), .A2(new_n742), .A3(new_n743), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n913), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n475), .B1(new_n729), .B2(new_n751), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n690), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n321), .A2(new_n699), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n909), .B2(new_n893), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n893), .A2(new_n899), .A3(new_n931), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n930), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n465), .A2(new_n879), .ZN(new_n936));
  INV_X1    g0736(.A(new_n823), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n727), .B2(new_n825), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n902), .A2(new_n903), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n909), .A2(new_n893), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n935), .A2(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n929), .A2(new_n943), .B1(new_n301), .B2(new_n693), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n929), .A2(new_n943), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n866), .B1(new_n944), .B2(new_n945), .ZN(G367));
  NAND2_X1  g0746(.A1(new_n607), .A2(new_n699), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n671), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n679), .A2(new_n699), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n712), .A2(new_n716), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n610), .B1(new_n948), .B2(new_n659), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n706), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n562), .A2(new_n706), .ZN(new_n957));
  MUX2_X1   g0757(.A(new_n747), .B(new_n664), .S(new_n957), .Z(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT110), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n956), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n950), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n715), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n960), .B1(new_n956), .B2(new_n962), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n966), .B1(new_n963), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n721), .B(KEYINPUT41), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n704), .A2(new_n716), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n712), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n752), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n712), .A2(new_n716), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n648), .A2(new_n706), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(KEYINPUT44), .A3(new_n964), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n717), .B2(new_n950), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n982));
  NAND3_X1  g0782(.A1(new_n717), .A2(new_n950), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n982), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n977), .B2(new_n964), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n981), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT112), .B1(new_n986), .B2(new_n714), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n985), .A2(new_n983), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT112), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n988), .A2(new_n715), .A3(new_n981), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n974), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n752), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n971), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n970), .B1(new_n993), .B2(new_n754), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n958), .A2(new_n804), .ZN(new_n995));
  INV_X1    g0795(.A(new_n810), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n237), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n806), .B1(new_n225), .B2(new_n560), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n756), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT113), .B(G311), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G294), .A2(new_n773), .B1(new_n782), .B2(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n792), .B2(new_n787), .C1(new_n477), .C2(new_n835), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n789), .A2(G116), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT46), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1003), .A2(new_n1004), .B1(G107), .B2(new_n767), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n437), .B1(new_n762), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G97), .B2(new_n841), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1005), .B(new_n1008), .C1(new_n1004), .C2(new_n1003), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n777), .A2(new_n201), .B1(new_n776), .B2(new_n295), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT114), .B(G137), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n437), .B(new_n1010), .C1(new_n790), .C2(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n202), .B2(new_n768), .C1(new_n835), .C2(new_n334), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G143), .A2(new_n782), .B1(new_n773), .B2(G159), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n243), .B2(new_n787), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1002), .A2(new_n1009), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT47), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n759), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n999), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n995), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n994), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(G387));
  NAND2_X1  g0824(.A1(new_n973), .A2(new_n755), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n996), .B1(new_n233), .B2(new_n272), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n719), .B2(new_n807), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n349), .A2(new_n243), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n494), .B1(new_n202), .B2(new_n295), .C1(new_n1028), .C2(KEYINPUT50), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n719), .B(new_n1029), .C1(KEYINPUT50), .C2(new_n1028), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1027), .A2(new_n1030), .B1(G107), .B2(new_n225), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n757), .B1(new_n1031), .B2(new_n806), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n782), .A2(G159), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT115), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n786), .A2(G68), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n767), .A2(new_n378), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n437), .B1(new_n841), .B2(G97), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n789), .A2(G77), .B1(new_n790), .B2(G150), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n243), .A2(new_n835), .B1(new_n774), .B2(new_n335), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1034), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G322), .A2(new_n782), .B1(new_n773), .B2(new_n1000), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n477), .B2(new_n787), .C1(new_n1006), .C2(new_n835), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT48), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n792), .B2(new_n768), .C1(new_n620), .C2(new_n777), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n251), .B1(new_n790), .B2(G326), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n513), .B2(new_n776), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1041), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1032), .B1(new_n712), .B2(new_n804), .C1(new_n1051), .C2(new_n759), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n974), .A2(new_n721), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n973), .A2(new_n752), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1025), .B(new_n1052), .C1(new_n1053), .C2(new_n1054), .ZN(G393));
  NAND2_X1  g0855(.A1(new_n987), .A2(new_n990), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n986), .A2(new_n714), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n974), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n721), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n991), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n987), .A2(new_n990), .B1(new_n714), .B2(new_n986), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n964), .A2(new_n803), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n242), .A2(new_n996), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n806), .B1(new_n553), .B2(new_n225), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n756), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n768), .A2(new_n295), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n437), .B1(new_n841), .B2(G87), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n834), .B2(new_n762), .C1(new_n209), .C2(new_n777), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(new_n349), .C2(new_n786), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G150), .A2(new_n782), .B1(new_n784), .B2(G159), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT51), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(new_n243), .C2(new_n774), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1072), .A2(KEYINPUT51), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n852), .A2(new_n835), .B1(new_n833), .B2(new_n1006), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT52), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n789), .A2(G283), .B1(new_n790), .B2(G322), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(KEYINPUT116), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(KEYINPUT116), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n437), .B1(new_n776), .B2(new_n368), .C1(new_n768), .C2(new_n513), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G294), .A2(new_n786), .B1(new_n773), .B2(G303), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1078), .A2(new_n1081), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1074), .A2(new_n1075), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1067), .B1(new_n1088), .B2(new_n758), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1063), .A2(new_n755), .B1(new_n1064), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1062), .A2(new_n1090), .ZN(G390));
  AND3_X1   g0891(.A1(new_n927), .A2(new_n690), .A3(new_n912), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n905), .A2(G330), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n937), .B1(new_n750), .B2(new_n822), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n742), .A2(G330), .A3(new_n743), .A4(new_n825), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n939), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n905), .A2(G330), .B1(new_n1095), .B2(new_n939), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n938), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT39), .B1(new_n918), .B2(new_n920), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n930), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n938), .B2(new_n939), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1103), .A3(new_n933), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n900), .B(new_n1102), .C1(new_n939), .C2(new_n1094), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1104), .A2(new_n1093), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1093), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1100), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1093), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n927), .A2(new_n690), .A3(new_n912), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1098), .A2(new_n938), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n1097), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1104), .A2(new_n1093), .A3(new_n1105), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1108), .A2(new_n1116), .A3(new_n721), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n829), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G97), .A2(new_n786), .B1(new_n782), .B2(G283), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n368), .B2(new_n774), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n835), .A2(new_n513), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n789), .A2(G87), .B1(new_n790), .B2(G294), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n437), .A3(new_n842), .ZN(new_n1123));
  NOR4_X1   g0923(.A1(new_n1120), .A2(new_n1068), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n251), .B1(new_n776), .B2(new_n243), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT117), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n777), .A2(new_n334), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n790), .A2(G125), .B1(new_n767), .B2(G159), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n787), .A2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(new_n773), .C2(new_n1011), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G128), .A2(new_n782), .B1(new_n784), .B2(G132), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT118), .Z(new_n1135));
  AOI21_X1  g0935(.A(new_n1124), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n756), .B1(new_n349), .B2(new_n1118), .C1(new_n1136), .C2(new_n759), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n932), .A2(new_n934), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n801), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n755), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1117), .A2(new_n1141), .ZN(G378));
  INV_X1    g0942(.A(KEYINPUT122), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n935), .B2(new_n942), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n689), .A2(new_n345), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n347), .A2(new_n353), .A3(new_n879), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT121), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n911), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT121), .B1(new_n923), .B2(G330), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1150), .B1(new_n1151), .B2(new_n911), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1145), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1148), .B(new_n1149), .Z(new_n1158));
  NAND2_X1  g0958(.A1(new_n911), .A2(new_n1151), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n921), .A2(new_n922), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1160), .A2(KEYINPUT121), .A3(G330), .A4(new_n906), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1158), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1162), .A2(new_n1144), .A3(new_n1155), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n755), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n756), .B1(G50), .B2(new_n1118), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n271), .A2(new_n251), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G50), .B(new_n1166), .C1(new_n261), .C2(new_n262), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n833), .A2(new_n513), .B1(new_n202), .B2(new_n768), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT119), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT119), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n251), .B(new_n271), .C1(new_n789), .C2(G77), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n201), .B2(new_n776), .C1(new_n792), .C2(new_n762), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G97), .B2(new_n773), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G107), .A2(new_n784), .B1(new_n786), .B2(new_n378), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1169), .A2(new_n1170), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1167), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n768), .A2(new_n334), .B1(new_n1131), .B2(new_n777), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G128), .A2(new_n784), .B1(new_n773), .B2(G132), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n832), .B2(new_n787), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G125), .C2(new_n782), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(G33), .B(G41), .C1(new_n790), .C2(G124), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n421), .B2(new_n776), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT120), .Z(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1177), .B1(new_n1176), .B2(new_n1175), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1165), .B1(new_n1189), .B2(new_n758), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1158), .B2(new_n802), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1154), .A2(new_n1145), .A3(new_n1156), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1144), .B1(new_n1162), .B2(new_n1155), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1192), .A2(new_n1193), .B1(new_n1092), .B2(new_n1116), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT57), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT57), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1116), .B2(new_n1092), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1154), .A2(new_n943), .A3(new_n1156), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n943), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1162), .B2(new_n1155), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n721), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1164), .B(new_n1191), .C1(new_n1195), .C2(new_n1202), .ZN(G375));
  AOI22_X1  g1003(.A1(G107), .A2(new_n786), .B1(new_n784), .B2(G283), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n513), .B2(new_n774), .C1(new_n620), .C2(new_n833), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n437), .B1(new_n776), .B2(new_n295), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT123), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT123), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n789), .A2(G97), .B1(new_n790), .B2(G303), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1207), .A2(new_n1036), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n777), .A2(new_n421), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n251), .B1(new_n776), .B2(new_n201), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G128), .C2(new_n790), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n243), .B2(new_n768), .C1(new_n787), .C2(new_n334), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n784), .A2(new_n1011), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n833), .B2(new_n839), .C1(new_n774), .C2(new_n1131), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1205), .A2(new_n1210), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n758), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1218), .B(new_n756), .C1(G68), .C2(new_n1118), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n939), .B2(new_n801), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1099), .B2(new_n755), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1100), .A2(new_n971), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(G381));
  NAND2_X1  g1024(.A1(new_n1164), .A2(new_n1191), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n943), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1162), .A2(new_n1199), .A3(new_n1155), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1060), .B1(new_n1228), .B2(new_n1197), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1116), .A2(new_n1092), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1196), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1225), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(G378), .ZN(new_n1234));
  OR2_X1    g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(G390), .A2(new_n1235), .A3(G384), .A4(G381), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1023), .A3(new_n1234), .A4(new_n1236), .ZN(G407));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(G343), .C2(new_n1238), .ZN(G409));
  AND2_X1   g1039(.A1(new_n698), .A2(G213), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1117), .A2(new_n1141), .A3(new_n1191), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1194), .B2(new_n971), .ZN(new_n1242));
  OAI21_X1  g1042(.A(KEYINPUT124), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1198), .A2(new_n1200), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n755), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1240), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1240), .A2(G2897), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1092), .B2(new_n1099), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1113), .A2(new_n1112), .A3(KEYINPUT60), .A4(new_n1097), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(new_n721), .A3(new_n1100), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1221), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(G384), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT125), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1250), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1255), .B1(new_n828), .B2(new_n856), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G384), .B1(new_n1254), .B2(new_n1221), .ZN(new_n1260));
  OAI211_X1 g1060(.A(KEYINPUT125), .B(new_n1249), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1258), .A2(new_n1261), .B1(new_n1257), .B2(new_n1256), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1248), .B2(new_n1262), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1247), .B(new_n1256), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT62), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G375), .A2(G378), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1256), .A4(new_n1247), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1263), .A2(new_n1265), .A3(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(G393), .B(new_n819), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1064), .A2(new_n1089), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1058), .B2(new_n754), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1274), .A2(new_n1022), .A3(new_n994), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n994), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G390), .B1(new_n1276), .B2(new_n1021), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1271), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1023), .A2(G390), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1274), .B1(new_n1022), .B2(new_n994), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1270), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1269), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1278), .A2(new_n1284), .A3(new_n1281), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1264), .B2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1256), .A4(new_n1247), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1248), .A2(new_n1262), .A3(KEYINPUT126), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT126), .B1(new_n1248), .B2(new_n1262), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1287), .B(new_n1288), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1283), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1283), .A2(new_n1291), .A3(KEYINPUT127), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G405));
  NAND2_X1  g1096(.A1(new_n1266), .A2(new_n1238), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1297), .B(new_n1256), .ZN(new_n1298));
  XOR2_X1   g1098(.A(new_n1298), .B(new_n1282), .Z(G402));
endmodule


