

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747;

  XNOR2_X1 U378 ( .A(n596), .B(n595), .ZN(n744) );
  XNOR2_X1 U379 ( .A(n424), .B(G110), .ZN(n423) );
  XNOR2_X2 U380 ( .A(n734), .B(n400), .ZN(n649) );
  XNOR2_X2 U381 ( .A(n383), .B(n591), .ZN(n594) );
  OR2_X2 U382 ( .A1(n714), .A2(n384), .ZN(n383) );
  NOR2_X2 U383 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X2 U384 ( .A(n417), .B(n416), .ZN(n745) );
  XNOR2_X2 U385 ( .A(n576), .B(n575), .ZN(n628) );
  NOR2_X2 U386 ( .A1(n747), .A2(n745), .ZN(n415) );
  XNOR2_X1 U387 ( .A(G116), .B(G113), .ZN(n463) );
  NAND2_X1 U388 ( .A1(n562), .A2(n561), .ZN(n679) );
  XNOR2_X1 U389 ( .A(G146), .B(KEYINPUT65), .ZN(n470) );
  INV_X2 U390 ( .A(G953), .ZN(n736) );
  AND2_X1 U391 ( .A1(n387), .A2(n361), .ZN(n402) );
  XNOR2_X1 U392 ( .A(n404), .B(n388), .ZN(n387) );
  XNOR2_X1 U393 ( .A(n538), .B(KEYINPUT74), .ZN(n660) );
  INV_X2 U394 ( .A(n619), .ZN(n605) );
  INV_X1 U395 ( .A(KEYINPUT16), .ZN(n391) );
  AND2_X1 U396 ( .A1(n711), .A2(n514), .ZN(n437) );
  NAND2_X1 U397 ( .A1(n574), .A2(n676), .ZN(n576) );
  XNOR2_X1 U398 ( .A(n402), .B(n401), .ZN(n407) );
  XNOR2_X1 U399 ( .A(KEYINPUT107), .B(n565), .ZN(n747) );
  NOR2_X1 U400 ( .A1(n683), .A2(n660), .ZN(n539) );
  XNOR2_X1 U401 ( .A(n431), .B(KEYINPUT42), .ZN(n565) );
  AND2_X1 U402 ( .A1(n618), .A2(n372), .ZN(n567) );
  XNOR2_X1 U403 ( .A(n534), .B(n533), .ZN(n558) );
  XNOR2_X1 U404 ( .A(n425), .B(n358), .ZN(n400) );
  XNOR2_X1 U405 ( .A(n394), .B(n357), .ZN(n464) );
  XNOR2_X1 U406 ( .A(n395), .B(n463), .ZN(n394) );
  XNOR2_X1 U407 ( .A(n481), .B(n480), .ZN(n502) );
  XNOR2_X1 U408 ( .A(n423), .B(n465), .ZN(n531) );
  XNOR2_X1 U409 ( .A(n470), .B(KEYINPUT4), .ZN(n501) );
  XNOR2_X1 U410 ( .A(n391), .B(G122), .ZN(n390) );
  INV_X1 U411 ( .A(G101), .ZN(n460) );
  INV_X1 U412 ( .A(KEYINPUT32), .ZN(n401) );
  INV_X2 U413 ( .A(KEYINPUT70), .ZN(n424) );
  XNOR2_X1 U414 ( .A(G104), .B(G107), .ZN(n465) );
  NOR2_X1 U415 ( .A1(KEYINPUT44), .A2(KEYINPUT81), .ZN(n608) );
  XNOR2_X2 U416 ( .A(n374), .B(n366), .ZN(n688) );
  XNOR2_X1 U417 ( .A(n531), .B(n390), .ZN(n389) );
  XNOR2_X1 U418 ( .A(n501), .B(n500), .ZN(n503) );
  INV_X1 U419 ( .A(G131), .ZN(n499) );
  AND2_X1 U420 ( .A1(n604), .A2(n546), .ZN(n615) );
  XNOR2_X1 U421 ( .A(n382), .B(G140), .ZN(n733) );
  XNOR2_X1 U422 ( .A(G125), .B(KEYINPUT10), .ZN(n382) );
  INV_X1 U423 ( .A(G469), .ZN(n533) );
  XNOR2_X1 U424 ( .A(n733), .B(n370), .ZN(n513) );
  INV_X1 U425 ( .A(G146), .ZN(n370) );
  AND2_X1 U426 ( .A1(n368), .A2(n614), .ZN(n582) );
  XNOR2_X1 U427 ( .A(n615), .B(n369), .ZN(n368) );
  INV_X1 U428 ( .A(KEYINPUT22), .ZN(n388) );
  NOR2_X1 U429 ( .A1(n393), .A2(n392), .ZN(n442) );
  AND2_X1 U430 ( .A1(n736), .A2(G227), .ZN(n421) );
  XNOR2_X1 U431 ( .A(n530), .B(G140), .ZN(n422) );
  INV_X1 U432 ( .A(KEYINPUT88), .ZN(n530) );
  XNOR2_X1 U433 ( .A(KEYINPUT87), .B(KEYINPUT18), .ZN(n466) );
  XOR2_X1 U434 ( .A(G125), .B(KEYINPUT71), .Z(n467) );
  NOR2_X1 U435 ( .A1(n679), .A2(n376), .ZN(n375) );
  NAND2_X1 U436 ( .A1(n462), .A2(n461), .ZN(n395) );
  XNOR2_X1 U437 ( .A(n450), .B(n449), .ZN(n448) );
  XNOR2_X1 U438 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n450) );
  XNOR2_X1 U439 ( .A(G119), .B(G110), .ZN(n449) );
  XNOR2_X1 U440 ( .A(n381), .B(n379), .ZN(n511) );
  XNOR2_X1 U441 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n381) );
  NOR2_X1 U442 ( .A1(n380), .A2(G953), .ZN(n379) );
  INV_X1 U443 ( .A(G234), .ZN(n380) );
  INV_X1 U444 ( .A(G134), .ZN(n480) );
  XNOR2_X1 U445 ( .A(G116), .B(G122), .ZN(n476) );
  XOR2_X1 U446 ( .A(KEYINPUT97), .B(G107), .Z(n477) );
  XOR2_X1 U447 ( .A(n491), .B(n513), .Z(n637) );
  XNOR2_X1 U448 ( .A(KEYINPUT1), .B(KEYINPUT64), .ZN(n440) );
  XNOR2_X1 U449 ( .A(n386), .B(KEYINPUT103), .ZN(n385) );
  AND2_X1 U450 ( .A1(n549), .A2(n548), .ZN(n372) );
  INV_X1 U451 ( .A(n547), .ZN(n548) );
  XNOR2_X1 U452 ( .A(n446), .B(n517), .ZN(n606) );
  OR2_X1 U453 ( .A1(n720), .A2(G902), .ZN(n446) );
  INV_X1 U454 ( .A(KEYINPUT0), .ZN(n414) );
  NOR2_X1 U455 ( .A1(n588), .A2(n706), .ZN(n451) );
  NOR2_X1 U456 ( .A1(n716), .A2(G902), .ZN(n482) );
  XNOR2_X1 U457 ( .A(n619), .B(n452), .ZN(n614) );
  XNOR2_X1 U458 ( .A(KEYINPUT98), .B(KEYINPUT6), .ZN(n452) );
  NAND2_X1 U459 ( .A1(n435), .A2(n434), .ZN(n412) );
  AND2_X1 U460 ( .A1(n713), .A2(n365), .ZN(n434) );
  INV_X1 U461 ( .A(KEYINPUT77), .ZN(n397) );
  INV_X1 U462 ( .A(KEYINPUT48), .ZN(n441) );
  NAND2_X1 U463 ( .A1(G234), .A2(G237), .ZN(n518) );
  NAND2_X1 U464 ( .A1(G953), .A2(G902), .ZN(n585) );
  XOR2_X1 U465 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n506) );
  INV_X1 U466 ( .A(KEYINPUT67), .ZN(n459) );
  XNOR2_X1 U467 ( .A(G143), .B(G113), .ZN(n483) );
  XOR2_X1 U468 ( .A(G104), .B(G122), .Z(n484) );
  XNOR2_X1 U469 ( .A(G131), .B(KEYINPUT11), .ZN(n485) );
  XOR2_X1 U470 ( .A(KEYINPUT96), .B(KEYINPUT12), .Z(n486) );
  NOR2_X1 U471 ( .A1(G953), .A2(G237), .ZN(n504) );
  INV_X1 U472 ( .A(KEYINPUT101), .ZN(n369) );
  OR2_X1 U473 ( .A1(G237), .A2(G902), .ZN(n497) );
  XNOR2_X1 U474 ( .A(n531), .B(n420), .ZN(n532) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n727), .B(n468), .ZN(n475) );
  XNOR2_X1 U477 ( .A(n399), .B(n398), .ZN(n710) );
  INV_X1 U478 ( .A(KEYINPUT78), .ZN(n398) );
  XNOR2_X1 U479 ( .A(n373), .B(n419), .ZN(n618) );
  INV_X1 U480 ( .A(KEYINPUT92), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n371), .B(n513), .ZN(n720) );
  XNOR2_X1 U482 ( .A(n447), .B(n512), .ZN(n371) );
  XNOR2_X1 U483 ( .A(n510), .B(n448), .ZN(n447) );
  AND2_X2 U484 ( .A1(n437), .A2(n632), .ZN(n718) );
  XNOR2_X1 U485 ( .A(n378), .B(n377), .ZN(n716) );
  XNOR2_X1 U486 ( .A(n479), .B(n359), .ZN(n377) );
  XNOR2_X1 U487 ( .A(n502), .B(n478), .ZN(n378) );
  NAND2_X1 U488 ( .A1(n718), .A2(G478), .ZN(n445) );
  NAND2_X1 U489 ( .A1(n718), .A2(G475), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n637), .B(n636), .ZN(n439) );
  INV_X1 U491 ( .A(KEYINPUT40), .ZN(n416) );
  XNOR2_X1 U492 ( .A(n569), .B(KEYINPUT108), .ZN(n556) );
  INV_X1 U493 ( .A(n697), .ZN(n413) );
  NOR2_X1 U494 ( .A1(n613), .A2(n614), .ZN(n651) );
  INV_X1 U495 ( .A(KEYINPUT53), .ZN(n409) );
  XNOR2_X1 U496 ( .A(n558), .B(n440), .ZN(n604) );
  XNOR2_X1 U497 ( .A(G119), .B(KEYINPUT3), .ZN(n357) );
  XOR2_X1 U498 ( .A(n506), .B(n505), .Z(n358) );
  XNOR2_X1 U499 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n359) );
  AND2_X1 U500 ( .A1(n561), .A2(n543), .ZN(n360) );
  NAND2_X1 U501 ( .A1(n606), .A2(n598), .ZN(n691) );
  AND2_X1 U502 ( .A1(n603), .A2(n432), .ZN(n361) );
  AND2_X1 U503 ( .A1(n619), .A2(n618), .ZN(n362) );
  AND2_X1 U504 ( .A1(n552), .A2(KEYINPUT47), .ZN(n363) );
  INV_X1 U505 ( .A(n604), .ZN(n692) );
  NOR2_X1 U506 ( .A1(n363), .A2(n664), .ZN(n364) );
  OR2_X1 U507 ( .A1(n715), .A2(n714), .ZN(n365) );
  XOR2_X1 U508 ( .A(n563), .B(KEYINPUT106), .Z(n366) );
  XNOR2_X1 U509 ( .A(n464), .B(n389), .ZN(n727) );
  NAND2_X1 U510 ( .A1(n367), .A2(n623), .ZN(n624) );
  NAND2_X1 U511 ( .A1(n611), .A2(n403), .ZN(n367) );
  NOR2_X1 U512 ( .A1(G902), .A2(n642), .ZN(n534) );
  NAND2_X1 U513 ( .A1(n546), .A2(n558), .ZN(n373) );
  INV_X1 U514 ( .A(n679), .ZN(n599) );
  NAND2_X1 U515 ( .A1(n375), .A2(n566), .ZN(n374) );
  INV_X1 U516 ( .A(n680), .ZN(n376) );
  INV_X1 U517 ( .A(n601), .ZN(n384) );
  XNOR2_X1 U518 ( .A(n582), .B(n583), .ZN(n714) );
  NAND2_X1 U519 ( .A1(n385), .A2(n360), .ZN(n569) );
  NAND2_X1 U520 ( .A1(n555), .A2(n614), .ZN(n386) );
  NAND2_X1 U521 ( .A1(n553), .A2(n673), .ZN(n393) );
  NAND2_X1 U522 ( .A1(n559), .A2(n604), .ZN(n673) );
  AND2_X1 U523 ( .A1(n387), .A2(n692), .ZN(n612) );
  NAND2_X1 U524 ( .A1(n396), .A2(n364), .ZN(n392) );
  OR2_X1 U525 ( .A1(KEYINPUT44), .A2(n744), .ZN(n611) );
  NAND2_X1 U526 ( .A1(n625), .A2(n708), .ZN(n711) );
  XNOR2_X1 U527 ( .A(n430), .B(n439), .ZN(n429) );
  XNOR2_X1 U528 ( .A(n581), .B(KEYINPUT79), .ZN(n625) );
  XNOR2_X1 U529 ( .A(n445), .B(n444), .ZN(n405) );
  NAND2_X1 U530 ( .A1(n628), .A2(n580), .ZN(n581) );
  XNOR2_X1 U531 ( .A(n436), .B(n397), .ZN(n396) );
  NAND2_X1 U532 ( .A1(n629), .A2(n630), .ZN(n399) );
  NOR2_X1 U533 ( .A1(n709), .A2(n710), .ZN(n712) );
  NAND2_X1 U534 ( .A1(n429), .A2(n717), .ZN(n428) );
  NAND2_X1 U535 ( .A1(n610), .A2(n744), .ZN(n403) );
  NAND2_X1 U536 ( .A1(n601), .A2(n600), .ZN(n404) );
  NAND2_X1 U537 ( .A1(n405), .A2(n717), .ZN(n443) );
  NOR2_X2 U538 ( .A1(G902), .A2(n649), .ZN(n508) );
  XNOR2_X1 U539 ( .A(n406), .B(n646), .ZN(G54) );
  NAND2_X1 U540 ( .A1(n645), .A2(n717), .ZN(n406) );
  NAND2_X1 U541 ( .A1(n442), .A2(n427), .ZN(n426) );
  NAND2_X1 U542 ( .A1(n407), .A2(n659), .ZN(n609) );
  XNOR2_X1 U543 ( .A(n407), .B(G119), .ZN(G21) );
  XNOR2_X1 U544 ( .A(n408), .B(KEYINPUT19), .ZN(n433) );
  NOR2_X1 U545 ( .A1(n556), .A2(n408), .ZN(n557) );
  XNOR2_X2 U546 ( .A(n498), .B(KEYINPUT82), .ZN(n408) );
  XNOR2_X1 U547 ( .A(n410), .B(n409), .ZN(G75) );
  NAND2_X1 U548 ( .A1(n411), .A2(n736), .ZN(n410) );
  XNOR2_X1 U549 ( .A(n412), .B(KEYINPUT119), .ZN(n411) );
  AND2_X1 U550 ( .A1(n601), .A2(n413), .ZN(n617) );
  AND2_X1 U551 ( .A1(n601), .A2(n362), .ZN(n656) );
  XNOR2_X2 U552 ( .A(n590), .B(n414), .ZN(n601) );
  XNOR2_X1 U553 ( .A(n415), .B(KEYINPUT46), .ZN(n427) );
  NAND2_X1 U554 ( .A1(n577), .A2(n360), .ZN(n417) );
  NAND2_X1 U555 ( .A1(n418), .A2(n708), .ZN(n631) );
  INV_X1 U556 ( .A(n629), .ZN(n418) );
  XNOR2_X1 U557 ( .A(n629), .B(n738), .ZN(n737) );
  INV_X1 U558 ( .A(n464), .ZN(n425) );
  XNOR2_X1 U559 ( .A(n426), .B(n441), .ZN(n574) );
  XNOR2_X1 U560 ( .A(n428), .B(n638), .ZN(G60) );
  NAND2_X1 U561 ( .A1(n688), .A2(n564), .ZN(n431) );
  INV_X1 U562 ( .A(n689), .ZN(n432) );
  NAND2_X1 U563 ( .A1(n433), .A2(n564), .ZN(n538) );
  NAND2_X1 U564 ( .A1(n433), .A2(n451), .ZN(n590) );
  NAND2_X1 U565 ( .A1(n712), .A2(n711), .ZN(n435) );
  NAND2_X1 U566 ( .A1(n660), .A2(KEYINPUT47), .ZN(n436) );
  XNOR2_X1 U567 ( .A(n443), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U568 ( .A(n734), .B(n438), .ZN(n642) );
  XNOR2_X2 U569 ( .A(n502), .B(n503), .ZN(n734) );
  XNOR2_X1 U570 ( .A(n532), .B(G101), .ZN(n438) );
  XNOR2_X2 U571 ( .A(G128), .B(KEYINPUT75), .ZN(n469) );
  INV_X1 U572 ( .A(n716), .ZN(n444) );
  INV_X1 U573 ( .A(n606), .ZN(n602) );
  XNOR2_X2 U574 ( .A(n469), .B(G143), .ZN(n481) );
  XNOR2_X2 U575 ( .A(n508), .B(n507), .ZN(n619) );
  NAND2_X1 U576 ( .A1(n453), .A2(n717), .ZN(n635) );
  XNOR2_X1 U577 ( .A(n455), .B(n454), .ZN(n453) );
  XNOR2_X1 U578 ( .A(n633), .B(KEYINPUT54), .ZN(n454) );
  NAND2_X1 U579 ( .A1(n718), .A2(G210), .ZN(n455) );
  XNOR2_X1 U580 ( .A(n456), .B(n650), .ZN(G57) );
  NAND2_X1 U581 ( .A1(n457), .A2(n717), .ZN(n456) );
  XNOR2_X1 U582 ( .A(n647), .B(n458), .ZN(n457) );
  XNOR2_X1 U583 ( .A(n649), .B(n648), .ZN(n458) );
  XNOR2_X1 U584 ( .A(n499), .B(G137), .ZN(n500) );
  INV_X1 U585 ( .A(KEYINPUT80), .ZN(n575) );
  INV_X1 U586 ( .A(KEYINPUT41), .ZN(n563) );
  XNOR2_X1 U587 ( .A(n481), .B(n473), .ZN(n474) );
  INV_X1 U588 ( .A(n743), .ZN(n627) );
  AND2_X1 U589 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U590 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U591 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X1 U592 ( .A1(n736), .A2(G952), .ZN(n722) );
  NAND2_X1 U593 ( .A1(G101), .A2(n459), .ZN(n462) );
  NAND2_X1 U594 ( .A1(n460), .A2(KEYINPUT67), .ZN(n461) );
  XNOR2_X1 U595 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U596 ( .A(n501), .B(KEYINPUT17), .Z(n472) );
  NAND2_X1 U597 ( .A1(G224), .A2(n736), .ZN(n471) );
  XNOR2_X1 U598 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U599 ( .A(n475), .B(n474), .ZN(n494) );
  XNOR2_X1 U600 ( .A(n494), .B(KEYINPUT55), .ZN(n633) );
  XNOR2_X1 U601 ( .A(n477), .B(n476), .ZN(n479) );
  NAND2_X1 U602 ( .A1(G217), .A2(n511), .ZN(n478) );
  XNOR2_X1 U603 ( .A(G478), .B(n482), .ZN(n561) );
  XNOR2_X1 U604 ( .A(KEYINPUT13), .B(G475), .ZN(n493) );
  XNOR2_X1 U605 ( .A(n484), .B(n483), .ZN(n488) );
  XNOR2_X1 U606 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U607 ( .A(n488), .B(n487), .Z(n490) );
  NAND2_X1 U608 ( .A1(n504), .A2(G214), .ZN(n489) );
  XNOR2_X1 U609 ( .A(n490), .B(n489), .ZN(n491) );
  NOR2_X1 U610 ( .A1(G902), .A2(n637), .ZN(n492) );
  XNOR2_X1 U611 ( .A(n493), .B(n492), .ZN(n543) );
  NOR2_X1 U612 ( .A1(n543), .A2(n561), .ZN(n669) );
  NOR2_X1 U613 ( .A1(n360), .A2(n669), .ZN(n683) );
  XOR2_X1 U614 ( .A(G902), .B(KEYINPUT15), .Z(n514) );
  NOR2_X1 U615 ( .A1(n514), .A2(n494), .ZN(n496) );
  NAND2_X1 U616 ( .A1(G210), .A2(n497), .ZN(n495) );
  XNOR2_X1 U617 ( .A(n496), .B(n495), .ZN(n542) );
  NAND2_X1 U618 ( .A1(G214), .A2(n497), .ZN(n680) );
  NAND2_X1 U619 ( .A1(n542), .A2(n680), .ZN(n498) );
  NAND2_X1 U620 ( .A1(n504), .A2(G210), .ZN(n505) );
  XNOR2_X1 U621 ( .A(KEYINPUT94), .B(G472), .ZN(n507) );
  XNOR2_X1 U622 ( .A(G128), .B(G137), .ZN(n509) );
  XNOR2_X1 U623 ( .A(n509), .B(KEYINPUT89), .ZN(n510) );
  NAND2_X1 U624 ( .A1(G221), .A2(n511), .ZN(n512) );
  INV_X1 U625 ( .A(n514), .ZN(n626) );
  NAND2_X1 U626 ( .A1(G234), .A2(n626), .ZN(n515) );
  XNOR2_X1 U627 ( .A(KEYINPUT20), .B(n515), .ZN(n523) );
  NAND2_X1 U628 ( .A1(n523), .A2(G217), .ZN(n516) );
  XOR2_X1 U629 ( .A(KEYINPUT25), .B(n516), .Z(n517) );
  XNOR2_X1 U630 ( .A(n518), .B(KEYINPUT14), .ZN(n589) );
  NOR2_X1 U631 ( .A1(G900), .A2(n585), .ZN(n519) );
  NAND2_X1 U632 ( .A1(n589), .A2(n519), .ZN(n520) );
  XOR2_X1 U633 ( .A(KEYINPUT102), .B(n520), .Z(n522) );
  INV_X1 U634 ( .A(n589), .ZN(n706) );
  NAND2_X1 U635 ( .A1(n736), .A2(G952), .ZN(n584) );
  NOR2_X1 U636 ( .A1(n706), .A2(n584), .ZN(n521) );
  NOR2_X1 U637 ( .A1(n522), .A2(n521), .ZN(n547) );
  XOR2_X1 U638 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n525) );
  NAND2_X1 U639 ( .A1(n523), .A2(G221), .ZN(n524) );
  XNOR2_X1 U640 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U641 ( .A(KEYINPUT90), .B(n526), .ZN(n597) );
  NOR2_X1 U642 ( .A1(n547), .A2(n597), .ZN(n527) );
  NAND2_X1 U643 ( .A1(n602), .A2(n527), .ZN(n554) );
  NOR2_X1 U644 ( .A1(n619), .A2(n554), .ZN(n529) );
  XNOR2_X1 U645 ( .A(KEYINPUT105), .B(KEYINPUT28), .ZN(n528) );
  XNOR2_X1 U646 ( .A(n529), .B(n528), .ZN(n537) );
  INV_X1 U647 ( .A(n558), .ZN(n535) );
  XNOR2_X1 U648 ( .A(KEYINPUT104), .B(n535), .ZN(n536) );
  NOR2_X1 U649 ( .A1(n537), .A2(n536), .ZN(n564) );
  XNOR2_X1 U650 ( .A(n539), .B(KEYINPUT68), .ZN(n541) );
  INV_X1 U651 ( .A(KEYINPUT47), .ZN(n540) );
  NAND2_X1 U652 ( .A1(n541), .A2(n540), .ZN(n553) );
  INV_X1 U653 ( .A(n542), .ZN(n572) );
  INV_X1 U654 ( .A(n543), .ZN(n562) );
  NOR2_X1 U655 ( .A1(n562), .A2(n561), .ZN(n592) );
  INV_X1 U656 ( .A(KEYINPUT30), .ZN(n545) );
  NAND2_X1 U657 ( .A1(n680), .A2(n605), .ZN(n544) );
  XNOR2_X1 U658 ( .A(n545), .B(n544), .ZN(n549) );
  INV_X1 U659 ( .A(n691), .ZN(n546) );
  NAND2_X1 U660 ( .A1(n592), .A2(n567), .ZN(n550) );
  NOR2_X1 U661 ( .A1(n572), .A2(n550), .ZN(n664) );
  INV_X1 U662 ( .A(n683), .ZN(n551) );
  NAND2_X1 U663 ( .A1(KEYINPUT68), .A2(n551), .ZN(n552) );
  INV_X1 U664 ( .A(n554), .ZN(n555) );
  XNOR2_X1 U665 ( .A(n557), .B(KEYINPUT36), .ZN(n559) );
  XOR2_X1 U666 ( .A(KEYINPUT69), .B(KEYINPUT38), .Z(n560) );
  XNOR2_X1 U667 ( .A(n572), .B(n560), .ZN(n566) );
  BUF_X1 U668 ( .A(n566), .Z(n681) );
  NAND2_X1 U669 ( .A1(n567), .A2(n681), .ZN(n568) );
  XNOR2_X2 U670 ( .A(n568), .B(KEYINPUT39), .ZN(n577) );
  NOR2_X1 U671 ( .A1(n604), .A2(n569), .ZN(n570) );
  NAND2_X1 U672 ( .A1(n570), .A2(n680), .ZN(n571) );
  XNOR2_X1 U673 ( .A(n571), .B(KEYINPUT43), .ZN(n573) );
  NAND2_X1 U674 ( .A1(n573), .A2(n572), .ZN(n676) );
  INV_X1 U675 ( .A(KEYINPUT2), .ZN(n630) );
  NAND2_X1 U676 ( .A1(n577), .A2(n669), .ZN(n578) );
  XNOR2_X1 U677 ( .A(KEYINPUT109), .B(n578), .ZN(n743) );
  OR2_X1 U678 ( .A1(n630), .A2(n743), .ZN(n579) );
  XOR2_X1 U679 ( .A(KEYINPUT76), .B(n579), .Z(n580) );
  XOR2_X1 U680 ( .A(KEYINPUT33), .B(KEYINPUT83), .Z(n583) );
  INV_X1 U681 ( .A(n584), .ZN(n587) );
  NOR2_X1 U682 ( .A1(G898), .A2(n585), .ZN(n586) );
  NOR2_X1 U683 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U684 ( .A(KEYINPUT34), .B(KEYINPUT73), .Z(n591) );
  INV_X1 U685 ( .A(n592), .ZN(n593) );
  XNOR2_X1 U686 ( .A(KEYINPUT35), .B(KEYINPUT72), .ZN(n595) );
  INV_X1 U687 ( .A(n597), .ZN(n598) );
  XNOR2_X1 U688 ( .A(n602), .B(KEYINPUT99), .ZN(n689) );
  NOR2_X1 U689 ( .A1(n692), .A2(n614), .ZN(n603) );
  NOR2_X1 U690 ( .A1(n605), .A2(n606), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n612), .A2(n607), .ZN(n659) );
  XNOR2_X1 U692 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n612), .A2(n689), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n615), .A2(n605), .ZN(n697) );
  XNOR2_X1 U695 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n617), .B(n616), .ZN(n670) );
  NOR2_X1 U697 ( .A1(n670), .A2(n656), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n683), .A2(n620), .ZN(n621) );
  NOR2_X1 U699 ( .A1(n651), .A2(n621), .ZN(n622) );
  XNOR2_X1 U700 ( .A(KEYINPUT100), .B(n622), .ZN(n623) );
  XNOR2_X2 U701 ( .A(n624), .B(KEYINPUT45), .ZN(n708) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n632) );
  INV_X1 U704 ( .A(n722), .ZN(n717) );
  INV_X1 U705 ( .A(KEYINPUT56), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(G51) );
  XOR2_X1 U707 ( .A(KEYINPUT59), .B(KEYINPUT85), .Z(n636) );
  INV_X1 U708 ( .A(KEYINPUT60), .ZN(n638) );
  INV_X1 U709 ( .A(KEYINPUT122), .ZN(n646) );
  NAND2_X1 U710 ( .A1(n718), .A2(G469), .ZN(n644) );
  XOR2_X1 U711 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n640) );
  XNOR2_X1 U712 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n641) );
  XOR2_X1 U714 ( .A(KEYINPUT62), .B(KEYINPUT84), .Z(n648) );
  NAND2_X1 U715 ( .A1(n718), .A2(G472), .ZN(n647) );
  XNOR2_X1 U716 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n650) );
  XOR2_X1 U717 ( .A(n651), .B(G101), .Z(G3) );
  NAND2_X1 U718 ( .A1(n656), .A2(n360), .ZN(n652) );
  XNOR2_X1 U719 ( .A(n652), .B(G104), .ZN(G6) );
  XOR2_X1 U720 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n654) );
  XNOR2_X1 U721 ( .A(G107), .B(KEYINPUT26), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(n655) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(n655), .Z(n658) );
  NAND2_X1 U724 ( .A1(n656), .A2(n669), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n658), .B(n657), .ZN(G9) );
  XNOR2_X1 U726 ( .A(G110), .B(n659), .ZN(G12) );
  XOR2_X1 U727 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n662) );
  INV_X1 U728 ( .A(n660), .ZN(n665) );
  NAND2_X1 U729 ( .A1(n669), .A2(n665), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(G128), .B(n663), .ZN(G30) );
  XOR2_X1 U732 ( .A(G143), .B(n664), .Z(G45) );
  XOR2_X1 U733 ( .A(G146), .B(KEYINPUT113), .Z(n667) );
  NAND2_X1 U734 ( .A1(n360), .A2(n665), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(G48) );
  NAND2_X1 U736 ( .A1(n670), .A2(n360), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n668), .B(G113), .ZN(G15) );
  NAND2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n671), .B(KEYINPUT114), .ZN(n672) );
  XNOR2_X1 U740 ( .A(G116), .B(n672), .ZN(G18) );
  XNOR2_X1 U741 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U743 ( .A(G125), .B(n675), .ZN(G27) );
  XNOR2_X1 U744 ( .A(G140), .B(KEYINPUT116), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n677), .B(n676), .ZN(G42) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n685) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U751 ( .A1(n714), .A2(n686), .ZN(n687) );
  XNOR2_X1 U752 ( .A(KEYINPUT118), .B(n687), .ZN(n703) );
  INV_X1 U753 ( .A(n688), .ZN(n715) );
  NOR2_X1 U754 ( .A1(n598), .A2(n689), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n690), .B(KEYINPUT49), .ZN(n696) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U757 ( .A(KEYINPUT50), .B(n693), .Z(n694) );
  NOR2_X1 U758 ( .A1(n605), .A2(n694), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n700) );
  XOR2_X1 U761 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n699) );
  XNOR2_X1 U762 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n715), .A2(n701), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U765 ( .A(n704), .B(KEYINPUT52), .ZN(n705) );
  NOR2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U767 ( .A1(G952), .A2(n707), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n708), .A2(KEYINPUT2), .ZN(n709) );
  NAND2_X1 U769 ( .A1(G217), .A2(n718), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U771 ( .A1(n722), .A2(n721), .ZN(G66) );
  NAND2_X1 U772 ( .A1(n736), .A2(n708), .ZN(n726) );
  NAND2_X1 U773 ( .A1(G953), .A2(G224), .ZN(n723) );
  XNOR2_X1 U774 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U775 ( .A1(n724), .A2(G898), .ZN(n725) );
  NAND2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U777 ( .A1(G898), .A2(n736), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n727), .A2(n728), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(n732) );
  XOR2_X1 U780 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n731) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(G69) );
  XNOR2_X1 U782 ( .A(n734), .B(n733), .ZN(n735) );
  XOR2_X1 U783 ( .A(n735), .B(KEYINPUT126), .Z(n738) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(n742) );
  XNOR2_X1 U785 ( .A(G227), .B(n738), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U787 ( .A1(G953), .A2(n740), .ZN(n741) );
  NAND2_X1 U788 ( .A1(n742), .A2(n741), .ZN(G72) );
  XOR2_X1 U789 ( .A(G134), .B(n743), .Z(G36) );
  XNOR2_X1 U790 ( .A(G122), .B(n744), .ZN(G24) );
  XNOR2_X1 U791 ( .A(G131), .B(KEYINPUT127), .ZN(n746) );
  XNOR2_X1 U792 ( .A(n746), .B(n745), .ZN(G33) );
  XOR2_X1 U793 ( .A(n747), .B(G137), .Z(G39) );
endmodule

