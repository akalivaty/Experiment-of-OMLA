//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT68), .A2(G119), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT68), .A2(G119), .ZN(new_n196));
  OAI21_X1  g010(.A(G128), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT24), .B(G110), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OR3_X1    g017(.A1(new_n201), .A2(KEYINPUT80), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT80), .B1(new_n201), .B2(new_n203), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n195), .A2(new_n196), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n208), .B1(new_n201), .B2(new_n206), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n204), .B(new_n205), .C1(G110), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G140), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT77), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G140), .ZN(new_n215));
  AND4_X1   g029(.A1(KEYINPUT77), .A2(new_n213), .A3(new_n215), .A4(G125), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n211), .A2(KEYINPUT76), .A3(G140), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(KEYINPUT76), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n217), .B(G146), .C1(new_n213), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(KEYINPUT78), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n215), .A2(G125), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n211), .A2(G140), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT76), .ZN(new_n228));
  OR3_X1    g042(.A1(new_n211), .A2(KEYINPUT76), .A3(G140), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n213), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT77), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n226), .B2(KEYINPUT16), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n212), .A2(KEYINPUT77), .A3(new_n213), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n222), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT79), .ZN(new_n236));
  INV_X1    g050(.A(new_n230), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT78), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G146), .A4(new_n217), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n240), .B(new_n222), .C1(new_n230), .C2(new_n234), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n225), .A2(new_n236), .A3(new_n239), .A4(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n209), .A2(G110), .B1(new_n201), .B2(new_n203), .ZN(new_n243));
  AOI221_X4 g057(.A(new_n194), .B1(new_n210), .B2(new_n224), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n243), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n210), .A2(new_n224), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n193), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT25), .B1(new_n248), .B2(new_n188), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n250));
  NOR4_X1   g064(.A1(new_n244), .A2(new_n247), .A3(new_n250), .A4(G902), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n189), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n245), .A2(new_n246), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n194), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n245), .A2(new_n246), .A3(new_n193), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n188), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n250), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n257), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT81), .A3(new_n189), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n189), .A2(G902), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n248), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n254), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G237), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n191), .A3(G210), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n267), .B(KEYINPUT27), .Z(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n198), .B2(G116), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n207), .B2(G116), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n198), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT68), .A2(G119), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n276), .A2(KEYINPUT69), .A3(G116), .A4(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n271), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT2), .A2(G113), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT67), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT2), .A2(G113), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n276), .A2(G116), .A3(new_n277), .ZN(new_n285));
  INV_X1    g099(.A(new_n273), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT70), .A3(new_n278), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n280), .A2(new_n284), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n278), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n282), .A3(new_n283), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n222), .A2(G143), .ZN(new_n293));
  INV_X1    g107(.A(G143), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G146), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT0), .A4(G128), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G143), .B(G146), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(KEYINPUT64), .A3(KEYINPUT0), .A4(G128), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n299), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT0), .B(G128), .Z(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n306));
  INV_X1    g120(.A(G134), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT11), .B1(new_n307), .B2(G137), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT11), .ZN(new_n309));
  INV_X1    g123(.A(G137), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G134), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n308), .A2(new_n311), .B1(new_n307), .B2(G137), .ZN(new_n312));
  INV_X1    g126(.A(G131), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n298), .A2(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n306), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT66), .ZN(new_n319));
  AOI21_X1  g133(.A(G128), .B1(new_n293), .B2(new_n295), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n294), .A2(KEYINPUT1), .A3(G146), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n321), .B(KEYINPUT66), .C1(new_n299), .C2(G128), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n299), .A2(new_n325), .A3(G128), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n312), .A2(new_n313), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n310), .B2(G134), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n307), .B2(G137), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n329), .A2(new_n310), .A3(G134), .ZN(new_n332));
  OAI21_X1  g146(.A(G131), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n292), .A2(new_n318), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n289), .A2(new_n291), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n312), .B(G131), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n334), .B1(new_n338), .B2(new_n305), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n292), .A2(new_n318), .A3(KEYINPUT28), .A4(new_n334), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n270), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n318), .A2(KEYINPUT30), .A3(new_n334), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n344));
  INV_X1    g158(.A(new_n334), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n338), .A2(new_n305), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n337), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n270), .A3(new_n335), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT31), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n348), .A2(KEYINPUT31), .A3(new_n270), .A4(new_n335), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n342), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n354));
  NOR2_X1   g168(.A1(G472), .A2(G902), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT72), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(new_n335), .ZN(new_n358));
  INV_X1    g172(.A(new_n270), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n335), .A2(new_n336), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n339), .A2(new_n337), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n363), .A2(new_n270), .A3(new_n341), .A4(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n358), .A2(KEYINPUT74), .A3(new_n359), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n335), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n292), .B1(new_n334), .B2(new_n318), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT28), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT75), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT75), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n374), .B(KEYINPUT28), .C1(new_n370), .C2(new_n371), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n359), .A2(new_n366), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n373), .A2(new_n363), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n369), .A2(new_n188), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n357), .B1(new_n378), .B2(G472), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n351), .A2(new_n352), .ZN(new_n380));
  INV_X1    g194(.A(new_n342), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT73), .ZN(new_n383));
  INV_X1    g197(.A(new_n356), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT73), .B1(new_n353), .B2(new_n356), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n354), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n265), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(new_n389), .B2(G107), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G104), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(G107), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n390), .A2(new_n393), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n389), .A2(G107), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n392), .A2(G104), .ZN(new_n398));
  OAI21_X1  g212(.A(G101), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n291), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G113), .B1(new_n285), .B2(KEYINPUT5), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n290), .B2(KEYINPUT5), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT5), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n280), .B2(new_n288), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n291), .B1(new_n407), .B2(new_n403), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n405), .B1(new_n408), .B2(new_n400), .ZN(new_n409));
  XNOR2_X1  g223(.A(G110), .B(G122), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n410), .B(KEYINPUT8), .Z(new_n411));
  OAI21_X1  g225(.A(KEYINPUT87), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n413));
  INV_X1    g227(.A(new_n411), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n287), .A2(KEYINPUT70), .A3(new_n278), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT70), .B1(new_n287), .B2(new_n278), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT5), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n403), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n401), .B1(new_n419), .B2(new_n291), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n413), .B(new_n414), .C1(new_n420), .C2(new_n405), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n291), .A3(new_n401), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n390), .A2(new_n393), .A3(new_n395), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G101), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT4), .A3(new_n396), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n426), .A3(G101), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n289), .B2(new_n291), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n422), .A2(new_n410), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n323), .A2(new_n324), .A3(new_n211), .A4(new_n326), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n432), .A2(KEYINPUT86), .B1(new_n315), .B2(new_n211), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n191), .A2(G224), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT7), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n438), .A2(KEYINPUT88), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(KEYINPUT88), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n434), .A2(new_n435), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n435), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT88), .B(new_n438), .C1(new_n442), .C2(new_n433), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n412), .A2(new_n421), .A3(new_n431), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n188), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(KEYINPUT89), .A3(new_n188), .ZN(new_n449));
  INV_X1    g263(.A(new_n410), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n402), .B1(new_n417), .B2(new_n418), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n429), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n431), .A2(new_n452), .A3(KEYINPUT6), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n442), .A2(new_n433), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n436), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n450), .C1(new_n451), .C2(new_n429), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n453), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n449), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G210), .B1(G237), .B2(G902), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(KEYINPUT91), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n458), .B1(new_n446), .B2(new_n447), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(KEYINPUT90), .A3(new_n449), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n464), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n468), .A3(new_n449), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G214), .B1(G237), .B2(G902), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT9), .B(G234), .Z(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT82), .ZN(new_n473));
  OAI21_X1  g287(.A(G221), .B1(new_n473), .B2(G902), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n474), .B(KEYINPUT83), .Z(new_n475));
  INV_X1    g289(.A(G469), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n188), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G140), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n191), .A2(G227), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT10), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n400), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n327), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n321), .B1(new_n299), .B2(G128), .ZN(new_n484));
  AND4_X1   g298(.A1(new_n325), .A2(new_n293), .A3(new_n295), .A4(G128), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n481), .B1(new_n486), .B2(new_n400), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n428), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n306), .A3(new_n317), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n489), .A2(new_n491), .A3(new_n338), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n338), .B1(new_n489), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n480), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n491), .A3(new_n338), .ZN(new_n495));
  INV_X1    g309(.A(new_n480), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n323), .A2(new_n400), .A3(new_n324), .A4(new_n326), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n326), .B(new_n321), .C1(G128), .C2(new_n299), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n498), .A2(new_n499), .B1(new_n401), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n485), .B1(new_n484), .B2(new_n319), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n502), .A2(KEYINPUT85), .A3(new_n324), .A4(new_n400), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n497), .B(new_n338), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(new_n499), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n401), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT12), .B1(new_n507), .B2(new_n314), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n495), .B(new_n496), .C1(new_n504), .C2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n494), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n477), .B1(new_n510), .B2(new_n476), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n495), .B1(new_n504), .B2(new_n508), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n480), .B(KEYINPUT84), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n315), .B(KEYINPUT71), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n488), .B1(new_n515), .B2(new_n490), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n480), .B1(new_n516), .B2(new_n338), .ZN(new_n517));
  INV_X1    g331(.A(new_n493), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n512), .A2(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G469), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n475), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G475), .A2(G902), .ZN(new_n523));
  XNOR2_X1  g337(.A(G113), .B(G122), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(new_n389), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n266), .A2(new_n191), .A3(G214), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n294), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n266), .A2(new_n191), .A3(G143), .A4(G214), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT18), .A2(G131), .ZN(new_n530));
  OR3_X1    g344(.A1(new_n529), .A2(KEYINPUT93), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n529), .B2(KEYINPUT93), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n220), .A2(G146), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n223), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n529), .A2(G131), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n527), .A2(new_n313), .A3(new_n528), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT17), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(KEYINPUT17), .B2(new_n537), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n525), .B(new_n536), .C1(new_n242), .C2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n219), .A2(KEYINPUT19), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n228), .A2(new_n229), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n544), .B2(KEYINPUT19), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G146), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n230), .A2(new_n234), .A3(new_n222), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT94), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n221), .B(new_n549), .C1(G146), .C2(new_n545), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n537), .A2(new_n538), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n525), .B1(new_n552), .B2(new_n536), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n523), .B1(new_n542), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n536), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n221), .B1(new_n545), .B2(G146), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n559), .A2(KEYINPUT94), .B1(new_n537), .B2(new_n538), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n560), .B2(new_n550), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n541), .B1(new_n561), .B2(new_n525), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT20), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n523), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G478), .ZN(new_n566));
  NOR2_X1   g380(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G122), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(G116), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n574), .A2(KEYINPUT14), .ZN(new_n575));
  OR2_X1    g389(.A1(KEYINPUT95), .A2(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(KEYINPUT95), .A2(G122), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G116), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(KEYINPUT14), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G107), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n294), .A2(G128), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n199), .A2(KEYINPUT97), .A3(G143), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT97), .B1(new_n199), .B2(G143), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G134), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n586), .A2(G134), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n579), .A2(new_n589), .A3(new_n574), .ZN(new_n590));
  INV_X1    g404(.A(G116), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n576), .B2(new_n577), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT96), .B1(new_n592), .B2(new_n573), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI221_X1 g408(.A(new_n582), .B1(new_n587), .B2(new_n588), .C1(new_n594), .C2(G107), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n584), .A2(new_n585), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n583), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n294), .A2(KEYINPUT13), .A3(G128), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(G134), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n587), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n590), .A2(new_n593), .A3(G107), .ZN(new_n605));
  AOI21_X1  g419(.A(G107), .B1(new_n590), .B2(new_n593), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n595), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n473), .A2(new_n187), .A3(G953), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n595), .A2(new_n607), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n571), .B1(new_n613), .B2(new_n188), .ZN(new_n614));
  AOI211_X1 g428(.A(G902), .B(new_n570), .C1(new_n611), .C2(new_n612), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n191), .A2(G952), .ZN(new_n617));
  NAND2_X1  g431(.A1(G234), .A2(G237), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT21), .B(G898), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(G902), .A3(G953), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n536), .B1(new_n242), .B2(new_n540), .ZN(new_n624));
  INV_X1    g438(.A(new_n525), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n188), .B1(new_n626), .B2(new_n542), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G475), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n565), .A2(new_n616), .A3(new_n623), .A4(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n557), .A2(new_n564), .B1(new_n627), .B2(G475), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n632), .A2(KEYINPUT100), .A3(new_n623), .A4(new_n616), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n522), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n388), .A2(new_n470), .A3(new_n471), .A4(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT101), .B(G101), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G3));
  INV_X1    g451(.A(new_n449), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT89), .B1(new_n445), .B2(new_n188), .ZN(new_n639));
  NOR4_X1   g453(.A1(new_n638), .A2(new_n639), .A3(new_n464), .A4(new_n458), .ZN(new_n640));
  INV_X1    g454(.A(new_n471), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT102), .B1(new_n460), .B2(new_n464), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n469), .A2(new_n471), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n613), .A2(KEYINPUT33), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n611), .A2(new_n648), .A3(new_n612), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(G478), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n612), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n609), .B1(new_n595), .B2(new_n607), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n566), .B(new_n188), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(G478), .A2(G902), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n632), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n646), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n521), .A2(new_n254), .A3(new_n262), .A4(new_n264), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n353), .B2(G902), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n385), .A2(new_n386), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n657), .A2(new_n623), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NAND3_X1  g478(.A1(new_n562), .A2(new_n523), .A3(new_n555), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n557), .A2(new_n665), .B1(G475), .B2(new_n627), .ZN(new_n666));
  INV_X1    g480(.A(new_n616), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n468), .B1(new_n465), .B2(new_n449), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n471), .B(new_n469), .C1(new_n669), .C2(KEYINPUT102), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n668), .B1(new_n670), .B2(new_n643), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n623), .A3(new_n661), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NOR2_X1   g488(.A1(new_n194), .A2(KEYINPUT36), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n255), .B(new_n675), .Z(new_n676));
  OR3_X1    g490(.A1(new_n676), .A2(G902), .A3(new_n189), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n254), .A2(new_n262), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n660), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n470), .A2(new_n679), .A3(new_n471), .A4(new_n634), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  NAND3_X1  g496(.A1(new_n254), .A2(new_n262), .A3(new_n677), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n622), .A2(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n619), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n475), .B(new_n686), .C1(new_n511), .C2(new_n520), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n387), .B2(new_n379), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n671), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XNOR2_X1  g505(.A(new_n470), .B(KEYINPUT38), .ZN(new_n692));
  INV_X1    g506(.A(new_n357), .ZN(new_n693));
  INV_X1    g507(.A(G472), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n358), .A2(new_n270), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n370), .A2(new_n371), .A3(new_n270), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n696), .A2(G902), .A3(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n387), .B(new_n693), .C1(new_n694), .C2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n685), .B(KEYINPUT39), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n522), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT40), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT40), .B1(new_n522), .B2(new_n701), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n554), .A2(KEYINPUT20), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n555), .B1(new_n562), .B2(new_n523), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n628), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n667), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n683), .A2(new_n709), .A3(new_n641), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n704), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n692), .A2(new_n699), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND2_X1  g527(.A1(new_n657), .A2(new_n689), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  NAND3_X1  g529(.A1(new_n646), .A2(new_n623), .A3(new_n656), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n510), .A2(new_n476), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n510), .A2(new_n476), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n475), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n388), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  INV_X1    g538(.A(new_n668), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n646), .A2(new_n623), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n721), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT103), .B(G116), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G18));
  NAND2_X1  g543(.A1(new_n631), .A2(new_n633), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(new_n683), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n362), .A2(new_n367), .A3(new_n368), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n377), .A2(new_n188), .ZN(new_n733));
  OAI21_X1  g547(.A(G472), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n387), .A2(new_n693), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n646), .A3(new_n735), .A4(new_n720), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  AND3_X1   g551(.A1(new_n254), .A2(new_n262), .A3(new_n264), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n318), .A2(new_n334), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n337), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n336), .B1(new_n740), .B2(new_n335), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n741), .A2(new_n374), .B1(new_n336), .B2(new_n335), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n270), .B1(new_n742), .B2(new_n373), .ZN(new_n743));
  INV_X1    g557(.A(new_n380), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n384), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n745), .A2(new_n659), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n738), .A2(new_n746), .A3(new_n623), .A4(new_n720), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n709), .B1(new_n670), .B2(new_n643), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  INV_X1    g564(.A(new_n720), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n670), .B2(new_n643), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n745), .A2(new_n659), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n656), .A2(new_n685), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n678), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n752), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  AOI21_X1  g575(.A(new_n468), .B1(new_n460), .B2(new_n461), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n641), .B(new_n640), .C1(new_n762), .C2(new_n466), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n754), .A2(KEYINPUT42), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n388), .A3(new_n521), .A4(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n467), .A2(new_n471), .A3(new_n469), .A4(new_n521), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n354), .B1(new_n353), .B2(new_n356), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n734), .A2(new_n693), .A3(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n632), .A2(new_n655), .A3(new_n686), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n738), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT42), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT105), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n765), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n313), .ZN(G33));
  AOI21_X1  g591(.A(new_n640), .B1(new_n762), .B2(new_n466), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n388), .A2(new_n778), .A3(new_n471), .A4(new_n521), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n668), .A2(new_n686), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT106), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n766), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n388), .A4(new_n780), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NAND2_X1  g601(.A1(new_n653), .A2(new_n654), .ZN(new_n788));
  INV_X1    g602(.A(new_n649), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n648), .B1(new_n611), .B2(new_n612), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n788), .B1(new_n791), .B2(G478), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(new_n632), .B2(KEYINPUT110), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n565), .A2(KEYINPUT110), .A3(new_n628), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT43), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n708), .A2(new_n655), .A3(KEYINPUT43), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n796), .A2(new_n660), .A3(new_n798), .A4(new_n683), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n708), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n792), .A3(new_n794), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n797), .B1(new_n804), .B2(KEYINPUT43), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(KEYINPUT44), .A3(new_n660), .A4(new_n683), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n467), .A2(new_n471), .A3(new_n469), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT111), .B1(new_n778), .B2(new_n471), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n808), .A2(new_n809), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n778), .A2(KEYINPUT111), .A3(new_n471), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n801), .A2(new_n814), .A3(new_n806), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n512), .A2(new_n514), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n517), .A2(new_n518), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT45), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT107), .B1(new_n822), .B2(new_n476), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT107), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n824), .B(G469), .C1(new_n519), .C2(KEYINPUT45), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n519), .A2(KEYINPUT45), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT108), .ZN(new_n828));
  OAI21_X1  g642(.A(G469), .B1(new_n519), .B2(KEYINPUT45), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n829), .A2(KEYINPUT107), .B1(KEYINPUT45), .B2(new_n519), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT108), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n825), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n477), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT46), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n827), .A2(KEYINPUT108), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n831), .B1(new_n830), .B2(new_n825), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT46), .B(new_n834), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n718), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT109), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(KEYINPUT109), .A3(new_n718), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n475), .B(new_n701), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n819), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G137), .ZN(G39));
  NOR4_X1   g659(.A1(new_n808), .A2(new_n735), .A3(new_n738), .A4(new_n754), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT47), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n847), .B(new_n475), .C1(new_n841), .C2(new_n842), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT46), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n849), .B(new_n477), .C1(new_n828), .C2(new_n832), .ZN(new_n850));
  INV_X1    g664(.A(new_n718), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n840), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n835), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n842), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n475), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT47), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n846), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(G140), .ZN(G42));
  NOR2_X1   g672(.A1(new_n808), .A2(new_n751), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n699), .A2(new_n265), .A3(new_n619), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n632), .A3(new_n655), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n746), .A2(new_n683), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n619), .B(new_n797), .C1(new_n804), .C2(KEYINPUT43), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n265), .A2(new_n753), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n778), .B(KEYINPUT38), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n641), .A3(new_n720), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(KEYINPUT116), .A3(new_n641), .A4(new_n720), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n873), .B(new_n874), .C1(KEYINPUT117), .C2(KEYINPUT50), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n867), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n719), .A2(new_n855), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n848), .A2(new_n856), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n869), .A2(new_n810), .A3(new_n811), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT115), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n879), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n879), .B(KEYINPUT51), .C1(new_n881), .C2(new_n883), .ZN(new_n887));
  INV_X1    g701(.A(new_n752), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n617), .B1(new_n869), .B2(new_n888), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n738), .A2(new_n859), .A3(new_n768), .A4(new_n865), .ZN(new_n890));
  XOR2_X1   g704(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n889), .B(new_n892), .C1(new_n656), .C2(new_n862), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n886), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n721), .B1(new_n716), .B2(new_n726), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n635), .A2(new_n680), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n746), .A2(new_n683), .A3(new_n769), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n766), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n666), .A2(new_n616), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n689), .A2(new_n900), .A3(new_n763), .A4(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n718), .A2(new_n520), .A3(new_n834), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n855), .A3(new_n685), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT81), .B1(new_n261), .B2(new_n189), .ZN(new_n905));
  INV_X1    g719(.A(new_n189), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n253), .B(new_n906), .C1(new_n259), .C2(new_n260), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n908), .B2(new_n677), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n735), .A3(new_n901), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT113), .B1(new_n910), .B2(new_n808), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n899), .B1(new_n902), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n708), .A2(new_n655), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n632), .A2(new_n616), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n623), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n470), .A2(new_n661), .A3(new_n471), .A4(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n749), .A2(new_n736), .A3(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n897), .A2(new_n786), .A3(new_n912), .A4(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n776), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT53), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n689), .B(new_n646), .C1(new_n656), .C2(new_n725), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n748), .A2(new_n678), .A3(new_n687), .A4(new_n699), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n752), .A2(new_n758), .A3(new_n755), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n758), .B1(new_n752), .B2(new_n755), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n921), .B(new_n922), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT52), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n760), .A2(KEYINPUT52), .A3(new_n921), .A4(new_n922), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT114), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT114), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n925), .A2(new_n930), .A3(new_n926), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n919), .A2(new_n920), .A3(new_n929), .A4(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n927), .A2(new_n928), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n765), .A2(new_n771), .A3(new_n774), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n774), .B1(new_n765), .B2(new_n771), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n749), .A2(new_n736), .A3(new_n916), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n937), .A2(new_n895), .A3(new_n896), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n936), .A2(new_n938), .A3(new_n786), .A4(new_n912), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT53), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n932), .A2(new_n940), .A3(KEYINPUT54), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n920), .B1(new_n933), .B2(new_n939), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n786), .A2(new_n912), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n388), .A2(new_n720), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(new_n623), .C1(new_n657), .C2(new_n671), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n735), .A2(new_n730), .A3(new_n683), .ZN(new_n947));
  AOI22_X1  g761(.A1(new_n947), .A2(new_n752), .B1(new_n747), .B2(new_n748), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n778), .A2(new_n641), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(new_n634), .C1(new_n388), .C2(new_n679), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n946), .A2(new_n916), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n765), .A2(new_n771), .A3(KEYINPUT53), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n944), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n929), .A3(new_n931), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n942), .A2(new_n943), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n894), .A2(new_n957), .B1(G952), .B2(G953), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n738), .A2(new_n471), .A3(new_n855), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n719), .B(KEYINPUT49), .ZN(new_n960));
  NOR4_X1   g774(.A1(new_n959), .A2(new_n699), .A3(new_n960), .A4(new_n804), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n870), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n962), .ZN(G75));
  NOR2_X1   g777(.A1(new_n191), .A2(G952), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n188), .B1(new_n942), .B2(new_n954), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT56), .B1(new_n966), .B2(new_n464), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n453), .A2(new_n457), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(new_n455), .Z(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT55), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n965), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n967), .B2(new_n971), .ZN(G51));
  NAND2_X1  g787(.A1(new_n942), .A2(new_n954), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n974), .A2(G902), .A3(new_n832), .A4(new_n828), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT119), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n477), .B(KEYINPUT57), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n942), .A2(new_n943), .A3(new_n954), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n943), .B1(new_n942), .B2(new_n954), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n494), .A2(new_n509), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n964), .B1(new_n976), .B2(new_n982), .ZN(G54));
  AND2_X1   g797(.A1(KEYINPUT58), .A2(G475), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n974), .A2(G902), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n562), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n966), .A2(new_n562), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n987), .A2(new_n965), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT120), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT120), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n987), .A2(new_n991), .A3(new_n965), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(G60));
  INV_X1    g807(.A(KEYINPUT122), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n791), .B(KEYINPUT121), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n654), .B(KEYINPUT59), .Z(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n953), .A2(new_n931), .A3(new_n929), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n927), .A2(new_n928), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT53), .B1(new_n919), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT54), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n998), .B1(new_n1002), .B2(new_n955), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n994), .B1(new_n1003), .B2(new_n964), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n997), .B1(new_n978), .B2(new_n979), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(KEYINPUT122), .A3(new_n965), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n995), .B1(new_n956), .B2(new_n996), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(G63));
  INV_X1    g822(.A(KEYINPUT61), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G217), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT60), .Z(new_n1011));
  NAND2_X1  g825(.A1(new_n974), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n248), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n965), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1012), .A2(new_n676), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n964), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1018), .B(KEYINPUT61), .C1(new_n676), .C2(new_n1012), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(G66));
  NAND3_X1  g834(.A1(new_n621), .A2(G224), .A3(G953), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1021), .B1(new_n951), .B2(G953), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n968), .B1(G898), .B2(new_n191), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT123), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1022), .B(new_n1024), .ZN(G69));
  NAND3_X1  g839(.A1(new_n748), .A2(new_n738), .A3(new_n768), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n813), .B2(new_n818), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n843), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n760), .A2(new_n921), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1028), .A2(new_n857), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT125), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1031), .B1(new_n936), .B2(new_n786), .ZN(new_n1032));
  AND4_X1   g846(.A1(new_n1031), .A2(new_n773), .A3(new_n786), .A4(new_n775), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(KEYINPUT126), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n773), .A2(new_n786), .A3(new_n775), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1036), .B(KEYINPUT125), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1029), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n1027), .B2(new_n843), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT126), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .A4(new_n857), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1035), .A2(new_n1041), .A3(new_n191), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n343), .A2(new_n347), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(new_n545), .Z(new_n1044));
  AOI21_X1  g858(.A(new_n1044), .B1(G900), .B2(G953), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT124), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n388), .A2(new_n914), .A3(new_n702), .A4(new_n913), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1048), .A2(new_n808), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1029), .A2(KEYINPUT62), .A3(new_n712), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n712), .A2(new_n760), .A3(new_n921), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT62), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1049), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1054), .A2(new_n844), .A3(new_n857), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1055), .A2(new_n191), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1047), .B1(new_n1056), .B2(new_n1044), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1046), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1059), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1046), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1060), .A2(new_n1062), .ZN(G72));
  NAND2_X1  g877(.A1(G472), .A2(G902), .ZN(new_n1064));
  XOR2_X1   g878(.A(new_n1064), .B(KEYINPUT63), .Z(new_n1065));
  OAI21_X1  g879(.A(new_n1065), .B1(new_n1055), .B2(new_n951), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1066), .A2(new_n696), .ZN(new_n1067));
  INV_X1    g881(.A(new_n349), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n362), .A2(new_n368), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1068), .B1(new_n1069), .B2(KEYINPUT127), .ZN(new_n1070));
  OAI21_X1  g884(.A(new_n1070), .B1(KEYINPUT127), .B2(new_n1069), .ZN(new_n1071));
  NAND4_X1  g885(.A1(new_n932), .A2(new_n940), .A3(new_n1065), .A4(new_n1071), .ZN(new_n1072));
  NAND3_X1  g886(.A1(new_n1067), .A2(new_n965), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g887(.A1(new_n1035), .A2(new_n1041), .A3(new_n938), .ZN(new_n1074));
  NAND2_X1  g888(.A1(new_n1074), .A2(new_n1065), .ZN(new_n1075));
  NOR2_X1   g889(.A1(new_n358), .A2(new_n270), .ZN(new_n1076));
  AOI21_X1  g890(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(G57));
endmodule


