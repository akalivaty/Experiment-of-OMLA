//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT35), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT27), .B(G183gat), .Z(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G190gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT28), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT27), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT27), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n210), .A2(new_n206), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  OR3_X1    g013(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n207), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n211), .ZN(new_n228));
  NAND3_X1  g027(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n224), .B1(new_n219), .B2(new_n225), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n237), .A3(new_n216), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n223), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n225), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n240), .A2(new_n228), .A3(new_n229), .ZN(new_n241));
  NAND3_X1  g040(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n235), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n223), .B1(new_n216), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  OR3_X1    g045(.A1(new_n241), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n222), .B1(new_n239), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249));
  AND2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(KEYINPUT24), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n240), .A2(KEYINPUT64), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(new_n226), .ZN(new_n253));
  INV_X1    g052(.A(new_n238), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n241), .A2(new_n243), .A3(new_n246), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT66), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n221), .B1(new_n248), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G113gat), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n262));
  NAND2_X1  g061(.A1(G113gat), .A2(G120gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(KEYINPUT68), .A3(new_n266), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n258), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n207), .A2(new_n220), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n239), .A2(new_n222), .A3(new_n247), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT66), .B1(new_n255), .B2(new_n256), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n264), .A2(KEYINPUT68), .A3(new_n266), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n266), .B1(new_n264), .B2(KEYINPUT68), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n271), .A2(new_n273), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT32), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT33), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G15gat), .B(G43gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(G71gat), .ZN(new_n287));
  INV_X1    g086(.A(G99gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n282), .B(KEYINPUT32), .C1(new_n284), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n273), .B1(new_n271), .B2(new_n281), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT34), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n277), .A2(new_n280), .ZN(new_n297));
  AOI211_X1 g096(.A(new_n270), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n298));
  OAI211_X1 g097(.A(KEYINPUT34), .B(new_n272), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n290), .A2(new_n303), .A3(new_n292), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n294), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n301), .A2(new_n290), .A3(new_n303), .A4(new_n292), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n308));
  XOR2_X1   g107(.A(KEYINPUT71), .B(G218gat), .Z(new_n309));
  AOI21_X1  g108(.A(KEYINPUT22), .B1(new_n309), .B2(G211gat), .ZN(new_n310));
  XOR2_X1   g109(.A(G197gat), .B(G204gat), .Z(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(G211gat), .B(G218gat), .Z(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT72), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n312), .A2(new_n314), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n308), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n312), .A2(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n314), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT73), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322));
  INV_X1    g121(.A(G141gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(G148gat), .ZN(new_n324));
  INV_X1    g123(.A(G148gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(G141gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR3_X1   g128(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n322), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n332), .ZN(new_n337));
  OR2_X1    g136(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n325), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n323), .B2(G148gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n325), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n337), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n333), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n321), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n345), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n318), .B2(new_n319), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(KEYINPUT3), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(G228gat), .A3(G233gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n312), .A2(new_n313), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n348), .B1(new_n312), .B2(new_n313), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n346), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n351), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n350), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G78gat), .B(G106gat), .Z(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(G22gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT31), .B(G50gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n355), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n355), .B2(new_n361), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n307), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n333), .B(new_n345), .C1(new_n278), .C2(new_n279), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n270), .A2(KEYINPUT78), .A3(new_n345), .A4(new_n333), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n372), .B1(new_n376), .B2(KEYINPUT4), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n351), .A2(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(new_n280), .A3(new_n347), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n280), .A2(new_n351), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n374), .A2(new_n375), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n382), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n388), .B2(KEYINPUT5), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT5), .ZN(new_n390));
  AOI211_X1 g189(.A(KEYINPUT79), .B(new_n390), .C1(new_n387), .C2(new_n382), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n384), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n376), .A2(KEYINPUT4), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n370), .A2(new_n371), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n380), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n390), .A3(new_n381), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(G85gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT0), .B(G57gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n392), .A2(new_n396), .A3(new_n401), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n392), .B2(new_n396), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n407), .A2(KEYINPUT84), .A3(KEYINPUT6), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT84), .B1(new_n407), .B2(KEYINPUT6), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G8gat), .B(G36gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(KEYINPUT29), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n239), .A2(new_n247), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n221), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n277), .B2(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n317), .A2(new_n320), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n221), .A2(new_n417), .A3(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n277), .B2(new_n416), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n321), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n413), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n424), .A3(new_n413), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT30), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n421), .A2(new_n424), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n430));
  INV_X1    g229(.A(new_n413), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n203), .B1(new_n369), .B2(new_n434), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n295), .A2(KEYINPUT34), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT69), .A3(new_n299), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n293), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n301), .A2(new_n290), .A3(KEYINPUT69), .A4(new_n292), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n366), .A2(new_n367), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n407), .A2(KEYINPUT6), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n406), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n442), .A2(KEYINPUT35), .A3(new_n444), .A4(new_n433), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n368), .B1(new_n444), .B2(new_n433), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT36), .B1(new_n305), .B2(new_n306), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n438), .A2(KEYINPUT36), .A3(new_n439), .ZN(new_n449));
  NOR4_X1   g248(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT80), .A4(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT36), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n307), .B2(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n392), .A2(new_n396), .A3(new_n401), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n454), .A2(new_n407), .A3(KEYINPUT6), .ZN(new_n455));
  INV_X1    g254(.A(new_n443), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n433), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n441), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n451), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n450), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n429), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  MUX2_X1   g264(.A(new_n419), .B(new_n423), .S(new_n420), .Z(new_n466));
  AOI21_X1  g265(.A(KEYINPUT38), .B1(new_n466), .B2(KEYINPUT37), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n429), .A2(new_n462), .A3(new_n463), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n413), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n426), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n461), .B1(new_n410), .B2(new_n470), .ZN(new_n471));
  AOI211_X1 g270(.A(KEYINPUT83), .B(KEYINPUT37), .C1(new_n421), .C2(new_n424), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n464), .A2(new_n472), .A3(new_n431), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n425), .B1(new_n473), .B2(new_n467), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n443), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n407), .A2(KEYINPUT84), .A3(KEYINPUT6), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n474), .A2(new_n478), .A3(KEYINPUT85), .A4(new_n406), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT38), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n429), .A2(new_n463), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n473), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n393), .A2(new_n394), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n381), .B1(new_n487), .B2(new_n379), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n376), .A2(new_n381), .A3(new_n386), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT39), .B(new_n491), .C1(new_n395), .C2(new_n381), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n401), .B1(KEYINPUT81), .B2(KEYINPUT40), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT40), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n432), .A3(new_n428), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n403), .B1(new_n495), .B2(new_n499), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n501), .A2(KEYINPUT82), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT82), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n441), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n446), .B1(new_n460), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n509));
  OR3_X1    g308(.A1(new_n509), .A2(G29gat), .A3(G36gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(G29gat), .B2(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G50gat), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n515), .A2(G43gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(G43gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT15), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT86), .B(G43gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n515), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(KEYINPUT87), .A3(new_n516), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n522), .B2(KEYINPUT87), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n518), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n520), .B1(new_n527), .B2(new_n514), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  AND2_X1   g329(.A1(G15gat), .A2(G22gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(G15gat), .A2(G22gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n531), .B2(new_n532), .ZN(new_n535));
  INV_X1    g334(.A(G1gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI221_X1 g336(.A(new_n534), .B1(new_n530), .B2(G1gat), .C1(new_n531), .C2(new_n532), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT91), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT90), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(G8gat), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT93), .ZN(new_n544));
  INV_X1    g343(.A(G8gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(KEYINPUT90), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n544), .B1(new_n543), .B2(new_n546), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n529), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n539), .A2(KEYINPUT90), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n542), .A2(G8gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT93), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n547), .A3(new_n528), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(KEYINPUT94), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT13), .Z(new_n558));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n554), .A2(new_n559), .A3(new_n547), .A4(new_n528), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n556), .A2(KEYINPUT95), .A3(new_n558), .A4(new_n560), .ZN(new_n564));
  INV_X1    g363(.A(new_n520), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n521), .A2(new_n515), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT87), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT15), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n519), .B1(new_n568), .B2(new_n523), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT88), .B(new_n565), .C1(new_n569), .C2(new_n513), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n528), .A2(KEYINPUT88), .A3(KEYINPUT17), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n553), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n543), .A2(KEYINPUT92), .A3(new_n546), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n557), .A3(new_n555), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT18), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n578), .A2(new_n581), .A3(new_n557), .A4(new_n555), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n563), .A2(new_n564), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584));
  INV_X1    g383(.A(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT11), .B(G169gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT12), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT96), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n563), .A2(new_n564), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n580), .A2(new_n582), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n583), .A2(new_n596), .A3(new_n589), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n583), .B2(new_n589), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n590), .B(new_n595), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n202), .B1(new_n508), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n435), .A2(new_n445), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n290), .A2(new_n303), .A3(new_n292), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n303), .B1(new_n290), .B2(new_n292), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n603), .A2(new_n604), .A3(new_n301), .ZN(new_n605));
  INV_X1    g404(.A(new_n306), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n452), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n449), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n458), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT80), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n453), .A2(new_n451), .A3(new_n458), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n484), .B1(new_n471), .B2(new_n479), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT82), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n493), .B1(new_n488), .B2(new_n489), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n498), .B1(new_n615), .B2(new_n492), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n433), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n502), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n368), .B1(new_n619), .B2(new_n503), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n602), .B1(new_n612), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(KEYINPUT98), .A3(new_n599), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n601), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G57gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n628));
  INV_X1    g427(.A(G64gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G71gat), .ZN(new_n631));
  INV_X1    g430(.A(G78gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT9), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n632), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT9), .B1(new_n627), .B2(new_n629), .ZN(new_n638));
  NOR2_X1   g437(.A1(G57gat), .A2(G64gat), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n554), .A2(new_n547), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n209), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI211_X1 g446(.A(G183gat), .B(new_n645), .C1(new_n554), .C2(new_n547), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n548), .B2(new_n549), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(G183gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(new_n209), .A3(new_n646), .ZN(new_n652));
  INV_X1    g451(.A(new_n643), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G127gat), .B(G155gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G211gat), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n649), .A2(new_n654), .B1(G231gat), .B2(G233gat), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n655), .A2(new_n656), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n649), .A2(new_n654), .A3(G231gat), .A4(G233gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n626), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n659), .B1(new_n657), .B2(new_n660), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n662), .A3(new_n664), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n625), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G190gat), .B(G218gat), .ZN(new_n670));
  INV_X1    g469(.A(G134gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(G85gat), .A2(G92gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT101), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(G85gat), .A3(G92gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n675), .A3(KEYINPUT7), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n676), .B(new_n677), .C1(KEYINPUT7), .C2(new_n672), .ZN(new_n679));
  NAND2_X1  g478(.A1(G99gat), .A2(G106gat), .ZN(new_n680));
  INV_X1    g479(.A(G85gat), .ZN(new_n681));
  INV_X1    g480(.A(G92gat), .ZN(new_n682));
  AOI22_X1  g481(.A1(KEYINPUT8), .A2(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G99gat), .B(G106gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n678), .A2(new_n679), .A3(new_n685), .A4(new_n683), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(KEYINPUT103), .A3(new_n688), .ZN(new_n689));
  OR3_X1    g488(.A1(new_n684), .A2(KEYINPUT103), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n572), .B2(new_n573), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n528), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n671), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n691), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n574), .A2(new_n698), .ZN(new_n699));
  AND4_X1   g498(.A1(new_n671), .A2(new_n699), .A3(new_n696), .A4(new_n693), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n670), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT100), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G162gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(new_n696), .A3(new_n693), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G134gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n695), .A2(new_n671), .A3(new_n696), .ZN(new_n707));
  INV_X1    g506(.A(new_n670), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n701), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n704), .B1(new_n701), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n666), .A2(new_n669), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n666), .A2(new_n712), .A3(KEYINPUT104), .A4(new_n669), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(G120gat), .B(G148gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(G176gat), .B(G204gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(G230gat), .ZN(new_n722));
  INV_X1    g521(.A(G233gat), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT105), .B1(new_n691), .B2(new_n642), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n689), .A2(new_n690), .A3(new_n725), .A4(new_n641), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n642), .A2(new_n687), .A3(new_n688), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n722), .B(new_n723), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n728), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT10), .B(new_n731), .C1(new_n724), .C2(new_n726), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT10), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n698), .A2(new_n733), .A3(new_n641), .ZN(new_n734));
  OAI22_X1  g533(.A1(new_n732), .A2(new_n734), .B1(new_n722), .B2(new_n723), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n721), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n722), .A2(new_n723), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n727), .A2(new_n733), .A3(new_n728), .ZN(new_n738));
  INV_X1    g537(.A(new_n734), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n740), .A2(new_n729), .A3(new_n720), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n624), .A2(new_n717), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n444), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(new_n536), .ZN(G1324gat));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n433), .ZN(new_n746));
  NAND2_X1  g545(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n530), .A2(new_n545), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n746), .A2(KEYINPUT42), .A3(new_n747), .A4(new_n748), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n751), .B(new_n752), .C1(new_n545), .C2(new_n746), .ZN(G1325gat));
  INV_X1    g552(.A(new_n743), .ZN(new_n754));
  INV_X1    g553(.A(new_n453), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(G15gat), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(G15gat), .B1(new_n754), .B2(new_n307), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(G1326gat));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n368), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT43), .B(G22gat), .Z(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1327gat));
  OAI211_X1 g560(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n508), .C2(new_n712), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n763));
  INV_X1    g562(.A(new_n712), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n622), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n613), .B2(new_n620), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n712), .B1(new_n768), .B2(new_n602), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n769), .B2(new_n763), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n762), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n666), .A2(new_n669), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n742), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n773), .A2(new_n600), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G29gat), .B1(new_n776), .B2(new_n444), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n773), .A2(new_n774), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n601), .A2(new_n764), .A3(new_n623), .A4(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n779), .A2(G29gat), .A3(new_n444), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n777), .B1(new_n785), .B2(new_n786), .ZN(G1328gat));
  NOR3_X1   g586(.A1(new_n779), .A2(G36gat), .A3(new_n433), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT46), .ZN(new_n789));
  OAI21_X1  g588(.A(G36gat), .B1(new_n776), .B2(new_n433), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1329gat));
  OAI21_X1  g590(.A(new_n521), .B1(new_n776), .B2(new_n453), .ZN(new_n792));
  INV_X1    g591(.A(new_n779), .ZN(new_n793));
  INV_X1    g592(.A(new_n307), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n521), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n793), .A2(KEYINPUT108), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT108), .B1(new_n793), .B2(new_n795), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1330gat));
  NAND3_X1  g602(.A1(new_n771), .A2(new_n441), .A3(new_n775), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G50gat), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n368), .B1(new_n779), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n515), .B1(new_n779), .B2(new_n806), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n805), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT48), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n808), .B2(new_n809), .ZN(new_n816));
  INV_X1    g615(.A(new_n809), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT112), .A3(new_n807), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT48), .A4(new_n805), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n810), .A2(KEYINPUT111), .A3(new_n811), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n814), .A2(new_n819), .A3(new_n820), .ZN(G1331gat));
  AND2_X1   g620(.A1(new_n717), .A2(new_n600), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n742), .B1(new_n768), .B2(new_n602), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n444), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(new_n627), .ZN(G1332gat));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n433), .ZN(new_n827));
  NOR2_X1   g626(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n828));
  AND2_X1   g627(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n827), .B2(new_n828), .ZN(G1333gat));
  OAI21_X1  g630(.A(G71gat), .B1(new_n824), .B2(new_n453), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n307), .A2(new_n631), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g634(.A1(new_n824), .A2(new_n368), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(new_n632), .ZN(G1335gat));
  NOR2_X1   g636(.A1(new_n773), .A2(new_n599), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n769), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n769), .A2(KEYINPUT51), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n742), .A2(G85gat), .A3(new_n444), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT114), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847));
  INV_X1    g646(.A(new_n838), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT44), .B(new_n712), .C1(new_n768), .C2(new_n602), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n610), .B(new_n611), .C1(new_n613), .C2(new_n620), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n712), .B1(new_n850), .B2(new_n602), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n849), .A2(new_n766), .B1(new_n851), .B2(new_n763), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n848), .B1(new_n852), .B2(new_n762), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n847), .B1(new_n853), .B2(new_n774), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AND4_X1   g654(.A1(new_n847), .A2(new_n771), .A3(new_n774), .A4(new_n838), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n444), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n846), .B1(new_n858), .B2(new_n681), .ZN(G1336gat));
  NAND2_X1  g658(.A1(new_n853), .A2(new_n774), .ZN(new_n860));
  OAI21_X1  g659(.A(G92gat), .B1(new_n860), .B2(new_n433), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n742), .A2(G92gat), .A3(new_n433), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT115), .Z(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n841), .B2(new_n842), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT52), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n433), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n854), .B2(new_n856), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(KEYINPUT52), .A3(G92gat), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n864), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(G1337gat));
  NAND4_X1  g672(.A1(new_n843), .A2(new_n288), .A3(new_n774), .A4(new_n307), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n453), .B1(new_n855), .B2(new_n857), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n288), .ZN(G1338gat));
  NAND2_X1  g675(.A1(new_n843), .A2(new_n774), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(G106gat), .A3(new_n368), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(KEYINPUT53), .ZN(new_n879));
  OAI21_X1  g678(.A(G106gat), .B1(new_n860), .B2(new_n368), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n441), .B1(new_n854), .B2(new_n856), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n882), .B2(G106gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(G1339gat));
  AND4_X1   g684(.A1(new_n715), .A2(new_n716), .A3(new_n742), .A4(new_n600), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n558), .B1(new_n556), .B2(new_n560), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n557), .B1(new_n578), .B2(new_n555), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n588), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n583), .A2(new_n589), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT97), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n583), .A2(new_n596), .A3(new_n589), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n721), .B1(new_n740), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n738), .A2(new_n737), .A3(new_n739), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n735), .A2(KEYINPUT54), .A3(new_n898), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n897), .A2(new_n899), .A3(KEYINPUT55), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT55), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n900), .A2(new_n901), .A3(new_n741), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n895), .A2(new_n902), .A3(new_n764), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n599), .A2(new_n902), .B1(new_n895), .B2(new_n774), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n764), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n886), .B1(new_n772), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n369), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n444), .A2(new_n868), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n259), .A3(new_n600), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n599), .A2(new_n902), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n774), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n764), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n903), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n772), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n715), .A2(new_n716), .A3(new_n742), .A4(new_n600), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n444), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n917), .A2(new_n433), .A3(new_n442), .ZN(new_n918));
  AOI21_X1  g717(.A(G113gat), .B1(new_n918), .B2(new_n599), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n910), .A2(new_n919), .ZN(G1340gat));
  OAI21_X1  g719(.A(G120gat), .B1(new_n909), .B2(new_n742), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n260), .A3(new_n774), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT118), .Z(G1341gat));
  OAI21_X1  g723(.A(G127gat), .B1(new_n909), .B2(new_n772), .ZN(new_n925));
  INV_X1    g724(.A(G127gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n918), .A2(new_n926), .A3(new_n773), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1342gat));
  NAND3_X1  g727(.A1(new_n918), .A2(new_n671), .A3(new_n764), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT56), .Z(new_n930));
  OAI21_X1  g729(.A(G134gat), .B1(new_n909), .B2(new_n712), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1343gat));
  NOR2_X1   g731(.A1(new_n755), .A2(new_n368), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT121), .Z(new_n934));
  NAND4_X1  g733(.A1(new_n917), .A2(new_n323), .A3(new_n433), .A4(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n600), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n906), .B2(new_n368), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n915), .A2(new_n916), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(KEYINPUT57), .A3(new_n441), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(KEYINPUT119), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n453), .A2(new_n908), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI211_X1 g742(.A(new_n937), .B(new_n368), .C1(new_n915), .C2(new_n916), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT119), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n941), .A2(new_n599), .A3(new_n943), .A4(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n338), .A2(new_n339), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n936), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT58), .B1(new_n936), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n953), .B(KEYINPUT58), .C1(new_n936), .C2(new_n950), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n949), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n947), .A2(new_n948), .ZN(new_n956));
  INV_X1    g755(.A(new_n936), .ZN(new_n957));
  AOI22_X1  g756(.A1(new_n952), .A2(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n955), .A2(new_n958), .ZN(G1344gat));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT57), .B1(new_n939), .B2(new_n441), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n774), .B(new_n943), .C1(new_n961), .C2(new_n944), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G148gat), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n941), .A2(new_n774), .A3(new_n943), .A4(new_n946), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n325), .A2(KEYINPUT59), .ZN(new_n965));
  AOI22_X1  g764(.A1(KEYINPUT59), .A2(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n917), .A2(new_n433), .ZN(new_n967));
  INV_X1    g766(.A(new_n934), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n969), .A2(new_n325), .A3(new_n774), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n960), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n964), .A2(new_n965), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT59), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n962), .B2(G148gat), .ZN(new_n975));
  OAI211_X1 g774(.A(KEYINPUT123), .B(new_n970), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n972), .A2(new_n976), .ZN(G1345gat));
  AOI21_X1  g776(.A(G155gat), .B1(new_n969), .B2(new_n773), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n941), .A2(new_n943), .A3(new_n946), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n772), .A2(new_n334), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1346gat));
  AOI21_X1  g780(.A(G162gat), .B1(new_n969), .B2(new_n764), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n712), .A2(new_n335), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n979), .B2(new_n983), .ZN(G1347gat));
  NAND2_X1  g783(.A1(new_n444), .A2(new_n868), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n907), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(G169gat), .B1(new_n987), .B2(new_n600), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n939), .A2(new_n442), .A3(new_n986), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n990), .A2(new_n233), .A3(new_n599), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n988), .A2(new_n991), .ZN(G1348gat));
  OAI21_X1  g791(.A(G176gat), .B1(new_n987), .B2(new_n742), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n774), .A2(new_n234), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT124), .ZN(G1349gat));
  OAI21_X1  g795(.A(G183gat), .B1(new_n987), .B2(new_n772), .ZN(new_n997));
  OR3_X1    g796(.A1(new_n989), .A2(new_n772), .A3(new_n204), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT60), .ZN(new_n999));
  AOI22_X1  g798(.A1(new_n997), .A2(new_n998), .B1(KEYINPUT125), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n999), .A2(KEYINPUT125), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1000), .B(new_n1001), .ZN(G1350gat));
  OAI21_X1  g801(.A(G190gat), .B1(new_n987), .B2(new_n712), .ZN(new_n1003));
  XNOR2_X1  g802(.A(new_n1003), .B(KEYINPUT61), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n990), .A2(new_n211), .A3(new_n764), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1351gat));
  NAND2_X1  g805(.A1(new_n938), .A2(new_n940), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n755), .A2(new_n985), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT126), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n1007), .A2(G197gat), .A3(new_n599), .A4(new_n1009), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n939), .A2(new_n441), .A3(new_n1008), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n1011), .A2(new_n599), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1010), .B1(G197gat), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT127), .ZN(G1352gat));
  INV_X1    g813(.A(G204gat), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1011), .A2(new_n1015), .A3(new_n774), .ZN(new_n1016));
  XOR2_X1   g815(.A(new_n1016), .B(KEYINPUT62), .Z(new_n1017));
  AND3_X1   g816(.A1(new_n1007), .A2(new_n774), .A3(new_n1009), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1017), .B1(new_n1015), .B2(new_n1018), .ZN(G1353gat));
  INV_X1    g818(.A(G211gat), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1011), .A2(new_n1020), .A3(new_n773), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1007), .A2(new_n773), .A3(new_n1008), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1022), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1023));
  AOI21_X1  g822(.A(KEYINPUT63), .B1(new_n1022), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(G1354gat));
  AOI21_X1  g824(.A(G218gat), .B1(new_n1011), .B2(new_n764), .ZN(new_n1026));
  AND3_X1   g825(.A1(new_n1007), .A2(new_n764), .A3(new_n309), .ZN(new_n1027));
  AOI21_X1  g826(.A(new_n1026), .B1(new_n1027), .B2(new_n1009), .ZN(G1355gat));
endmodule


