//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n192), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT66), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n199), .A3(G131), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT0), .B1(new_n206), .B2(G128), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT0), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n204), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n202), .B2(G143), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n204), .A2(KEYINPUT65), .A3(G146), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n208), .B1(new_n213), .B2(G128), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n207), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT69), .B1(new_n201), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n212), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(G128), .A3(new_n203), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT0), .A3(new_n216), .ZN(new_n221));
  INV_X1    g035(.A(new_n207), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n200), .A4(new_n198), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G116), .B(G119), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT2), .B(G113), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n193), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n189), .A2(G137), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n213), .A2(new_n236), .A3(G128), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n206), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n215), .B1(new_n240), .B2(KEYINPUT67), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n236), .B1(G143), .B2(new_n202), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n239), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n197), .B(new_n235), .C1(new_n238), .C2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n226), .A2(KEYINPUT28), .A3(new_n232), .A4(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n223), .A2(new_n200), .A3(new_n198), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n246), .ZN(new_n249));
  INV_X1    g063(.A(new_n232), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n249), .B2(new_n250), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n255), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n226), .A2(KEYINPUT30), .A3(new_n246), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT68), .B1(new_n249), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n268));
  AOI211_X1 g082(.A(new_n268), .B(new_n265), .C1(new_n248), .C2(new_n246), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n264), .B(new_n250), .C1(new_n267), .C2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n226), .A2(new_n246), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n232), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n260), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n270), .A2(KEYINPUT31), .A3(new_n272), .A4(new_n260), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n263), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(G472), .A2(G902), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n187), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n276), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n262), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT32), .B1(new_n282), .B2(new_n278), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n277), .A2(new_n284), .A3(new_n279), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n280), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(new_n278), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n187), .A3(KEYINPUT32), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n226), .A2(new_n246), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT72), .B1(new_n289), .B2(new_n250), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n272), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n271), .A2(KEYINPUT72), .A3(new_n232), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(KEYINPUT28), .A3(new_n292), .ZN(new_n293));
  AND4_X1   g107(.A1(KEYINPUT29), .A2(new_n293), .A3(new_n260), .A4(new_n253), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n260), .B1(new_n270), .B2(new_n272), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n254), .B2(new_n261), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G472), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n286), .A2(new_n288), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n302));
  INV_X1    g116(.A(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n215), .A2(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT24), .B(G110), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT75), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT23), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n305), .B(new_n311), .Z(new_n312));
  OAI211_X1 g126(.A(new_n312), .B(new_n304), .C1(new_n310), .C2(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n309), .B1(new_n313), .B2(G110), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(G125), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(G146), .B(new_n317), .C1(new_n321), .C2(new_n315), .ZN(new_n322));
  XNOR2_X1  g136(.A(G125), .B(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n202), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n314), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(KEYINPUT74), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n317), .B1(new_n321), .B2(new_n315), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n202), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n326), .B(new_n328), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n306), .A2(new_n307), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n313), .A2(G110), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT76), .B(KEYINPUT77), .Z(new_n334));
  INV_X1    g148(.A(G953), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(G221), .A3(G234), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G137), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n325), .A2(new_n332), .A3(new_n339), .ZN(new_n342));
  AOI21_X1  g156(.A(G902), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n302), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n342), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n339), .B1(new_n325), .B2(new_n332), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n295), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n349));
  INV_X1    g163(.A(G217), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(G234), .B2(new_n295), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n341), .A2(new_n342), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n351), .A2(G902), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G469), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G140), .ZN(new_n359));
  INV_X1    g173(.A(G227), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G953), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n359), .B(new_n361), .Z(new_n362));
  INV_X1    g176(.A(G104), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G107), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(G107), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT81), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n366), .A2(new_n368), .A3(KEYINPUT81), .A4(G104), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n364), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT80), .B(KEYINPUT3), .C1(new_n363), .C2(G107), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(G104), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT80), .B1(new_n374), .B2(KEYINPUT3), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G101), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT84), .B(KEYINPUT4), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n366), .A2(new_n368), .A3(G104), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n384), .A2(new_n369), .B1(new_n363), .B2(G107), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n365), .B2(new_n366), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n372), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n381), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n381), .A3(new_n388), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n390), .B(G101), .C1(new_n371), .C2(new_n376), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n390), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n377), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n389), .B2(new_n390), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT83), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n223), .B(new_n380), .C1(new_n396), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n219), .A2(new_n203), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n215), .B2(new_n242), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n237), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n374), .A2(new_n364), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G101), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n391), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n238), .A2(new_n245), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n391), .A2(new_n407), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n411), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n201), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n402), .A2(new_n201), .A3(new_n410), .A4(new_n413), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n362), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n411), .A2(new_n412), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n201), .B1(new_n420), .B2(new_n408), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT12), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n201), .B2(KEYINPUT85), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n421), .A2(new_n423), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n419), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n421), .A2(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n421), .A2(new_n423), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(KEYINPUT86), .A3(new_n428), .ZN(new_n429));
  AND4_X1   g243(.A1(new_n417), .A2(new_n362), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n358), .B(new_n295), .C1(new_n418), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(G469), .A2(G902), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n416), .A2(new_n417), .A3(new_n362), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n428), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n417), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n362), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n437), .A3(G469), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n431), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT9), .B(G234), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G221), .B1(new_n441), .B2(G902), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT79), .Z(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT17), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n204), .ZN(new_n451));
  NOR2_X1   g265(.A1(KEYINPUT90), .A2(G143), .ZN(new_n452));
  OAI211_X1 g266(.A(G214), .B(new_n256), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n256), .A2(G214), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n450), .B2(new_n204), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n453), .A2(new_n455), .A3(new_n196), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n196), .B1(new_n453), .B2(new_n455), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n455), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n460), .A2(KEYINPUT91), .A3(G131), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n449), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n326), .B(new_n328), .Z(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(G131), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(new_n449), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G113), .B(G122), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT93), .B(G104), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n460), .A2(KEYINPUT18), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n457), .A2(KEYINPUT18), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n453), .A2(new_n455), .A3(new_n196), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n321), .A2(G146), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n324), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n471), .B1(new_n467), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n295), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(KEYINPUT94), .B(new_n295), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(G475), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n321), .A2(KEYINPUT19), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT19), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n323), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT92), .B1(new_n489), .B2(new_n202), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT92), .A4(new_n202), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n322), .ZN(new_n492));
  NOR4_X1   g306(.A1(new_n459), .A2(new_n490), .A3(new_n461), .A4(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n477), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n470), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n478), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G475), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n295), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT20), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n496), .A2(new_n500), .A3(new_n497), .A4(new_n295), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G952), .ZN(new_n503));
  AOI211_X1 g317(.A(G953), .B(new_n503), .C1(G234), .C2(G237), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT21), .B(G898), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n295), .B(new_n335), .C1(G234), .C2(G237), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G478), .ZN(new_n510));
  NOR2_X1   g324(.A1(KEYINPUT98), .A2(KEYINPUT15), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(KEYINPUT98), .A2(KEYINPUT15), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  XOR2_X1   g329(.A(G116), .B(G122), .Z(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT95), .ZN(new_n517));
  XNOR2_X1  g331(.A(G116), .B(G122), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n520), .A3(new_n368), .ZN(new_n521));
  INV_X1    g335(.A(G116), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(KEYINPUT14), .A3(G122), .ZN(new_n523));
  OAI211_X1 g337(.A(G107), .B(new_n523), .C1(new_n516), .C2(KEYINPUT14), .ZN(new_n524));
  XNOR2_X1  g338(.A(G128), .B(G143), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n525), .A2(new_n189), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n189), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n521), .B(new_n524), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n520), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G107), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n521), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT97), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT96), .B(KEYINPUT13), .Z(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n525), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n215), .A2(G143), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n189), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n526), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n531), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n532), .B1(new_n531), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n528), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n441), .A2(new_n350), .A3(G953), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n528), .B(new_n542), .C1(new_n539), .C2(new_n540), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n515), .B1(new_n546), .B2(new_n295), .ZN(new_n547));
  AOI211_X1 g361(.A(G902), .B(new_n514), .C1(new_n544), .C2(new_n545), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n485), .A2(new_n502), .A3(new_n509), .A4(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(G110), .B(G122), .Z(new_n551));
  OAI21_X1  g365(.A(new_n395), .B1(new_n392), .B2(new_n394), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n398), .A2(KEYINPUT83), .A3(new_n400), .ZN(new_n553));
  AOI211_X1 g367(.A(new_n232), .B(new_n379), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT5), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n303), .A3(G116), .ZN(new_n556));
  OAI211_X1 g370(.A(G113), .B(new_n556), .C1(new_n228), .C2(new_n555), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n230), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n412), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n551), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n250), .B(new_n380), .C1(new_n396), .C2(new_n401), .ZN(new_n561));
  INV_X1    g375(.A(new_n559), .ZN(new_n562));
  INV_X1    g376(.A(new_n551), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(KEYINPUT6), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n223), .A2(G125), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(G125), .B2(new_n411), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n335), .A2(G224), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT6), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n570), .B(new_n551), .C1(new_n554), .C2(new_n559), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n568), .B1(KEYINPUT88), .B2(KEYINPUT7), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(KEYINPUT88), .B2(KEYINPUT7), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT89), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n567), .A2(KEYINPUT7), .A3(new_n568), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n551), .B(KEYINPUT8), .Z(new_n578));
  NAND2_X1  g392(.A1(new_n412), .A2(new_n558), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT87), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n578), .B1(new_n580), .B2(new_n559), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n576), .A2(new_n564), .A3(new_n577), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n572), .A2(new_n295), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G210), .B1(G237), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n572), .A2(new_n295), .A3(new_n584), .A4(new_n582), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n448), .B(new_n550), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n301), .A2(new_n357), .A3(new_n446), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  OAI21_X1  g404(.A(G472), .B1(new_n277), .B2(G902), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n287), .A2(new_n591), .A3(new_n357), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n445), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n448), .B1(new_n586), .B2(new_n587), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n485), .A2(new_n502), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n544), .B2(new_n545), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(KEYINPUT33), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n597), .B(new_n600), .C1(new_n544), .C2(new_n545), .ZN(new_n601));
  OAI211_X1 g415(.A(G478), .B(new_n295), .C1(new_n599), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n546), .A2(new_n295), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n510), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n593), .A2(new_n509), .A3(new_n594), .A4(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  NOR2_X1   g423(.A1(new_n595), .A2(new_n549), .ZN(new_n610));
  AND4_X1   g424(.A1(new_n509), .A2(new_n593), .A3(new_n594), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT35), .B(G107), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  NAND2_X1  g427(.A1(new_n287), .A2(new_n591), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n339), .A2(KEYINPUT36), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n333), .B(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n617), .B2(new_n354), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n333), .B1(KEYINPUT36), .B2(new_n339), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n616), .A2(new_n325), .A3(new_n332), .ZN(new_n620));
  AND4_X1   g434(.A1(new_n615), .A2(new_n619), .A3(new_n354), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(new_n352), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  AND4_X1   g438(.A1(new_n444), .A2(new_n588), .A3(new_n439), .A4(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G110), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(G12));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n504), .B1(new_n507), .B2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n595), .A2(new_n549), .A3(new_n630), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n448), .B(new_n623), .C1(new_n586), .C2(new_n587), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n301), .A2(new_n446), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G128), .ZN(G30));
  XNOR2_X1  g448(.A(new_n630), .B(KEYINPUT39), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n446), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT40), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n637), .A2(KEYINPUT40), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n291), .A2(new_n261), .A3(new_n292), .ZN(new_n640));
  INV_X1    g454(.A(new_n273), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n295), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(G472), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n286), .A2(new_n643), .A3(new_n288), .ZN(new_n644));
  INV_X1    g458(.A(new_n549), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n623), .A2(new_n645), .A3(new_n595), .A4(new_n447), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n586), .A2(new_n587), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT38), .B1(new_n586), .B2(new_n587), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n649), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n656), .B1(new_n649), .B2(new_n655), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n638), .B(new_n639), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NOR3_X1   g474(.A1(new_n596), .A2(new_n605), .A3(new_n630), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n301), .A2(new_n446), .A3(new_n632), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G146), .ZN(G48));
  OAI21_X1  g477(.A(new_n295), .B1(new_n418), .B2(new_n430), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G469), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n665), .A2(new_n444), .A3(new_n431), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n301), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n594), .A2(new_n509), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n668), .A2(new_n596), .A3(new_n605), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n669), .A3(new_n357), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT41), .B(G113), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G15));
  NOR3_X1   g486(.A1(new_n668), .A2(new_n549), .A3(new_n595), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n667), .A2(new_n673), .A3(new_n357), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  NAND2_X1  g489(.A1(new_n622), .A2(new_n352), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n667), .A2(new_n588), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  NAND2_X1  g492(.A1(new_n595), .A2(new_n645), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n275), .A2(new_n276), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n260), .B1(new_n293), .B2(new_n253), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n278), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT104), .B(G472), .Z(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n277), .B2(G902), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n356), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n666), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  NOR2_X1   g503(.A1(new_n686), .A2(new_n623), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(new_n594), .A3(new_n661), .A4(new_n666), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G125), .ZN(G27));
  OAI21_X1  g506(.A(KEYINPUT105), .B1(new_n283), .B2(new_n285), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n278), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n284), .B1(new_n277), .B2(new_n279), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n693), .A2(new_n300), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(KEYINPUT42), .A3(new_n357), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n630), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n606), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n586), .A2(new_n447), .A3(new_n587), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n700), .A2(KEYINPUT106), .A3(new_n446), .A4(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n704), .A2(new_n698), .A3(KEYINPUT42), .A4(new_n357), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n706), .B1(new_n707), .B2(new_n445), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n586), .A2(new_n447), .A3(new_n587), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n301), .A2(new_n357), .A3(new_n446), .A4(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n710), .B1(new_n712), .B2(new_n702), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT107), .B(G131), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G33));
  INV_X1    g530(.A(new_n712), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n631), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G134), .ZN(G36));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n605), .B2(new_n595), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n602), .A2(new_n604), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n596), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n614), .A3(new_n676), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n724), .A2(KEYINPUT44), .A3(new_n614), .A4(new_n676), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n711), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n433), .A2(new_n437), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n433), .A2(new_n437), .A3(KEYINPUT45), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(G469), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n432), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(KEYINPUT46), .A3(new_n432), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n431), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n444), .A3(new_n636), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT108), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n732), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT110), .B(G137), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G39));
  NOR4_X1   g561(.A1(new_n301), .A2(new_n357), .A3(new_n702), .A4(new_n703), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n741), .A2(new_n431), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT46), .B1(new_n737), .B2(new_n432), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n750), .B(new_n444), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n750), .B1(new_n742), .B2(new_n444), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G140), .ZN(G42));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n670), .A2(new_n674), .A3(new_n677), .A4(new_n688), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n446), .A2(new_n690), .A3(new_n711), .A4(new_n661), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n623), .A2(new_n595), .A3(new_n645), .A4(new_n630), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n301), .A2(new_n446), .A3(new_n711), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n631), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n763), .B(new_n765), .C1(new_n712), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n709), .B2(new_n713), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n589), .A2(new_n769), .A3(new_n607), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n769), .B1(new_n589), .B2(new_n607), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n611), .A2(new_n625), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT115), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n589), .A2(new_n607), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT114), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n589), .A2(new_n769), .A3(new_n607), .ZN(new_n777));
  AND4_X1   g591(.A1(KEYINPUT115), .A2(new_n776), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n762), .B(new_n768), .C1(new_n774), .C2(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n633), .A2(new_n691), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n448), .B(new_n679), .C1(new_n586), .C2(new_n587), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n676), .A2(KEYINPUT116), .A3(new_n630), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT116), .B1(new_n676), .B2(new_n630), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n783), .A2(new_n439), .A3(new_n444), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(new_n644), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n780), .A2(KEYINPUT117), .A3(new_n662), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n785), .A2(new_n633), .A3(new_n662), .A4(new_n691), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n760), .B1(new_n779), .B2(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n787), .B1(new_n786), .B2(new_n790), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n772), .A2(KEYINPUT115), .A3(new_n773), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n776), .A2(new_n773), .A3(new_n777), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n761), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n797), .A2(new_n802), .A3(KEYINPUT53), .A4(new_n768), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT54), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n795), .A2(new_n796), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n760), .B1(new_n806), .B2(new_n779), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n808));
  INV_X1    g622(.A(new_n793), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n802), .A3(KEYINPUT53), .A4(new_n768), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n687), .A2(new_n504), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n720), .A2(new_n723), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n665), .A2(new_n444), .A3(new_n431), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n652), .A2(new_n654), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n448), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n815), .A2(new_n817), .A3(KEYINPUT50), .A4(new_n448), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n711), .A2(KEYINPUT118), .A3(new_n666), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n703), .B2(new_n814), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n823), .A2(new_n504), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n644), .A2(new_n356), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n596), .A3(new_n605), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(new_n690), .A3(new_n724), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n665), .ZN(new_n836));
  INV_X1    g650(.A(new_n431), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n443), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n754), .B2(new_n755), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n812), .A2(new_n813), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n711), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n844), .A2(KEYINPUT51), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT120), .B(new_n822), .C1(new_n831), .C2(new_n832), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n835), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n826), .A2(new_n606), .A3(new_n827), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n503), .A2(G953), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT48), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT121), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(KEYINPUT121), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n823), .A2(new_n504), .A3(new_n825), .A4(new_n724), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n698), .A2(new_n357), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n849), .B(new_n855), .C1(new_n856), .C2(new_n851), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n844), .A2(new_n822), .A3(new_n830), .A4(new_n828), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  AOI211_X1 g673(.A(new_n848), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n843), .A2(new_n594), .A3(new_n666), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n847), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n805), .A2(new_n811), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT122), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n503), .A2(new_n335), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n805), .A2(new_n862), .A3(new_n866), .A4(new_n811), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT49), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n840), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n840), .A2(new_n869), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n596), .A2(new_n722), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n816), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n444), .A3(new_n447), .A4(new_n827), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT113), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n868), .A2(new_n875), .ZN(G75));
  NAND2_X1  g690(.A1(new_n807), .A2(new_n810), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n877), .A2(G210), .A3(G902), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n565), .A2(new_n571), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(new_n569), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT55), .Z(new_n881));
  NOR3_X1   g695(.A1(new_n878), .A2(KEYINPUT56), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n335), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n881), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n295), .B1(new_n807), .B2(new_n810), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(G210), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n882), .A2(new_n883), .A3(new_n888), .ZN(G51));
  NAND2_X1  g703(.A1(new_n432), .A2(KEYINPUT57), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n432), .A2(KEYINPUT57), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n808), .B1(new_n807), .B2(new_n810), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n890), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n418), .A2(new_n430), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n737), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n885), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n883), .B1(new_n896), .B2(new_n898), .ZN(G54));
  NAND3_X1  g713(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n478), .A3(new_n495), .ZN(new_n901));
  INV_X1    g715(.A(new_n883), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .A4(new_n496), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G60));
  OR2_X1    g718(.A1(new_n599), .A2(new_n601), .ZN(new_n905));
  NAND2_X1  g719(.A1(G478), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT59), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n905), .B(new_n908), .C1(new_n892), .C2(new_n893), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n805), .B2(new_n811), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n909), .B(new_n902), .C1(new_n910), .C2(new_n905), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(G63));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n350), .A2(new_n295), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n877), .A2(new_n617), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n902), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n353), .B1(new_n877), .B2(new_n916), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n913), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n919), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(KEYINPUT61), .A3(new_n902), .A4(new_n917), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(G66));
  INV_X1    g737(.A(G224), .ZN(new_n924));
  OAI21_X1  g738(.A(G953), .B1(new_n506), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n802), .B2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n879), .B1(G898), .B2(new_n335), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(G69));
  NAND3_X1  g742(.A1(new_n781), .A2(new_n698), .A3(new_n357), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n731), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n744), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n780), .A2(new_n662), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n758), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n931), .A2(new_n714), .A3(new_n718), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n335), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n264), .B1(new_n267), .B2(new_n269), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT124), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n489), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n629), .B2(G953), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n758), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n659), .A2(new_n932), .ZN(new_n942));
  XOR2_X1   g756(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n659), .B(new_n932), .C1(KEYINPUT125), .C2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n717), .B(new_n636), .C1(new_n606), .C2(new_n610), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n745), .A2(new_n944), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n335), .A3(new_n938), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n360), .B2(new_n629), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G72));
  NAND2_X1  g766(.A1(G472), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT63), .Z(new_n954));
  INV_X1    g768(.A(new_n802), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n270), .A2(new_n272), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n261), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n883), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n934), .B2(new_n955), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n261), .A3(new_n958), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n804), .B(new_n954), .C1(new_n641), .C2(new_n296), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n960), .A2(new_n962), .A3(KEYINPUT127), .A4(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G57));
endmodule


