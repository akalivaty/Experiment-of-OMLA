

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U319 ( .A(n442), .B(n441), .ZN(n494) );
  XNOR2_X1 U320 ( .A(n392), .B(n391), .ZN(n503) );
  INV_X1 U321 ( .A(KEYINPUT92), .ZN(n394) );
  XNOR2_X1 U322 ( .A(n394), .B(KEYINPUT25), .ZN(n395) );
  XNOR2_X1 U323 ( .A(n396), .B(n395), .ZN(n399) );
  NOR2_X1 U324 ( .A1(n514), .A2(n400), .ZN(n401) );
  XNOR2_X1 U325 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n382) );
  XNOR2_X1 U326 ( .A(n428), .B(KEYINPUT67), .ZN(n429) );
  XNOR2_X1 U327 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U328 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U329 ( .A(n438), .B(n437), .ZN(n439) );
  INV_X1 U330 ( .A(n560), .ZN(n562) );
  XNOR2_X1 U331 ( .A(n440), .B(n439), .ZN(n573) );
  XNOR2_X1 U332 ( .A(n466), .B(KEYINPUT119), .ZN(n560) );
  INV_X1 U333 ( .A(G36GAT), .ZN(n443) );
  XNOR2_X1 U334 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U335 ( .A(n443), .B(KEYINPUT102), .ZN(n444) );
  XNOR2_X1 U336 ( .A(n472), .B(n471), .ZN(G1349GAT) );
  XNOR2_X1 U337 ( .A(n445), .B(n444), .ZN(G1329GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT38), .B(KEYINPUT99), .Z(n442) );
  INV_X1 U339 ( .A(G218GAT), .ZN(n287) );
  NAND2_X1 U340 ( .A1(n287), .A2(G92GAT), .ZN(n290) );
  INV_X1 U341 ( .A(G92GAT), .ZN(n288) );
  NAND2_X1 U342 ( .A1(n288), .A2(G218GAT), .ZN(n289) );
  NAND2_X1 U343 ( .A1(n290), .A2(n289), .ZN(n292) );
  XNOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n383) );
  XOR2_X1 U346 ( .A(KEYINPUT72), .B(n383), .Z(n294) );
  NAND2_X1 U347 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n303) );
  XOR2_X1 U349 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n296) );
  XNOR2_X1 U350 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(G134GAT), .B(KEYINPUT73), .Z(n328) );
  XOR2_X1 U353 ( .A(n297), .B(n328), .Z(n301) );
  XOR2_X1 U354 ( .A(G29GAT), .B(G43GAT), .Z(n299) );
  XNOR2_X1 U355 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n417) );
  XOR2_X1 U357 ( .A(G50GAT), .B(G162GAT), .Z(n346) );
  XNOR2_X1 U358 ( .A(n417), .B(n346), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U361 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n305) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(G85GAT), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U364 ( .A(G99GAT), .B(n306), .Z(n433) );
  XOR2_X1 U365 ( .A(n307), .B(n433), .Z(n552) );
  XNOR2_X1 U366 ( .A(KEYINPUT74), .B(n552), .ZN(n561) );
  XNOR2_X1 U367 ( .A(KEYINPUT36), .B(n561), .ZN(n579) );
  XOR2_X1 U368 ( .A(G57GAT), .B(KEYINPUT13), .Z(n424) );
  XOR2_X1 U369 ( .A(G78GAT), .B(G211GAT), .Z(n309) );
  XNOR2_X1 U370 ( .A(G183GAT), .B(G155GAT), .ZN(n308) );
  XNOR2_X1 U371 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U372 ( .A(n424), .B(n310), .Z(n312) );
  NAND2_X1 U373 ( .A1(G231GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U375 ( .A(n313), .B(KEYINPUT77), .Z(n316) );
  XNOR2_X1 U376 ( .A(G22GAT), .B(G15GAT), .ZN(n314) );
  XNOR2_X1 U377 ( .A(n314), .B(G1GAT), .ZN(n416) );
  XNOR2_X1 U378 ( .A(n416), .B(KEYINPUT14), .ZN(n315) );
  XNOR2_X1 U379 ( .A(n316), .B(n315), .ZN(n324) );
  XOR2_X1 U380 ( .A(G64GAT), .B(G71GAT), .Z(n318) );
  XNOR2_X1 U381 ( .A(G8GAT), .B(G127GAT), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U383 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n320) );
  XNOR2_X1 U384 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U386 ( .A(n322), .B(n321), .Z(n323) );
  XOR2_X1 U387 ( .A(n324), .B(n323), .Z(n557) );
  INV_X1 U388 ( .A(n557), .ZN(n577) );
  XOR2_X1 U389 ( .A(G85GAT), .B(G148GAT), .Z(n326) );
  XNOR2_X1 U390 ( .A(G29GAT), .B(G162GAT), .ZN(n325) );
  XNOR2_X1 U391 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U392 ( .A(n328), .B(n327), .Z(n330) );
  NAND2_X1 U393 ( .A1(G225GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n344) );
  XOR2_X1 U395 ( .A(KEYINPUT1), .B(KEYINPUT87), .Z(n332) );
  XNOR2_X1 U396 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U398 ( .A(KEYINPUT4), .B(G57GAT), .Z(n334) );
  XNOR2_X1 U399 ( .A(G120GAT), .B(KEYINPUT6), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U401 ( .A(n336), .B(n335), .Z(n342) );
  XOR2_X1 U402 ( .A(G127GAT), .B(KEYINPUT78), .Z(n338) );
  XNOR2_X1 U403 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n367) );
  XOR2_X1 U405 ( .A(G155GAT), .B(KEYINPUT2), .Z(n340) );
  XNOR2_X1 U406 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n339) );
  XNOR2_X1 U407 ( .A(n340), .B(n339), .ZN(n357) );
  XNOR2_X1 U408 ( .A(n367), .B(n357), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U410 ( .A(n344), .B(n343), .ZN(n514) );
  XNOR2_X1 U411 ( .A(G78GAT), .B(G204GAT), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n345), .B(G148GAT), .ZN(n430) );
  XOR2_X1 U413 ( .A(n430), .B(n346), .Z(n348) );
  NAND2_X1 U414 ( .A1(G228GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n348), .B(n347), .ZN(n361) );
  XOR2_X1 U416 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n350) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n349) );
  XNOR2_X1 U418 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U419 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n352) );
  XNOR2_X1 U420 ( .A(G218GAT), .B(G106GAT), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U422 ( .A(n354), .B(n353), .Z(n359) );
  XOR2_X1 U423 ( .A(G211GAT), .B(KEYINPUT84), .Z(n356) );
  XNOR2_X1 U424 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n386) );
  XNOR2_X1 U426 ( .A(n357), .B(n386), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n463) );
  XOR2_X1 U429 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n363) );
  NAND2_X1 U430 ( .A1(G227GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U431 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U432 ( .A(n364), .B(KEYINPUT82), .Z(n369) );
  XOR2_X1 U433 ( .A(G183GAT), .B(KEYINPUT19), .Z(n366) );
  XNOR2_X1 U434 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n387) );
  XNOR2_X1 U436 ( .A(n387), .B(n367), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n380) );
  XOR2_X1 U438 ( .A(KEYINPUT81), .B(G176GAT), .Z(n371) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(KEYINPUT80), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n378) );
  XOR2_X1 U441 ( .A(KEYINPUT79), .B(G99GAT), .Z(n373) );
  XNOR2_X1 U442 ( .A(G15GAT), .B(G190GAT), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U444 ( .A(n374), .B(G134GAT), .Z(n376) );
  XOR2_X1 U445 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U446 ( .A(G43GAT), .B(n434), .ZN(n375) );
  XNOR2_X1 U447 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U448 ( .A(n378), .B(n377), .Z(n379) );
  XOR2_X1 U449 ( .A(n380), .B(n379), .Z(n518) );
  INV_X1 U450 ( .A(n518), .ZN(n525) );
  XOR2_X1 U451 ( .A(G169GAT), .B(G8GAT), .Z(n421) );
  XNOR2_X1 U452 ( .A(G204GAT), .B(KEYINPUT90), .ZN(n381) );
  XOR2_X1 U453 ( .A(G176GAT), .B(G64GAT), .Z(n425) );
  XNOR2_X1 U454 ( .A(n381), .B(n425), .ZN(n385) );
  XOR2_X1 U455 ( .A(n385), .B(n384), .Z(n389) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n421), .B(n390), .ZN(n392) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  NOR2_X1 U460 ( .A1(n525), .A2(n503), .ZN(n393) );
  NOR2_X1 U461 ( .A1(n463), .A2(n393), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n503), .B(KEYINPUT27), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n463), .A2(n525), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n397), .B(KEYINPUT26), .ZN(n566) );
  NOR2_X1 U465 ( .A1(n402), .A2(n566), .ZN(n398) );
  NOR2_X1 U466 ( .A1(n399), .A2(n398), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(KEYINPUT93), .ZN(n406) );
  XOR2_X1 U468 ( .A(KEYINPUT28), .B(n463), .Z(n507) );
  INV_X1 U469 ( .A(n507), .ZN(n526) );
  INV_X1 U470 ( .A(n514), .ZN(n499) );
  NOR2_X1 U471 ( .A1(n499), .A2(n402), .ZN(n403) );
  XOR2_X1 U472 ( .A(KEYINPUT91), .B(n403), .Z(n528) );
  NAND2_X1 U473 ( .A1(n528), .A2(n525), .ZN(n404) );
  OR2_X1 U474 ( .A1(n526), .A2(n404), .ZN(n405) );
  AND2_X1 U475 ( .A1(n406), .A2(n405), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n407), .B(KEYINPUT94), .ZN(n475) );
  NOR2_X1 U477 ( .A1(n577), .A2(n475), .ZN(n408) );
  NAND2_X1 U478 ( .A1(n579), .A2(n408), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n409), .B(KEYINPUT37), .ZN(n511) );
  XOR2_X1 U480 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n411) );
  XNOR2_X1 U481 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n410) );
  XNOR2_X1 U482 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U483 ( .A(G197GAT), .B(G141GAT), .Z(n413) );
  XNOR2_X1 U484 ( .A(G50GAT), .B(G36GAT), .ZN(n412) );
  XNOR2_X1 U485 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U486 ( .A(n415), .B(n414), .Z(n419) );
  XNOR2_X1 U487 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U488 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U489 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U490 ( .A1(G229GAT), .A2(G233GAT), .ZN(n422) );
  XOR2_X1 U491 ( .A(n423), .B(n422), .Z(n568) );
  INV_X1 U492 ( .A(n568), .ZN(n555) );
  XOR2_X1 U493 ( .A(KEYINPUT33), .B(n424), .Z(n427) );
  XNOR2_X1 U494 ( .A(n425), .B(G92GAT), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n432) );
  AND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n428) );
  XOR2_X1 U497 ( .A(n432), .B(n431), .Z(n440) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U499 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n436) );
  XNOR2_X1 U500 ( .A(KEYINPUT70), .B(KEYINPUT32), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  NOR2_X1 U502 ( .A1(n555), .A2(n573), .ZN(n477) );
  NAND2_X1 U503 ( .A1(n511), .A2(n477), .ZN(n441) );
  NOR2_X1 U504 ( .A1(n494), .A2(n503), .ZN(n445) );
  XNOR2_X1 U505 ( .A(KEYINPUT41), .B(n573), .ZN(n544) );
  INV_X1 U506 ( .A(n503), .ZN(n516) );
  NOR2_X1 U507 ( .A1(n555), .A2(n544), .ZN(n447) );
  XNOR2_X1 U508 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  NOR2_X1 U510 ( .A1(n448), .A2(n577), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n449), .B(KEYINPUT111), .ZN(n450) );
  NOR2_X1 U512 ( .A1(n552), .A2(n450), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n451), .B(KEYINPUT47), .ZN(n457) );
  XOR2_X1 U514 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n453) );
  NAND2_X1 U515 ( .A1(n577), .A2(n579), .ZN(n452) );
  XNOR2_X1 U516 ( .A(n453), .B(n452), .ZN(n454) );
  NOR2_X1 U517 ( .A1(n454), .A2(n573), .ZN(n455) );
  NAND2_X1 U518 ( .A1(n455), .A2(n555), .ZN(n456) );
  NAND2_X1 U519 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n458), .B(KEYINPUT48), .ZN(n527) );
  NAND2_X1 U521 ( .A1(n516), .A2(n527), .ZN(n461) );
  XNOR2_X1 U522 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n459) );
  XNOR2_X1 U523 ( .A(n459), .B(KEYINPUT54), .ZN(n460) );
  XNOR2_X1 U524 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U525 ( .A1(n462), .A2(n499), .ZN(n565) );
  NOR2_X1 U526 ( .A1(n463), .A2(n565), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n464), .B(KEYINPUT55), .ZN(n465) );
  NOR2_X1 U528 ( .A1(n525), .A2(n465), .ZN(n466) );
  NOR2_X1 U529 ( .A1(n544), .A2(n560), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n468) );
  XNOR2_X1 U531 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n467) );
  XNOR2_X1 U532 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U533 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n469) );
  NOR2_X1 U534 ( .A1(n561), .A2(n557), .ZN(n473) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U536 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U537 ( .A(KEYINPUT95), .B(n476), .Z(n498) );
  NAND2_X1 U538 ( .A1(n477), .A2(n498), .ZN(n486) );
  NOR2_X1 U539 ( .A1(n499), .A2(n486), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  NOR2_X1 U543 ( .A1(n503), .A2(n486), .ZN(n481) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n486), .A2(n525), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n483) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U548 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NOR2_X1 U550 ( .A1(n507), .A2(n486), .ZN(n487) );
  XOR2_X1 U551 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  NOR2_X1 U552 ( .A1(n499), .A2(n494), .ZN(n491) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n489) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U555 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n494), .A2(n525), .ZN(n492) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(n492), .Z(n493) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NOR2_X1 U560 ( .A1(n494), .A2(n507), .ZN(n496) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n496), .B(n495), .ZN(G1331GAT) );
  NOR2_X1 U563 ( .A1(n568), .A2(n544), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n497), .B(KEYINPUT104), .ZN(n512) );
  NAND2_X1 U565 ( .A1(n498), .A2(n512), .ZN(n506) );
  NOR2_X1 U566 ( .A1(n499), .A2(n506), .ZN(n501) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT105), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n503), .A2(n506), .ZN(n504) );
  XOR2_X1 U571 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U572 ( .A1(n525), .A2(n506), .ZN(n505) );
  XOR2_X1 U573 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U574 ( .A1(n507), .A2(n506), .ZN(n509) );
  XNOR2_X1 U575 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(KEYINPUT107), .ZN(n520) );
  NAND2_X1 U580 ( .A1(n520), .A2(n514), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n520), .A2(n516), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n524) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n522) );
  NAND2_X1 U588 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(G1339GAT) );
  OR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n530) );
  NAND2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U593 ( .A(KEYINPUT112), .B(n529), .ZN(n542) );
  NOR2_X1 U594 ( .A1(n530), .A2(n542), .ZN(n539) );
  INV_X1 U595 ( .A(n539), .ZN(n536) );
  NOR2_X1 U596 ( .A1(n555), .A2(n536), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1340GAT) );
  NOR2_X1 U599 ( .A1(n544), .A2(n536), .ZN(n534) );
  XNOR2_X1 U600 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G120GAT), .B(n535), .ZN(G1341GAT) );
  NOR2_X1 U603 ( .A1(n557), .A2(n536), .ZN(n537) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(n537), .Z(n538) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U607 ( .A1(n539), .A2(n561), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U609 ( .A1(n566), .A2(n542), .ZN(n551) );
  INV_X1 U610 ( .A(n551), .ZN(n549) );
  NOR2_X1 U611 ( .A1(n555), .A2(n549), .ZN(n543) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n549), .A2(n544), .ZN(n548) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT115), .ZN(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n557), .A2(n549), .ZN(n550) );
  XOR2_X1 U619 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n553), .B(KEYINPUT116), .ZN(n554) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n560), .ZN(n556) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n556), .Z(G1348GAT) );
  NOR2_X1 U625 ( .A1(n557), .A2(n560), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1350GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT58), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT124), .B(n567), .ZN(n580) );
  AND2_X1 U633 ( .A1(n580), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n580), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n582) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

