//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0007(.A1(G97), .A2(G107), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT65), .Z(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n216), .A2(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G58), .B2(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n222), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(G87), .B2(G250), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT66), .B(G244), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G77), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n221), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G238), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n203), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n215), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT1), .Z(new_n234));
  NOR2_X1   g0034(.A1(new_n215), .A2(G13), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G250), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(new_n223), .B2(new_n225), .ZN(new_n237));
  NAND2_X1  g0037(.A1(G1), .A2(G13), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n238), .A2(new_n213), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n204), .A2(new_n205), .ZN(new_n240));
  NOR2_X1   g0040(.A1(new_n240), .A2(new_n216), .ZN(new_n241));
  AOI22_X1  g0041(.A1(new_n237), .A2(KEYINPUT0), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  OAI211_X1 g0042(.A(new_n234), .B(new_n242), .C1(KEYINPUT0), .C2(new_n237), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(G361));
  XOR2_X1   g0044(.A(G238), .B(G244), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT2), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n217), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G250), .B(G257), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G264), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n219), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G358));
  XNOR2_X1  g0052(.A(G50), .B(G68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G87), .B(G97), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(G107), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(new_n218), .ZN(new_n258));
  XOR2_X1   g0058(.A(new_n255), .B(new_n258), .Z(G351));
  OAI21_X1  g0059(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G150), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT69), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n213), .A2(KEYINPUT69), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT8), .B(G58), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n260), .B(new_n262), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n238), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n270), .A2(new_n272), .B1(new_n216), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n272), .B1(new_n212), .B2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n275), .B1(new_n216), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT9), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G222), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G77), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n282), .B1(new_n283), .B2(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n238), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT67), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n287), .B2(new_n238), .ZN(new_n292));
  AND2_X1   g0092(.A1(G1), .A2(G13), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(KEYINPUT67), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n290), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G41), .ZN(new_n297));
  INV_X1    g0097(.A(G45), .ZN(new_n298));
  AOI21_X1  g0098(.A(G1), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n292), .B2(new_n295), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT68), .B(G226), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n289), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(G200), .B2(new_n304), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n279), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT10), .B1(new_n307), .B2(KEYINPUT70), .ZN(new_n309));
  XOR2_X1   g0109(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n278), .B(new_n312), .C1(G179), .C2(new_n304), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT7), .B1(new_n317), .B2(new_n213), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT7), .ZN(new_n319));
  NOR4_X1   g0119(.A1(new_n315), .A2(new_n316), .A3(new_n319), .A4(G20), .ZN(new_n320));
  OAI21_X1  g0120(.A(G68), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n261), .A2(G159), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n202), .A2(new_n203), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n240), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT16), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n321), .A2(KEYINPUT16), .A3(new_n322), .A4(new_n324), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n272), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT77), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n327), .A2(KEYINPUT77), .A3(new_n272), .A4(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n269), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n274), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n277), .B2(new_n334), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n301), .A2(G232), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n280), .A2(G223), .A3(new_n281), .ZN(new_n341));
  INV_X1    g0141(.A(G87), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n341), .B1(new_n264), .B2(new_n342), .C1(new_n284), .C2(new_n217), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n288), .B1(new_n299), .B2(new_n296), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G200), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n340), .A2(G190), .A3(new_n344), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n333), .A2(new_n337), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT17), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n336), .B1(new_n331), .B2(new_n332), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT17), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n346), .A4(new_n347), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n333), .A2(new_n337), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n311), .B1(new_n340), .B2(new_n344), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n355), .B1(new_n356), .B2(new_n345), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(KEYINPUT18), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n345), .A2(new_n356), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n354), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n350), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n349), .A2(new_n352), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n231), .B1(new_n301), .B2(KEYINPUT73), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(KEYINPUT73), .B2(new_n301), .ZN(new_n365));
  OAI211_X1 g0165(.A(G232), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT71), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n280), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n280), .A2(G226), .A3(new_n281), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G97), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n372), .A2(KEYINPUT72), .A3(new_n288), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT72), .B1(new_n372), .B2(new_n288), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n300), .B(new_n365), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n305), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n267), .A2(G77), .B1(G50), .B2(new_n261), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n213), .B2(G68), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n272), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT11), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT11), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n384), .A3(new_n272), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n383), .A2(new_n385), .B1(G68), .B2(new_n276), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n274), .A2(KEYINPUT74), .A3(new_n203), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT12), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT74), .B1(new_n274), .B2(new_n203), .ZN(new_n389));
  XOR2_X1   g0189(.A(new_n388), .B(new_n389), .Z(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G200), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n376), .B2(new_n377), .ZN(new_n395));
  OR3_X1    g0195(.A1(new_n379), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n314), .A2(new_n363), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n398), .B(G169), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n378), .A2(new_n398), .A3(new_n403), .A4(G169), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n376), .A2(G179), .A3(new_n377), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n393), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n317), .B1(G232), .B2(new_n281), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n231), .B2(new_n281), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n409), .B(new_n288), .C1(G107), .C2(new_n280), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n301), .A2(new_n228), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n300), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n311), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n334), .A2(new_n261), .ZN(new_n414));
  XOR2_X1   g0214(.A(KEYINPUT15), .B(G87), .Z(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n414), .B1(new_n213), .B2(new_n283), .C1(new_n268), .C2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n272), .B1(new_n283), .B2(new_n274), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n283), .B2(new_n277), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n413), .B(new_n419), .C1(G179), .C2(new_n412), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n407), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(G200), .B2(new_n412), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n305), .B2(new_n412), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n397), .A2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n213), .A2(KEYINPUT23), .A3(G107), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT23), .B1(new_n213), .B2(G107), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT86), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n213), .C2(G107), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n213), .A2(G33), .A3(G116), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n213), .B(G87), .C1(new_n315), .C2(new_n316), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT22), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n280), .A2(KEYINPUT22), .A3(new_n213), .A4(G87), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n431), .A2(new_n432), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n437), .A2(KEYINPUT24), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(KEYINPUT24), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n272), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT87), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT87), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(new_n272), .C1(new_n438), .C2(new_n439), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT25), .B1(new_n274), .B2(new_n224), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n274), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n212), .A2(G33), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n273), .A2(new_n448), .A3(new_n238), .A4(new_n271), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n446), .A2(new_n447), .B1(G107), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n280), .A2(G250), .A3(new_n281), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n284), .B2(new_n223), .ZN(new_n454));
  INV_X1    g0254(.A(G294), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n264), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n288), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n212), .A2(G45), .ZN(new_n458));
  OR2_X1    g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  NAND2_X1  g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n287), .A2(new_n291), .A3(new_n238), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT67), .B1(new_n293), .B2(new_n294), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n461), .B(G274), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n298), .A2(G1), .ZN(new_n465));
  INV_X1    g0265(.A(new_n460), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G264), .B(new_n468), .C1(new_n462), .C2(new_n463), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n457), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G169), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT88), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n457), .A2(new_n469), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(G179), .A3(new_n464), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n470), .A2(KEYINPUT88), .A3(new_n356), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n452), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G244), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT82), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n280), .A2(new_n483), .A3(G244), .A4(G1698), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G116), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n280), .A2(G238), .A3(new_n281), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n482), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n288), .ZN(new_n488));
  OAI211_X1 g0288(.A(G250), .B(new_n458), .C1(new_n462), .C2(new_n463), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n465), .A2(new_n291), .A3(G274), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n356), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n415), .A2(new_n273), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n280), .A2(new_n213), .A3(G68), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT19), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n213), .B1(new_n371), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G87), .B2(new_n209), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n222), .B1(new_n265), .B2(new_n266), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n494), .B(new_n497), .C1(new_n498), .C2(KEYINPUT19), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n493), .B1(new_n499), .B2(new_n272), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n450), .A2(new_n415), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n489), .A2(new_n490), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(new_n288), .B2(new_n487), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n492), .B(new_n502), .C1(new_n504), .C2(G169), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n488), .A2(G190), .A3(new_n491), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n449), .A2(new_n342), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n493), .B(new_n507), .C1(new_n499), .C2(new_n272), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n506), .B(new_n508), .C1(new_n504), .C2(new_n394), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n505), .A2(new_n509), .A3(KEYINPUT83), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT83), .B1(new_n505), .B2(new_n509), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G257), .B(new_n281), .C1(new_n315), .C2(new_n316), .ZN(new_n513));
  OAI211_X1 g0313(.A(G264), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n514));
  INV_X1    g0314(.A(G303), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n280), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(new_n288), .B1(new_n296), .B2(new_n461), .ZN(new_n517));
  OAI211_X1 g0317(.A(G270), .B(new_n468), .C1(new_n462), .C2(new_n463), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(KEYINPUT21), .A3(G169), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n288), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n521), .A2(G179), .A3(new_n464), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n274), .A2(new_n218), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G283), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n525), .B(new_n213), .C1(G33), .C2(new_n222), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n272), .C1(new_n213), .C2(G116), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT20), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  OAI221_X1 g0330(.A(new_n524), .B1(new_n218), .B2(new_n449), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G169), .A3(new_n519), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT84), .B(KEYINPUT21), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n523), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n480), .A2(new_n512), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n470), .A2(G200), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n474), .A2(G190), .A3(new_n464), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n444), .A2(new_n451), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(G257), .B(new_n468), .C1(new_n462), .C2(new_n463), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n464), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT80), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT80), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n464), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(new_n281), .C1(new_n315), .C2(new_n316), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n525), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n288), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT81), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n464), .A2(new_n539), .A3(new_n542), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n542), .B1(new_n464), .B2(new_n539), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n551), .B(KEYINPUT81), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G190), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(G107), .B1(new_n318), .B2(new_n320), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n222), .A2(new_n224), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n208), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n563), .B2(KEYINPUT6), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G20), .ZN(new_n565));
  OAI211_X1 g0365(.A(KEYINPUT79), .B(G107), .C1(new_n318), .C2(new_n320), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n261), .A2(G77), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n560), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n272), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n274), .A2(new_n222), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n449), .B2(new_n222), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G200), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n557), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n541), .A2(new_n543), .B1(new_n288), .B2(new_n550), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n569), .A2(new_n572), .B1(new_n578), .B2(new_n356), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT81), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n311), .A3(new_n555), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n531), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n517), .A2(G190), .A3(new_n518), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n519), .A2(G200), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT85), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n584), .A2(new_n586), .A3(new_n589), .A4(new_n585), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n538), .A2(new_n577), .A3(new_n583), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n535), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n425), .A2(new_n593), .ZN(G372));
  NAND2_X1  g0394(.A1(new_n349), .A2(new_n352), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n379), .A2(new_n393), .A3(new_n395), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n421), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n358), .A2(new_n362), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n310), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n601), .A2(new_n313), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n505), .A2(new_n509), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT26), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n582), .A4(new_n579), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n605), .A2(new_n505), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n505), .A2(new_n509), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT83), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n505), .A2(new_n509), .A3(KEYINPUT83), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n582), .A4(new_n579), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT26), .ZN(new_n612));
  INV_X1    g0412(.A(new_n451), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n441), .B2(new_n443), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n477), .B1(new_n473), .B2(new_n475), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n534), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n603), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n538), .A2(new_n577), .A3(new_n583), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n606), .B(new_n612), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n425), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n602), .A2(new_n620), .ZN(G369));
  INV_X1    g0421(.A(G13), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(G20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n212), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G213), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n480), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n629), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n538), .B1(new_n614), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n630), .B1(new_n480), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G330), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n591), .B(new_n534), .C1(new_n584), .C2(new_n631), .ZN(new_n635));
  OR3_X1    g0435(.A1(new_n534), .A2(new_n584), .A3(new_n631), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n480), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n534), .A2(new_n629), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n630), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(new_n641), .ZN(G399));
  INV_X1    g0442(.A(new_n235), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G41), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n208), .A2(new_n342), .A3(new_n218), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT89), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(G1), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n241), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n645), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT28), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n611), .A2(KEYINPUT26), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT26), .B1(new_n583), .B2(new_n607), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n505), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT94), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n581), .A2(new_n555), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n573), .B1(new_n656), .B2(G190), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n576), .B1(new_n582), .B2(new_n579), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n658), .A2(new_n603), .A3(new_n616), .A4(new_n538), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT94), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n652), .A2(new_n660), .A3(new_n505), .A4(new_n653), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n655), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(KEYINPUT29), .A3(new_n631), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n605), .A2(new_n505), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(KEYINPUT26), .B2(new_n611), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n629), .B1(new_n665), .B2(new_n659), .ZN(new_n666));
  XNOR2_X1  g0466(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n522), .A2(KEYINPUT90), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n517), .A2(new_n670), .A3(G179), .A4(new_n518), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n669), .A2(new_n474), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n656), .A2(new_n672), .A3(new_n504), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n504), .ZN(new_n676));
  AOI21_X1  g0476(.A(G179), .B1(new_n517), .B2(new_n518), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n575), .A3(new_n470), .A4(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n656), .A2(new_n672), .A3(KEYINPUT30), .A4(new_n504), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT31), .B1(new_n680), .B2(new_n629), .ZN(new_n683));
  OR3_X1    g0483(.A1(new_n682), .A2(KEYINPUT91), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT91), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT92), .B1(new_n593), .B2(new_n631), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT92), .ZN(new_n687));
  NOR4_X1   g0487(.A1(new_n535), .A2(new_n592), .A3(new_n687), .A4(new_n629), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n684), .B(new_n685), .C1(new_n686), .C2(new_n688), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n663), .A2(new_n668), .B1(new_n689), .B2(G330), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n651), .B1(new_n690), .B2(G1), .ZN(G364));
  AOI21_X1  g0491(.A(new_n238), .B1(G20), .B2(new_n311), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n213), .A2(new_n356), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n305), .A3(G200), .ZN(new_n694));
  XOR2_X1   g0494(.A(KEYINPUT33), .B(G317), .Z(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n213), .A2(G190), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n394), .A2(G179), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n356), .A2(G200), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n697), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(G283), .A2(new_n700), .B1(new_n703), .B2(G311), .ZN(new_n704));
  NOR2_X1   g0504(.A1(G179), .A2(G200), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G329), .ZN(new_n708));
  INV_X1    g0508(.A(G322), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n213), .A2(new_n305), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n701), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n704), .B(new_n708), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n693), .A2(G190), .A3(G200), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI211_X1 g0514(.A(new_n696), .B(new_n712), .C1(G326), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n710), .A2(new_n698), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n317), .B1(new_n716), .B2(new_n515), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT99), .Z(new_n718));
  AOI21_X1  g0518(.A(new_n213), .B1(new_n705), .B2(G190), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n715), .B(new_n718), .C1(new_n455), .C2(new_n719), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT100), .Z(new_n721));
  OR2_X1    g0521(.A1(new_n703), .A2(KEYINPUT98), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n703), .A2(KEYINPUT98), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G77), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n280), .B1(new_n716), .B2(new_n342), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n694), .A2(new_n203), .B1(new_n713), .B2(new_n216), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n727), .B(new_n728), .C1(G107), .C2(new_n700), .ZN(new_n729));
  INV_X1    g0529(.A(G159), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n706), .A2(KEYINPUT32), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT32), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n707), .B2(G159), .ZN(new_n733));
  INV_X1    g0533(.A(new_n719), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n731), .B(new_n733), .C1(G97), .C2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n726), .A2(new_n729), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n711), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(G58), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n692), .B1(new_n721), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n622), .A2(new_n264), .A3(KEYINPUT97), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT97), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(G13), .B2(G33), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n692), .ZN(new_n746));
  XNOR2_X1  g0546(.A(G355), .B(KEYINPUT95), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n643), .A2(new_n317), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n747), .A2(new_n748), .B1(new_n218), .B2(new_n643), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT96), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n643), .A2(new_n280), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n649), .A2(G45), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n752), .B(new_n753), .C1(new_n255), .C2(G45), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n746), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n635), .A2(new_n636), .ZN(new_n756));
  INV_X1    g0556(.A(new_n745), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n739), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n212), .B1(new_n623), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n644), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n761), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n756), .A2(G330), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n637), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT101), .Z(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(G396));
  NAND2_X1  g0568(.A1(new_n689), .A2(G330), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n420), .A2(new_n629), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n419), .A2(new_n629), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT104), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n423), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(new_n773), .B2(new_n420), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n619), .A2(new_n631), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT105), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT105), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n619), .A2(new_n777), .A3(new_n631), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n666), .B2(new_n774), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n769), .B(new_n780), .Z(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n763), .ZN(new_n782));
  INV_X1    g0582(.A(new_n694), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n783), .A2(G150), .B1(new_n714), .B2(G137), .ZN(new_n784));
  INV_X1    g0584(.A(G143), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n784), .B1(new_n785), .B2(new_n711), .C1(new_n724), .C2(new_n730), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT34), .ZN(new_n787));
  INV_X1    g0587(.A(new_n716), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G50), .A2(new_n788), .B1(new_n700), .B2(G68), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n280), .B1(new_n202), .B2(new_n719), .C1(new_n789), .C2(KEYINPUT103), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(KEYINPUT103), .B2(new_n789), .ZN(new_n791));
  INV_X1    g0591(.A(G132), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n787), .B(new_n791), .C1(new_n792), .C2(new_n706), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n706), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n724), .A2(new_n218), .B1(new_n796), .B2(new_n694), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(KEYINPUT102), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT102), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n713), .A2(new_n515), .B1(new_n719), .B2(new_n222), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n716), .A2(new_n224), .B1(new_n699), .B2(new_n342), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n317), .B1(new_n711), .B2(new_n455), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n798), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n793), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n763), .B1(new_n805), .B2(new_n692), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n743), .A2(new_n692), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n283), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(new_n744), .C2(new_n774), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n782), .A2(new_n809), .ZN(G384));
  NOR2_X1   g0610(.A1(new_n407), .A2(new_n629), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT39), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n329), .A2(new_n337), .ZN(new_n814));
  INV_X1    g0614(.A(new_n627), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n357), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n813), .B1(new_n816), .B2(new_n348), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n350), .B1(new_n361), .B2(new_n627), .ZN(new_n818));
  INV_X1    g0618(.A(new_n348), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n817), .B1(new_n820), .B2(new_n813), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT107), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n595), .A2(new_n599), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n814), .A2(new_n815), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n823), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(KEYINPUT107), .B(new_n825), .C1(new_n595), .C2(new_n599), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(KEYINPUT38), .B(new_n822), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n812), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n820), .A2(new_n813), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT37), .B1(new_n818), .B2(new_n819), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n350), .A2(new_n627), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n824), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT38), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n840), .A2(new_n832), .A3(new_n812), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n811), .B1(new_n833), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n831), .A2(new_n832), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n393), .A2(new_n629), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n407), .A2(new_n396), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n393), .B(new_n629), .C1(new_n597), .C2(new_n406), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT106), .ZN(new_n848));
  INV_X1    g0648(.A(new_n770), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n779), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g0650(.A(KEYINPUT106), .B(new_n770), .C1(new_n776), .C2(new_n778), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n843), .B(new_n847), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n600), .A2(new_n627), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n842), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n425), .A2(new_n663), .A3(new_n668), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n602), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n854), .B(new_n856), .Z(new_n857));
  AOI21_X1  g0657(.A(new_n683), .B1(KEYINPUT108), .B2(new_n681), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n681), .A2(KEYINPUT108), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(new_n859), .C1(new_n686), .C2(new_n688), .ZN(new_n860));
  INV_X1    g0660(.A(new_n774), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n845), .B2(new_n846), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT40), .B1(new_n843), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT107), .B1(new_n363), .B2(new_n825), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n824), .A2(new_n823), .A3(new_n826), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n821), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n839), .B1(new_n867), .B2(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n860), .A2(new_n862), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT40), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n425), .A2(new_n860), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(G330), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n857), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n212), .B2(new_n623), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n218), .B1(new_n564), .B2(KEYINPUT35), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n878), .B(new_n239), .C1(KEYINPUT35), .C2(new_n564), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT36), .ZN(new_n880));
  OAI21_X1  g0680(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n649), .A2(new_n881), .B1(G50), .B2(new_n203), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(G1), .A3(new_n622), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n877), .A2(new_n880), .A3(new_n883), .ZN(G367));
  OAI21_X1  g0684(.A(new_n658), .B1(new_n574), .B2(new_n631), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n633), .A2(new_n640), .A3(new_n886), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n887), .A2(KEYINPUT42), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n888), .A2(KEYINPUT111), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(KEYINPUT42), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(KEYINPUT111), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n480), .B1(new_n576), .B2(new_n657), .ZN(new_n892));
  INV_X1    g0692(.A(new_n583), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n631), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n889), .A2(new_n890), .A3(new_n891), .A4(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n508), .A2(new_n631), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT109), .Z(new_n897));
  MUX2_X1   g0697(.A(new_n505), .B(new_n607), .S(new_n897), .Z(new_n898));
  INV_X1    g0698(.A(KEYINPUT43), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT112), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT113), .ZN(new_n903));
  INV_X1    g0703(.A(new_n638), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n885), .B1(new_n583), .B2(new_n631), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT114), .Z(new_n907));
  XNOR2_X1  g0707(.A(new_n903), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n898), .B(KEYINPUT110), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n899), .B(new_n909), .C1(new_n902), .C2(KEYINPUT113), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n910), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n644), .B(KEYINPUT41), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n641), .A2(new_n905), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT45), .Z(new_n916));
  NOR2_X1   g0716(.A1(new_n641), .A2(new_n905), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT44), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n904), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n904), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n633), .B(new_n640), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(new_n637), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n690), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n914), .B1(new_n928), .B2(new_n690), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n911), .B(new_n912), .C1(new_n760), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n898), .A2(new_n745), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n746), .B1(new_n235), .B2(new_n416), .C1(new_n251), .C2(new_n752), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n280), .B1(new_n694), .B2(new_n730), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n734), .A2(G68), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n785), .B2(new_n713), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(G137), .C2(new_n707), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n788), .A2(G58), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n725), .A2(G50), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n699), .A2(new_n283), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G150), .B2(new_n737), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n936), .A2(new_n937), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n716), .A2(new_n218), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT46), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G311), .B2(new_n714), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n694), .A2(new_n455), .B1(new_n719), .B2(new_n224), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n711), .A2(new_n515), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n699), .A2(new_n222), .ZN(new_n947));
  NOR4_X1   g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n280), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n944), .B(new_n948), .C1(new_n796), .C2(new_n724), .ZN(new_n949));
  INV_X1    g0749(.A(G317), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n706), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n941), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n763), .B1(new_n953), .B2(new_n692), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n931), .A2(new_n932), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n930), .A2(new_n955), .ZN(G387));
  NAND2_X1  g0756(.A1(new_n925), .A2(new_n760), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n783), .A2(G311), .B1(new_n714), .B2(G322), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n950), .B2(new_n711), .C1(new_n724), .C2(new_n515), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT48), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n796), .B2(new_n719), .C1(new_n455), .C2(new_n716), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT49), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n707), .A2(G326), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n962), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n280), .B1(new_n700), .B2(G116), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n716), .A2(new_n283), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G150), .B2(new_n707), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n203), .B2(new_n702), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n947), .B(new_n970), .C1(G50), .C2(new_n737), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n783), .A2(new_n334), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n416), .A2(new_n719), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G159), .B2(new_n714), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n971), .A2(new_n280), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n967), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n763), .B1(new_n976), .B2(new_n692), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n647), .B(new_n298), .C1(new_n203), .C2(new_n283), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT115), .Z(new_n979));
  NOR2_X1   g0779(.A1(new_n269), .A2(G50), .ZN(new_n980));
  XOR2_X1   g0780(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n751), .B1(new_n979), .B2(new_n982), .C1(new_n248), .C2(new_n298), .ZN(new_n983));
  INV_X1    g0783(.A(new_n748), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(G107), .B2(new_n235), .C1(new_n647), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n746), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n977), .B(new_n986), .C1(new_n633), .C2(new_n757), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n644), .B1(new_n690), .B2(new_n925), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n957), .B(new_n987), .C1(new_n927), .C2(new_n988), .ZN(G393));
  INV_X1    g0789(.A(new_n922), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n920), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n759), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n905), .A2(new_n757), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n746), .B1(new_n222), .B2(new_n235), .C1(new_n258), .C2(new_n752), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n724), .A2(new_n269), .B1(new_n216), .B2(new_n694), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT117), .Z(new_n996));
  INV_X1    g0796(.A(G150), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n713), .A2(new_n997), .B1(new_n711), .B2(new_n730), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT51), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n280), .B1(new_n699), .B2(new_n342), .C1(new_n203), .C2(new_n716), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n719), .A2(new_n283), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n996), .B(new_n1004), .C1(new_n785), .C2(new_n706), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n713), .A2(new_n950), .B1(new_n711), .B2(new_n794), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT52), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n694), .A2(new_n515), .B1(new_n699), .B2(new_n224), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n716), .A2(new_n796), .B1(new_n706), .B2(new_n709), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n317), .B1(new_n719), .B2(new_n218), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1007), .B(new_n1011), .C1(new_n455), .C2(new_n702), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1005), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n763), .B1(new_n1013), .B2(new_n692), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n993), .A2(new_n994), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT118), .B1(new_n992), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT118), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1018), .B(new_n1015), .C1(new_n991), .C2(new_n759), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n991), .A2(new_n926), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n928), .A2(new_n1021), .A3(new_n644), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(G390));
  NAND3_X1  g0823(.A1(new_n425), .A2(G330), .A3(new_n860), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n602), .A2(new_n855), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n861), .A2(new_n634), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n847), .B1(new_n689), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n860), .A2(new_n1026), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n847), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1027), .A2(new_n1030), .B1(new_n850), .B2(new_n851), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT119), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n773), .A2(new_n420), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n662), .A2(new_n631), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n849), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n689), .A2(new_n847), .A3(new_n1026), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1028), .A2(KEYINPUT119), .A3(new_n1029), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1034), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1025), .B1(new_n1031), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n865), .A2(new_n866), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT38), .B1(new_n1043), .B2(new_n822), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n830), .B(new_n821), .C1(new_n865), .C2(new_n866), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT39), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n868), .A2(new_n812), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n811), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1037), .A2(new_n847), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n868), .A2(new_n811), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1051), .A2(new_n1055), .A3(new_n1039), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n833), .A2(new_n841), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n777), .B1(new_n666), .B2(new_n774), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n778), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n849), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT106), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n779), .A2(new_n848), .A3(new_n849), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1029), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1057), .B1(new_n1063), .B2(new_n811), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1030), .B1(new_n1064), .B2(new_n1054), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1042), .B1(new_n1056), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1030), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1041), .A2(new_n1031), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1025), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1039), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1064), .A2(new_n1054), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1068), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1066), .A2(new_n644), .A3(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n694), .A2(new_n224), .B1(new_n713), .B2(new_n796), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n317), .B1(new_n699), .B2(new_n203), .C1(new_n342), .C2(new_n716), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n725), .C2(G97), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1003), .B1(G116), .B2(new_n737), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT121), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n455), .C2(new_n706), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT122), .Z(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT54), .B(G143), .Z(new_n1083));
  NAND2_X1  g0883(.A1(new_n725), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(G128), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n713), .A2(new_n1085), .B1(new_n711), .B2(new_n792), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT120), .ZN(new_n1087));
  INV_X1    g0887(.A(G125), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n280), .B1(new_n706), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G137), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n694), .A2(new_n1090), .B1(new_n719), .B2(new_n730), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(G50), .C2(new_n700), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1084), .A2(new_n1087), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n788), .A2(G150), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1082), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n763), .B1(new_n1096), .B2(new_n692), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1048), .B2(new_n744), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n269), .B2(new_n807), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n760), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1075), .A2(new_n1101), .ZN(G378));
  INV_X1    g0902(.A(KEYINPUT57), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n864), .A2(new_n871), .A3(new_n634), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n854), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT56), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n278), .A2(new_n815), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n314), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT55), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n314), .A2(new_n1107), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1106), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT55), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(KEYINPUT56), .A3(new_n1111), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n840), .A2(new_n832), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n863), .A2(KEYINPUT40), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n869), .B1(new_n832), .B2(new_n831), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1120), .B(G330), .C1(new_n1121), .C2(KEYINPUT40), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1122), .A2(new_n853), .A3(new_n852), .A4(new_n842), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n1105), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1118), .B1(new_n1105), .B2(new_n1123), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1025), .B1(new_n1100), .B2(new_n1069), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1103), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1105), .A2(new_n1123), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1118), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1105), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1129), .A2(new_n1134), .A3(KEYINPUT57), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1128), .A2(new_n1135), .A3(new_n644), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n760), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n807), .A2(new_n216), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n934), .B1(new_n222), .B2(new_n694), .C1(new_n218), .C2(new_n713), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n1139), .A2(G41), .A3(new_n280), .A4(new_n968), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n416), .A2(new_n702), .B1(new_n699), .B2(new_n202), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G107), .B2(new_n737), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n796), .C2(new_n706), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT58), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n216), .B1(new_n315), .B2(G41), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n711), .A2(new_n1085), .B1(new_n702), .B2(new_n1090), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n788), .B2(new_n1083), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n783), .A2(G132), .B1(new_n714), .B2(G125), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n997), .C2(new_n719), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT59), .Z(new_n1150));
  AOI21_X1  g0950(.A(G41), .B1(new_n707), .B2(G124), .ZN(new_n1151));
  AOI21_X1  g0951(.A(G33), .B1(new_n700), .B2(G159), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1144), .A2(new_n1145), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n763), .B1(new_n1154), .B2(new_n692), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1138), .B(new_n1155), .C1(new_n1131), .C2(new_n744), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1137), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1136), .A2(new_n1158), .ZN(G375));
  AOI21_X1  g0959(.A(new_n759), .B1(new_n1041), .B2(new_n1031), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(KEYINPUT123), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1029), .A2(new_n743), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n807), .A2(new_n203), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n724), .A2(new_n224), .B1(new_n218), .B2(new_n694), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT124), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n711), .A2(new_n796), .B1(new_n706), .B2(new_n515), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1167), .B(new_n973), .C1(G97), .C2(new_n788), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1165), .A2(KEYINPUT124), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n280), .B(new_n939), .C1(G294), .C2(new_n714), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n711), .A2(new_n1090), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n783), .A2(new_n1083), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n216), .B2(new_n719), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G132), .B2(new_n714), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n280), .B1(new_n702), .B2(new_n997), .C1(new_n202), .C2(new_n699), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n716), .A2(new_n730), .B1(new_n706), .B2(new_n1085), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1176), .B1(KEYINPUT125), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1175), .B(new_n1178), .C1(KEYINPUT125), .C2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1171), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n763), .B1(new_n1180), .B2(new_n692), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1163), .A2(new_n1164), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1160), .A2(KEYINPUT123), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1162), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1025), .A2(new_n1041), .A3(new_n1031), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1185), .A2(new_n913), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n1071), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(G381));
  INV_X1    g0988(.A(G390), .ZN(new_n1189));
  INV_X1    g0989(.A(G384), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(G387), .A2(new_n1191), .A3(G396), .A4(G393), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n1101), .A2(new_n1075), .A3(new_n1137), .A4(new_n1156), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n1136), .A3(new_n1187), .A4(new_n1193), .ZN(G407));
  NAND2_X1  g0994(.A1(new_n1136), .A2(new_n1193), .ZN(new_n1195));
  OAI211_X1 g0995(.A(G407), .B(G213), .C1(G343), .C2(new_n1195), .ZN(G409));
  INV_X1    g0996(.A(G213), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(G343), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1129), .A2(new_n1134), .A3(new_n913), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT60), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n645), .B1(new_n1185), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1071), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1185), .A2(new_n1201), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1205), .A2(new_n1184), .A3(new_n1190), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1183), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1182), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1207), .A2(new_n1161), .A3(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1202), .B(new_n1071), .C1(new_n1201), .C2(new_n1185), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G384), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1206), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(G378), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1071), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1214), .A2(new_n1025), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n645), .B1(new_n1215), .B2(new_n1103), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1157), .B1(new_n1216), .B2(new_n1135), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1200), .B(new_n1212), .C1(new_n1213), .C2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1198), .A2(G2897), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1190), .B1(new_n1205), .B2(new_n1184), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1209), .A2(new_n1210), .A3(G384), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n1219), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G375), .A2(G378), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n1200), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT63), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1218), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(G393), .B(G396), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1189), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1189), .A2(new_n1230), .ZN(new_n1232));
  AND4_X1   g1032(.A1(new_n955), .A2(new_n1231), .A3(new_n930), .A4(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1231), .A2(new_n1232), .B1(new_n930), .B2(new_n955), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1233), .A2(new_n1234), .A3(KEYINPUT61), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT126), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1218), .B2(new_n1228), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1198), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1075), .A2(new_n1137), .A3(new_n1156), .A4(new_n1101), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1215), .A2(new_n914), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G375), .B2(G378), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1242), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1212), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1229), .A2(new_n1235), .A3(new_n1237), .A4(new_n1243), .ZN(new_n1244));
  XOR2_X1   g1044(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1245));
  NAND2_X1  g1045(.A1(new_n1193), .A2(new_n1199), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1238), .B(new_n1246), .C1(new_n1217), .C2(new_n1213), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1218), .A2(KEYINPUT62), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1242), .A2(new_n1251), .A3(new_n1212), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1244), .A2(new_n1256), .ZN(G405));
  NAND2_X1  g1057(.A1(new_n1226), .A2(new_n1195), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1212), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1226), .B(new_n1195), .C1(new_n1211), .C2(new_n1206), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1254), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1254), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(G402));
endmodule


