//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n440, new_n441, new_n445, new_n446, new_n447,
    new_n453, new_n457, new_n458, new_n459, new_n460, new_n461, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n439));
  OR2_X1    g014(.A1(new_n439), .A2(G69), .ZN(new_n440));
  NAND2_X1  g015(.A1(new_n439), .A2(G69), .ZN(new_n441));
  NAND2_X1  g016(.A1(new_n440), .A2(new_n441), .ZN(G235));
  INV_X1    g017(.A(G120), .ZN(G236));
  INV_X1    g018(.A(G57), .ZN(G237));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n445));
  OR2_X1    g020(.A1(new_n445), .A2(G108), .ZN(new_n446));
  NAND2_X1  g021(.A1(new_n445), .A2(G108), .ZN(new_n447));
  NAND2_X1  g022(.A1(new_n446), .A2(new_n447), .ZN(G238));
  NAND4_X1  g023(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g024(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g025(.A(G452), .Z(G391));
  AND2_X1   g026(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g027(.A1(G7), .A2(G661), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g029(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g030(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g031(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT2), .Z(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR4_X1   g034(.A1(G235), .A2(G238), .A3(G237), .A4(G236), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(G325));
  INV_X1    g037(.A(G325), .ZN(G261));
  NAND2_X1  g038(.A1(new_n461), .A2(G567), .ZN(new_n464));
  INV_X1    g039(.A(G2106), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n458), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  XNOR2_X1  g042(.A(KEYINPUT67), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT3), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n469), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n484), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n485));
  OR2_X1    g060(.A1(new_n485), .A2(new_n480), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  OAI211_X1 g063(.A(new_n480), .B(new_n476), .C1(new_n468), .C2(new_n475), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n476), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n470), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n493), .B1(new_n496), .B2(KEYINPUT3), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n492), .A2(G136), .B1(G124), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(G100), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(new_n480), .B2(G112), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XOR2_X1   g078(.A(new_n503), .B(KEYINPUT69), .Z(G162));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR4_X1   g080(.A1(new_n483), .A2(KEYINPUT4), .A3(new_n505), .A4(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n489), .B2(new_n505), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n474), .A2(G138), .A3(new_n480), .A4(new_n476), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT70), .A3(KEYINPUT4), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n506), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n480), .A2(G102), .A3(G2104), .ZN(new_n513));
  NAND2_X1  g088(.A1(G114), .A2(G2104), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n497), .B2(G126), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n516), .B2(new_n480), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n512), .A2(new_n517), .ZN(G164));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(KEYINPUT72), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT71), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  AND2_X1   g101(.A1(G75), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(G543), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT5), .B(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n525), .A2(G88), .ZN(new_n530));
  AND2_X1   g105(.A1(G62), .A2(G651), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  AND2_X1   g109(.A1(new_n529), .A2(KEYINPUT73), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n529), .A2(KEYINPUT73), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G63), .ZN(new_n538));
  NAND2_X1  g113(.A1(G76), .A2(G543), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n522), .A2(G543), .A3(new_n523), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G51), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n522), .A2(new_n523), .A3(new_n529), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT75), .B(G89), .Z(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n540), .B1(new_n520), .B2(new_n539), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n542), .A2(new_n545), .A3(new_n549), .A4(new_n550), .ZN(G286));
  INV_X1    g126(.A(G286), .ZN(G168));
  INV_X1    g127(.A(new_n537), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n520), .ZN(new_n555));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  INV_X1    g131(.A(G90), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n556), .A2(new_n543), .B1(new_n546), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(G171));
  AOI22_X1  g134(.A1(new_n553), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n520), .ZN(new_n561));
  INV_X1    g136(.A(G43), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n543), .B1(new_n546), .B2(new_n563), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(G188));
  AOI21_X1  g147(.A(KEYINPUT9), .B1(new_n544), .B2(G53), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  NOR3_X1   g150(.A1(new_n543), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  XOR2_X1   g153(.A(KEYINPUT5), .B(G543), .Z(new_n579));
  XNOR2_X1  g154(.A(KEYINPUT76), .B(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n547), .A2(G91), .B1(G651), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n585), .A2(new_n543), .B1(new_n546), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n520), .B1(new_n537), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  AND2_X1   g166(.A1(new_n529), .A2(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT77), .Z(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n546), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G48), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n543), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  AOI22_X1  g176(.A1(new_n553), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n520), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n604), .A2(new_n543), .B1(new_n546), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n579), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n544), .A2(G54), .B1(G651), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OR3_X1    g188(.A1(new_n546), .A2(KEYINPUT10), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT10), .B1(new_n546), .B2(new_n613), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G171), .B2(new_n617), .ZN(G284));
  OAI21_X1  g194(.A(new_n618), .B1(G171), .B2(new_n617), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(G299), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G297));
  OAI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(new_n616), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n565), .A2(new_n617), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n616), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n499), .A2(G123), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT78), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n492), .A2(G135), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT79), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G111), .B2(new_n480), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n633), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NOR3_X1   g214(.A1(new_n483), .A2(new_n496), .A3(G2105), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT12), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2435), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2438), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(G14), .ZN(G401));
  XNOR2_X1  g232(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(G2096), .Z(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(new_n658), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT81), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n682), .A2(new_n675), .A3(new_n677), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n683), .C1(new_n677), .C2(new_n682), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT22), .B(G1981), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NOR2_X1   g267(.A1(G286), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n694), .B(KEYINPUT91), .C1(G16), .C2(G21), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(KEYINPUT91), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1966), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(G29), .A2(G32), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n492), .A2(G141), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n499), .A2(G129), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n468), .A2(G105), .A3(new_n480), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT26), .Z(new_n704));
  NAND4_X1  g279(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n699), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT27), .B(G1996), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n698), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT28), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n706), .A2(G26), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n492), .A2(G140), .B1(G128), .B2(new_n499), .ZN(new_n712));
  OR2_X1    g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AOI211_X1 g290(.A(new_n710), .B(new_n711), .C1(new_n715), .C2(G29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n710), .B2(new_n711), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT89), .B(G2067), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n707), .A2(new_n708), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n692), .A2(KEYINPUT23), .A3(G20), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n723));
  INV_X1    g298(.A(G20), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G16), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n725), .C1(new_n622), .C2(new_n692), .ZN(new_n726));
  INV_X1    g301(.A(G1956), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n566), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G16), .B2(G19), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n728), .B1(G1341), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G164), .A2(new_n706), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G27), .B2(new_n706), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR4_X1   g311(.A1(new_n709), .A2(new_n721), .A3(new_n732), .A4(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n706), .A2(G33), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  INV_X1    g314(.A(G127), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n483), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2105), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT25), .Z(new_n746));
  INV_X1    g321(.A(G139), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n746), .C1(new_n747), .C2(new_n491), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n738), .B1(new_n748), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G2072), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n731), .A2(G1341), .ZN(new_n752));
  NOR2_X1   g327(.A1(G5), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G171), .B2(G16), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G1961), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n638), .A2(new_n706), .B1(new_n749), .B2(new_n750), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT92), .B(G28), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT30), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n754), .A2(G1961), .B1(new_n706), .B2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n760), .A2(new_n706), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n706), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n752), .A2(new_n755), .A3(new_n756), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n734), .A2(new_n735), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n737), .A2(new_n751), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G22), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G166), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1971), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n692), .A2(G23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n590), .B2(new_n692), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT86), .B(KEYINPUT33), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1976), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n775), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n692), .A2(G6), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n600), .B2(new_n692), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT85), .B(G1981), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n780), .B(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n773), .A2(new_n778), .A3(new_n783), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT87), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT34), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n492), .A2(G131), .B1(G119), .B2(new_n499), .ZN(new_n787));
  OR2_X1    g362(.A1(G95), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G107), .C2(new_n480), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT84), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(KEYINPUT84), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(new_n706), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G25), .B2(new_n706), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT35), .B(G1991), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n692), .A2(G24), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n607), .B2(new_n692), .ZN(new_n801));
  INV_X1    g376(.A(G1986), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n796), .A2(new_n798), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n786), .A2(new_n799), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT36), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT36), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n769), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G29), .A2(G35), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G162), .B2(G29), .ZN(new_n810));
  INV_X1    g385(.A(G2090), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G4), .A2(G16), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n625), .B2(G16), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT88), .B(G1348), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT31), .B(G11), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n808), .A2(new_n815), .A3(new_n820), .A4(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  AOI22_X1  g398(.A1(G55), .A2(new_n544), .B1(new_n547), .B2(G93), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n553), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n520), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n829), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n566), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n565), .A2(new_n826), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n625), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT39), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n828), .B1(new_n839), .B2(G860), .ZN(G145));
  NAND2_X1  g415(.A1(new_n748), .A2(KEYINPUT97), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n641), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(new_n513), .C1(new_n516), .C2(new_n480), .ZN(new_n844));
  OAI211_X1 g419(.A(G126), .B(new_n476), .C1(new_n468), .C2(new_n475), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n480), .B1(new_n845), .B2(new_n514), .ZN(new_n846));
  INV_X1    g421(.A(new_n513), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT96), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n506), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n510), .A2(KEYINPUT70), .A3(KEYINPUT4), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT70), .B1(new_n510), .B2(KEYINPUT4), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n715), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n842), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n705), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n492), .A2(G142), .B1(G130), .B2(new_n499), .ZN(new_n858));
  NOR2_X1   g433(.A1(G106), .A2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(new_n480), .B2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n793), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n638), .B(new_n487), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G162), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT98), .Z(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n863), .B2(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g445(.A1(new_n826), .A2(new_n617), .ZN(new_n871));
  XNOR2_X1  g446(.A(G303), .B(new_n590), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G290), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n600), .B(KEYINPUT101), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT42), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n622), .A2(new_n616), .ZN(new_n877));
  NAND2_X1  g452(.A1(G299), .A2(new_n625), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT99), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(KEYINPUT41), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n879), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(KEYINPUT100), .A3(KEYINPUT41), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n834), .B(new_n629), .ZN(new_n887));
  MUX2_X1   g462(.A(new_n880), .B(new_n886), .S(new_n887), .Z(new_n888));
  XOR2_X1   g463(.A(new_n876), .B(new_n888), .Z(new_n889));
  OAI21_X1  g464(.A(new_n871), .B1(new_n889), .B2(new_n617), .ZN(G295));
  OAI21_X1  g465(.A(new_n871), .B1(new_n889), .B2(new_n617), .ZN(G331));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  XNOR2_X1  g467(.A(G168), .B(G171), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n834), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n895), .B(new_n896), .C1(new_n884), .C2(new_n894), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n886), .A2(KEYINPUT102), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n875), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n881), .B2(new_n894), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n880), .B2(new_n894), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT103), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n901), .A2(new_n907), .A3(new_n902), .A4(new_n904), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n892), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n897), .A2(new_n875), .A3(new_n898), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n901), .A2(new_n902), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT44), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n901), .A2(new_n892), .A3(new_n902), .A4(new_n904), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n911), .B2(new_n892), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(G397));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT45), .B1(new_n854), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G40), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n487), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n793), .A2(new_n797), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n715), .A2(G2067), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n715), .A2(G2067), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1996), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n705), .B(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n924), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n930), .B2(new_n925), .ZN(new_n931));
  INV_X1    g506(.A(new_n923), .ZN(new_n932));
  INV_X1    g507(.A(new_n927), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n705), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(KEYINPUT46), .A3(new_n928), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n923), .B2(G1996), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n794), .A2(new_n798), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n927), .A2(new_n929), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n941), .A2(new_n942), .A3(new_n924), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(new_n923), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT126), .ZN(new_n945));
  NOR2_X1   g520(.A1(G290), .A2(G1986), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n932), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT48), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n931), .B(new_n940), .C1(new_n945), .C2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT122), .ZN(new_n950));
  OAI211_X1 g525(.A(KEYINPUT45), .B(new_n919), .C1(new_n512), .C2(new_n517), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n922), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n697), .B1(new_n952), .B2(new_n920), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n919), .B1(new_n512), .B2(new_n517), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT50), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n854), .A2(new_n956), .A3(new_n919), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n955), .A2(new_n957), .A3(new_n764), .A4(new_n922), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(G168), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT51), .B1(new_n959), .B2(G8), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n953), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n953), .B2(new_n958), .ZN(new_n963));
  OAI21_X1  g538(.A(G8), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G286), .A2(G8), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT117), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n960), .B1(new_n967), .B2(KEYINPUT51), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n962), .A2(new_n963), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n969), .A2(new_n965), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT121), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G2078), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n920), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n849), .B2(new_n853), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n921), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n481), .B(KEYINPUT119), .Z(new_n979));
  NAND4_X1  g554(.A1(new_n976), .A2(new_n486), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n954), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n854), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n735), .A4(new_n922), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n973), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n955), .A2(new_n957), .A3(new_n922), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT118), .B(G1961), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n980), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G171), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n984), .A2(new_n973), .B1(new_n986), .B2(new_n987), .ZN(new_n991));
  INV_X1    g566(.A(new_n920), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(new_n922), .A3(new_n951), .A4(new_n974), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(G301), .A3(new_n993), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n972), .A2(new_n990), .A3(KEYINPUT54), .A4(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n989), .B2(G171), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n972), .B1(new_n997), .B2(new_n994), .ZN(new_n998));
  OAI22_X1  g573(.A1(new_n968), .A2(new_n971), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n922), .B1(new_n977), .B2(new_n956), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT107), .B(new_n922), .C1(new_n977), .C2(new_n956), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1003), .A2(new_n811), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n982), .A2(new_n983), .A3(new_n922), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n772), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1000), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G303), .A2(G8), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT104), .B(KEYINPUT55), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1010), .B(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n982), .A2(new_n983), .A3(new_n922), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n1015), .A2(G1971), .B1(new_n986), .B2(G2090), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(new_n1013), .A3(G8), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1000), .B1(new_n977), .B2(new_n922), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G288), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n590), .A2(G1976), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT49), .B1(new_n600), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1027), .B(G1981), .C1(new_n597), .C2(new_n599), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT106), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n600), .A2(new_n1025), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1030), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1019), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n854), .A2(new_n922), .A3(new_n919), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(G8), .A3(new_n1023), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT105), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT52), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1037), .B2(KEYINPUT52), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1024), .B(new_n1035), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1014), .A2(new_n1018), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n985), .A2(new_n993), .A3(new_n988), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G171), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n991), .A2(G301), .A3(new_n980), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1043), .B1(new_n1047), .B2(new_n996), .ZN(new_n1048));
  AOI211_X1 g623(.A(KEYINPUT120), .B(KEYINPUT54), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1042), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n950), .B1(new_n999), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1036), .A2(G2067), .ZN(new_n1052));
  INV_X1    g627(.A(G1348), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n986), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT60), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n616), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(KEYINPUT115), .B(new_n625), .C1(new_n1054), .C2(KEYINPUT60), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1057), .A2(new_n1058), .B1(new_n1056), .B2(new_n1055), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1054), .A2(KEYINPUT60), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n577), .B(KEYINPUT110), .ZN(new_n1063));
  XOR2_X1   g638(.A(new_n582), .B(KEYINPUT111), .Z(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT112), .B(new_n1062), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1067), .B(new_n1068), .C1(new_n1062), .C2(G299), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n727), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT109), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(KEYINPUT109), .A3(new_n727), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n982), .A2(new_n983), .A3(new_n922), .A4(new_n1075), .ZN(new_n1076));
  XOR2_X1   g651(.A(new_n1076), .B(KEYINPUT113), .Z(new_n1077));
  NAND4_X1  g652(.A1(new_n1069), .A2(new_n1073), .A3(new_n1074), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT61), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1036), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1007), .B2(G1996), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(KEYINPUT114), .A3(new_n566), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT59), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1074), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT109), .B1(new_n1070), .B2(new_n727), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n1069), .A4(new_n1077), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1061), .A2(new_n1079), .A3(new_n1084), .A4(new_n1089), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1073), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1091), .A2(new_n1069), .B1(new_n616), .B2(new_n1054), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1078), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1041), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(new_n1017), .C1(new_n1009), .C2(new_n1013), .ZN(new_n1096));
  AND4_X1   g671(.A1(G301), .A2(new_n980), .A3(new_n985), .A4(new_n988), .ZN(new_n1097));
  AOI21_X1  g672(.A(G301), .B1(new_n991), .B2(new_n993), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n996), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT120), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1047), .A2(new_n1043), .A3(new_n996), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(new_n964), .B2(new_n966), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n970), .B1(new_n1104), .B2(new_n960), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n997), .A2(new_n994), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT121), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n997), .A2(new_n972), .A3(new_n994), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1102), .A2(KEYINPUT122), .A3(new_n1105), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1051), .A2(new_n1094), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1035), .A2(new_n1021), .A3(new_n590), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1031), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1019), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1017), .B2(new_n1041), .ZN(new_n1115));
  AOI211_X1 g690(.A(new_n1000), .B(G286), .C1(new_n953), .C2(new_n958), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1042), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1118), .A2(KEYINPUT108), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(KEYINPUT108), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1013), .B1(new_n1016), .B2(G8), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n1118), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(new_n1017), .A3(new_n1095), .A4(new_n1116), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1115), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(new_n970), .C1(new_n1104), .C2(new_n960), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1096), .A2(new_n1045), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT123), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1105), .A2(KEYINPUT62), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1111), .A2(new_n1125), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n943), .B1(new_n802), .B2(new_n607), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n932), .B1(new_n1136), .B2(new_n946), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1135), .A2(KEYINPUT124), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT124), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n949), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT127), .B(new_n949), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g719(.A1(new_n915), .A2(G319), .A3(new_n690), .ZN(new_n1146));
  NOR2_X1   g720(.A1(G401), .A2(G227), .ZN(new_n1147));
  NAND2_X1  g721(.A1(new_n869), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1148), .ZN(G308));
  OR2_X1    g723(.A1(new_n1146), .A2(new_n1148), .ZN(G225));
endmodule


