//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202));
  INV_X1    g001(.A(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(G228gat), .ZN(new_n204));
  INV_X1    g003(.A(G233gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G141gat), .B(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT72), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT72), .B1(new_n217), .B2(new_n209), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n208), .B(new_n210), .C1(new_n214), .C2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n209), .B(new_n217), .C1(new_n207), .C2(KEYINPUT2), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n222), .A2(KEYINPUT80), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT80), .B1(new_n222), .B2(new_n223), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT22), .ZN(new_n227));
  INV_X1    g026(.A(G211gat), .ZN(new_n228));
  INV_X1    g027(.A(G218gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G211gat), .B(G218gat), .Z(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n224), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n233), .B2(new_n223), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n221), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n206), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n206), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n235), .B2(new_n237), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n233), .B1(new_n222), .B2(new_n223), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n203), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n223), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n233), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n222), .A2(KEYINPUT80), .A3(new_n223), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n235), .A2(new_n237), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n240), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n253), .A2(G22gat), .A3(new_n243), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n202), .B1(new_n245), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n203), .A3(new_n244), .ZN(new_n256));
  OAI21_X1  g055(.A(G22gat), .B1(new_n253), .B2(new_n243), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT81), .ZN(new_n258));
  XNOR2_X1  g057(.A(G78gat), .B(G106gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT79), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT31), .B(G50gat), .Z(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  NAND3_X1  g061(.A1(new_n255), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n202), .B(new_n264), .C1(new_n245), .C2(new_n254), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT40), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  INV_X1    g069(.A(G113gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(G120gat), .ZN(new_n272));
  INV_X1    g071(.A(G120gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(G113gat), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n269), .B(new_n270), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G113gat), .B(G120gat), .ZN(new_n276));
  INV_X1    g075(.A(G127gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(G134gat), .ZN(new_n278));
  INV_X1    g077(.A(G134gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(G127gat), .ZN(new_n280));
  OAI22_X1  g079(.A1(new_n276), .A2(KEYINPUT1), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n219), .A2(new_n221), .A3(new_n275), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT4), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n275), .A2(new_n281), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n284), .A2(new_n221), .A3(new_n219), .A4(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(KEYINPUT75), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n282), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n288), .A2(KEYINPUT76), .A3(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n222), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT73), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n296), .A2(new_n300), .A3(new_n297), .A4(new_n222), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n294), .A2(new_n295), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT39), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n236), .A2(new_n297), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n306), .A2(new_n282), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n303), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n304), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G1gat), .B(G29gat), .ZN(new_n312));
  INV_X1    g111(.A(G85gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT0), .B(G57gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n299), .A2(new_n301), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n288), .A2(KEYINPUT76), .A3(new_n291), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT76), .B1(new_n288), .B2(new_n291), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n309), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n317), .B1(new_n322), .B2(KEYINPUT39), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n268), .B1(new_n311), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n304), .B2(new_n305), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n322), .B(KEYINPUT39), .C1(new_n309), .C2(new_n308), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(new_n326), .C1(new_n267), .C2(KEYINPUT40), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  AND2_X1   g128(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT65), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT64), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT27), .B(G183gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(new_n329), .ZN(new_n336));
  OAI211_X1 g135(.A(KEYINPUT28), .B(new_n333), .C1(new_n336), .C2(KEYINPUT65), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(G169gat), .B2(G176gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT26), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n339), .A2(KEYINPUT66), .A3(new_n340), .A4(new_n342), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT65), .B1(new_n332), .B2(KEYINPUT64), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n337), .A2(new_n345), .A3(new_n346), .A4(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n352), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n340), .A2(KEYINPUT24), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n359), .A4(new_n360), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n366), .A2(new_n223), .B1(G226gat), .B2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(G226gat), .A3(G233gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT70), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n366), .A2(new_n371), .A3(G226gat), .A4(G233gat), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n368), .A2(new_n370), .A3(new_n249), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n369), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n233), .B1(new_n374), .B2(new_n367), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(KEYINPUT30), .A3(new_n380), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n376), .A2(KEYINPUT71), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT71), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n373), .A2(new_n387), .A3(new_n375), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n388), .A3(new_n379), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n302), .A2(new_n390), .A3(new_n391), .A4(new_n303), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n391), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT77), .B1(new_n393), .B2(new_n309), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n309), .B1(new_n289), .B2(KEYINPUT4), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n318), .B(new_n395), .C1(new_n289), .C2(new_n285), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n396), .B(KEYINPUT5), .C1(new_n303), .C2(new_n307), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n385), .A2(new_n389), .B1(new_n398), .B2(new_n316), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n266), .B1(new_n328), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT37), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n380), .B1(new_n376), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT38), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n368), .A2(new_n249), .A3(new_n369), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n368), .A2(new_n370), .A3(new_n372), .ZN(new_n405));
  OAI211_X1 g204(.A(KEYINPUT37), .B(new_n404), .C1(new_n405), .C2(new_n249), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n398), .B2(new_n316), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n392), .A2(new_n394), .A3(new_n397), .A4(new_n317), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n409), .A2(new_n412), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n386), .A2(KEYINPUT37), .A3(new_n388), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n402), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(KEYINPUT38), .ZN(new_n419));
  AOI211_X1 g218(.A(KEYINPUT83), .B(new_n403), .C1(new_n417), .C2(new_n402), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n381), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n400), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n366), .A2(new_n297), .ZN(new_n423));
  NAND2_X1  g222(.A1(G227gat), .A2(G233gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n350), .A2(new_n365), .A3(new_n284), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n424), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n350), .A2(new_n284), .A3(new_n365), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n284), .B1(new_n350), .B2(new_n365), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT32), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G15gat), .B(G43gat), .ZN(new_n438));
  INV_X1    g237(.A(G71gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT67), .ZN(new_n441));
  INV_X1    g240(.A(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n435), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n443), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n434), .B(KEYINPUT32), .C1(new_n445), .C2(new_n436), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n430), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n430), .A3(new_n446), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT69), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT69), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT36), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n444), .A2(new_n430), .A3(new_n446), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n447), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n456), .A2(KEYINPUT36), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n398), .A2(new_n316), .ZN(new_n459));
  INV_X1    g258(.A(new_n408), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n410), .A2(new_n411), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n409), .A2(new_n412), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n389), .A2(new_n384), .A3(new_n383), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n266), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n422), .A2(new_n458), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n413), .A2(new_n414), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  AND4_X1   g271(.A1(new_n472), .A2(new_n456), .A3(new_n263), .A4(new_n265), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n470), .A2(new_n471), .A3(new_n466), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n266), .B1(new_n452), .B2(new_n450), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(new_n463), .A3(new_n464), .A4(new_n466), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT35), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n463), .A2(new_n473), .A3(new_n464), .A4(new_n466), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n469), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G64gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(G57gat), .ZN(new_n483));
  INV_X1    g282(.A(G57gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n484), .A2(G64gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT89), .ZN(new_n486));
  OAI22_X1  g285(.A1(new_n483), .A2(new_n485), .B1(new_n486), .B2(KEYINPUT9), .ZN(new_n487));
  NAND2_X1  g286(.A1(G71gat), .A2(G78gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT89), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n487), .B(new_n489), .C1(G71gat), .C2(G78gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n482), .A2(KEYINPUT91), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n482), .A2(KEYINPUT91), .ZN(new_n494));
  OAI21_X1  g293(.A(G57gat), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(KEYINPUT92), .C1(G57gat), .C2(new_n482), .ZN(new_n496));
  INV_X1    g295(.A(G78gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n439), .A2(new_n497), .A3(KEYINPUT9), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n488), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n496), .B(new_n499), .C1(KEYINPUT92), .C2(new_n495), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT21), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(G1gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT16), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(G1gat), .B2(new_n504), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(G8gat), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n502), .A2(new_n503), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n503), .B1(new_n502), .B2(new_n510), .ZN(new_n513));
  OAI211_X1 g312(.A(G231gat), .B(G233gat), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n513), .ZN(new_n515));
  NAND2_X1  g314(.A1(G231gat), .A2(G233gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n511), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G183gat), .B(G211gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n501), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G127gat), .B(G155gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n521), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n514), .A2(new_n527), .A3(new_n517), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n522), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n522), .B2(new_n528), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G134gat), .B(G162gat), .Z(new_n533));
  NAND3_X1  g332(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT96), .B(G92gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n313), .ZN(new_n537));
  INV_X1    g336(.A(G106gat), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT8), .B1(new_n442), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G99gat), .B(G106gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT97), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n535), .A2(new_n537), .A3(new_n541), .A4(new_n539), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n544), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G43gat), .B(G50gat), .Z(new_n549));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n549), .A2(new_n550), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  NOR3_X1   g352(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n551), .B(new_n553), .C1(new_n556), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G29gat), .A2(G36gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n558), .B2(new_n554), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT15), .A3(new_n552), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n548), .A2(new_n563), .B1(KEYINPUT41), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n563), .B(KEYINPUT17), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n547), .A3(new_n546), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n564), .A2(KEYINPUT41), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n571), .B1(new_n567), .B2(new_n569), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n533), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n574), .ZN(new_n576));
  INV_X1    g375(.A(new_n533), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n575), .A2(new_n578), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n532), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n481), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n492), .A2(new_n500), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n548), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n543), .A2(new_n545), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n492), .A2(new_n591), .A3(new_n500), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT10), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n501), .A2(KEYINPUT10), .A3(new_n548), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n588), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n588), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT99), .B(G120gat), .Z(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT100), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n595), .B2(new_n597), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n563), .A2(KEYINPUT17), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n559), .B2(new_n562), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n510), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n509), .A2(new_n563), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT18), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n509), .B(new_n563), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n614), .B(KEYINPUT13), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n612), .B1(new_n568), .B2(new_n510), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT18), .B1(new_n620), .B2(new_n614), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n621), .B2(KEYINPUT88), .ZN(new_n622));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623));
  INV_X1    g422(.A(G197gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT11), .B(G169gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n614), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT18), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT88), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n619), .A2(KEYINPUT87), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT87), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n615), .A2(new_n635), .A3(new_n618), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n628), .B(KEYINPUT85), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n622), .A2(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n607), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n587), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n470), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n505), .ZN(G1324gat));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n467), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(G8gat), .B1(new_n641), .B2(new_n466), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(G1325gat));
  AOI21_X1  g450(.A(G15gat), .B1(new_n644), .B2(new_n456), .ZN(new_n652));
  INV_X1    g451(.A(new_n458), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n458), .A2(KEYINPUT101), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(G15gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT102), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n652), .B1(new_n644), .B2(new_n659), .ZN(G1326gat));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n266), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n661), .B(KEYINPUT103), .ZN(new_n666));
  INV_X1    g465(.A(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(G1327gat));
  AOI21_X1  g468(.A(new_n584), .B1(new_n469), .B2(new_n480), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n532), .A2(new_n640), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n465), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G29gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n670), .A2(new_n674), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n470), .A2(G29gat), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n677), .A2(KEYINPUT45), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT45), .B1(new_n677), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT104), .ZN(G1328gat));
  NAND3_X1  g482(.A1(new_n672), .A2(new_n467), .A3(new_n674), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G36gat), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n677), .A2(G36gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n467), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n688), .B2(KEYINPUT46), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(KEYINPUT46), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n687), .A2(KEYINPUT105), .A3(new_n691), .A4(new_n467), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n685), .A2(new_n689), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n684), .A2(G36gat), .B1(KEYINPUT46), .B2(new_n688), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n696), .A2(KEYINPUT106), .A3(new_n689), .A4(new_n692), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1329gat));
  NAND3_X1  g497(.A1(new_n672), .A2(new_n653), .A3(new_n674), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G43gat), .ZN(new_n700));
  INV_X1    g499(.A(new_n456), .ZN(new_n701));
  OR3_X1    g500(.A1(new_n677), .A2(G43gat), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(KEYINPUT47), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n671), .B1(new_n481), .B2(new_n585), .ZN(new_n704));
  AOI211_X1 g503(.A(KEYINPUT44), .B(new_n584), .C1(new_n469), .C2(new_n480), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n657), .B(new_n674), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G43gat), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT47), .B1(new_n707), .B2(new_n702), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n710), .B(KEYINPUT47), .C1(new_n707), .C2(new_n702), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n703), .B1(new_n709), .B2(new_n711), .ZN(G1330gat));
  NAND3_X1  g511(.A1(new_n672), .A2(new_n266), .A3(new_n674), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT108), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n672), .A2(new_n715), .A3(new_n266), .A4(new_n674), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(G50gat), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(G50gat), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n670), .A2(new_n718), .A3(new_n266), .A4(new_n674), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(KEYINPUT48), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n713), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n721), .B2(new_n718), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(G1331gat));
  NAND4_X1  g524(.A1(new_n481), .A2(new_n607), .A3(new_n639), .A4(new_n586), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n470), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n484), .ZN(G1332gat));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n726), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n467), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT49), .B(G64gat), .Z(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(G1333gat));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n726), .A2(G71gat), .A3(new_n701), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n730), .A2(new_n657), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n735), .B(new_n737), .C1(new_n738), .C2(new_n439), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n439), .B1(new_n730), .B2(new_n657), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT50), .B1(new_n740), .B2(new_n736), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n730), .A2(new_n266), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g543(.A1(new_n633), .A2(new_n622), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n637), .A2(new_n638), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n531), .A2(new_n747), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n670), .A2(KEYINPUT51), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT51), .B1(new_n670), .B2(new_n748), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n606), .ZN(new_n752));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n465), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n531), .A2(new_n606), .A3(new_n747), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n704), .B2(new_n705), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT110), .B(new_n754), .C1(new_n704), .C2(new_n705), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n470), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n753), .B1(G85gat), .B2(new_n759), .ZN(G1336gat));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n758), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n536), .B1(new_n761), .B2(new_n467), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n466), .A2(G92gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n749), .B2(new_n750), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n750), .A2(new_n765), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n606), .B(new_n764), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT52), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n672), .A2(new_n467), .A3(new_n754), .ZN(new_n770));
  INV_X1    g569(.A(new_n536), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n607), .B(new_n763), .C1(new_n749), .C2(new_n750), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n776), .ZN(G1337gat));
  NAND3_X1  g576(.A1(new_n752), .A2(new_n442), .A3(new_n456), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n655), .A2(new_n656), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n757), .B2(new_n758), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n780), .B2(new_n442), .ZN(G1338gat));
  INV_X1    g580(.A(new_n266), .ZN(new_n782));
  OAI21_X1  g581(.A(G106gat), .B1(new_n755), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n782), .A2(G106gat), .A3(new_n606), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n783), .B(new_n784), .C1(new_n751), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n766), .B2(new_n767), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n761), .A2(new_n266), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(G106gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n790), .B2(new_n784), .ZN(G1339gat));
  AND4_X1   g590(.A1(new_n606), .A2(new_n531), .A3(new_n584), .A4(new_n639), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT10), .ZN(new_n794));
  INV_X1    g593(.A(new_n592), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n492), .A2(new_n500), .B1(new_n546), .B2(new_n547), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n501), .A2(KEYINPUT10), .A3(new_n548), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n596), .A3(new_n798), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n595), .A2(new_n799), .A3(KEYINPUT54), .ZN(new_n800));
  INV_X1    g599(.A(new_n602), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n595), .B2(KEYINPUT54), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n793), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n596), .B1(new_n797), .B2(new_n798), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n602), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n595), .A2(new_n799), .A3(KEYINPUT54), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT55), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(new_n603), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n620), .A2(new_n614), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n616), .A2(new_n617), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n627), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n745), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n810), .A2(new_n582), .A3(new_n583), .A4(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n745), .B(new_n813), .C1(new_n605), .C2(new_n604), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT113), .B(new_n816), .C1(new_n809), .C2(new_n639), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n584), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n747), .A2(new_n603), .A3(new_n808), .A4(new_n803), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT113), .B1(new_n819), .B2(new_n816), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n815), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n792), .B1(new_n821), .B2(new_n532), .ZN(new_n822));
  INV_X1    g621(.A(new_n475), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n470), .A3(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(KEYINPUT115), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n466), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n829), .A2(new_n271), .A3(new_n747), .A4(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n822), .A2(new_n470), .A3(new_n467), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n701), .A2(new_n266), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n639), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT114), .Z(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(G1340gat));
  NOR3_X1   g636(.A1(new_n834), .A2(new_n273), .A3(new_n606), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n829), .A2(new_n607), .A3(new_n830), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n273), .ZN(G1341gat));
  NOR3_X1   g639(.A1(new_n834), .A2(new_n277), .A3(new_n532), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n827), .A2(new_n532), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n277), .ZN(G1342gat));
  NAND2_X1  g642(.A1(new_n585), .A2(new_n279), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n827), .A2(KEYINPUT56), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n834), .B2(new_n584), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT56), .B1(new_n827), .B2(new_n844), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n822), .B2(new_n782), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT117), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n816), .B1(new_n809), .B2(new_n639), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n815), .B1(new_n585), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n792), .B1(new_n854), .B2(new_n532), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n782), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT57), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n858), .B(new_n849), .C1(new_n822), .C2(new_n782), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n851), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n653), .A2(new_n470), .A3(new_n467), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n860), .A2(G141gat), .A3(new_n747), .A4(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(G141gat), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n657), .A2(new_n782), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n832), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n639), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT118), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n867), .B(new_n868), .ZN(G1344gat));
  INV_X1    g668(.A(new_n865), .ZN(new_n870));
  INV_X1    g669(.A(G148gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n607), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n849), .B1(new_n855), .B2(new_n782), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n852), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n584), .A3(new_n817), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n531), .B1(new_n876), .B2(new_n815), .ZN(new_n877));
  OAI211_X1 g676(.A(KEYINPUT57), .B(new_n266), .C1(new_n877), .C2(new_n792), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n606), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n871), .B1(new_n879), .B2(new_n861), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n880), .A2(KEYINPUT119), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT119), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n860), .A2(new_n861), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n885), .B2(new_n606), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n871), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n872), .B1(new_n884), .B2(new_n887), .ZN(G1345gat));
  OAI21_X1  g687(.A(new_n215), .B1(new_n865), .B2(new_n532), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n860), .A2(G155gat), .A3(new_n861), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n532), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT120), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n870), .B2(new_n585), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n885), .A2(new_n216), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n585), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n465), .A2(new_n466), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n833), .B(new_n896), .C1(new_n877), .C2(new_n792), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n639), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n822), .A2(new_n465), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n475), .A2(new_n467), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT121), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(G169gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n898), .B1(new_n903), .B2(new_n639), .ZN(G1348gat));
  INV_X1    g703(.A(new_n902), .ZN(new_n905));
  AOI21_X1  g704(.A(G176gat), .B1(new_n905), .B2(new_n607), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n897), .A2(new_n606), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(G176gat), .B2(new_n907), .ZN(G1349gat));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n531), .A3(new_n335), .ZN(new_n909));
  OAI21_X1  g708(.A(G183gat), .B1(new_n897), .B2(new_n532), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n897), .B2(new_n584), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT61), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n905), .A2(new_n329), .A3(new_n585), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1351gat));
  NAND2_X1  g715(.A1(new_n779), .A2(new_n896), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n779), .A2(new_n919), .A3(new_n896), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n873), .ZN(new_n922));
  INV_X1    g721(.A(new_n878), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n624), .A3(new_n639), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n917), .A2(new_n782), .A3(new_n822), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n747), .ZN(new_n928));
  OR3_X1    g727(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n925), .B2(new_n928), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1352gat));
  INV_X1    g730(.A(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n927), .A2(new_n932), .A3(new_n607), .ZN(new_n933));
  XNOR2_X1  g732(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n921), .A2(new_n879), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n935), .B(new_n936), .C1(new_n932), .C2(new_n937), .ZN(G1353gat));
  OAI211_X1 g737(.A(new_n921), .B(new_n531), .C1(new_n922), .C2(new_n923), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G211gat), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(KEYINPUT125), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n940), .A2(new_n945), .A3(new_n941), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n927), .A2(new_n228), .A3(new_n531), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(G1354gat));
  AOI21_X1  g747(.A(G218gat), .B1(new_n927), .B2(new_n585), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT126), .Z(new_n950));
  NOR2_X1   g749(.A1(new_n924), .A2(KEYINPUT127), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n229), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n584), .B1(new_n924), .B2(KEYINPUT127), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1355gat));
endmodule


