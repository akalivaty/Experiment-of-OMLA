//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  OR2_X1    g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT91), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n208), .A2(KEYINPUT91), .ZN(new_n211));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n212), .A2(KEYINPUT92), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(new_n212), .B2(KEYINPUT92), .ZN(new_n216));
  OAI221_X1 g015(.A(new_n207), .B1(new_n210), .B2(new_n211), .C1(new_n213), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n208), .A2(new_n207), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(KEYINPUT94), .ZN(new_n219));
  INV_X1    g018(.A(G64gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G57gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT93), .B(G57gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(new_n220), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(KEYINPUT94), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n219), .A2(new_n215), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n206), .B1(new_n227), .B2(KEYINPUT21), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G127gat), .B(G155gat), .Z(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT20), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n230), .B(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n227), .A2(KEYINPUT21), .ZN(new_n234));
  NAND2_X1  g033(.A1(G231gat), .A2(G233gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(G183gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G211gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n234), .B(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT15), .ZN(new_n243));
  OR2_X1    g042(.A1(G43gat), .A2(G50gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(G43gat), .A2(G50gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT86), .B(G43gat), .Z(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT87), .B(G50gat), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n247), .A2(G50gat), .B1(new_n248), .B2(G43gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n249), .B2(new_n243), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NOR3_X1   g051(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n253));
  INV_X1    g052(.A(G29gat), .ZN(new_n254));
  INV_X1    g053(.A(G36gat), .ZN(new_n255));
  OAI22_X1  g054(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n246), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n256), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n260), .A2(KEYINPUT17), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(KEYINPUT17), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n263));
  NAND2_X1  g062(.A1(G85gat), .A2(G92gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G99gat), .ZN(new_n266));
  INV_X1    g065(.A(G106gat), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT8), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G99gat), .B(G106gat), .ZN(new_n269));
  OAI221_X1 g068(.A(new_n268), .B1(G85gat), .B2(G92gat), .C1(new_n269), .C2(KEYINPUT98), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(KEYINPUT98), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n271), .B(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n261), .A2(new_n262), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n271), .B(new_n272), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(new_n257), .A3(new_n259), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT99), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n278), .B1(new_n277), .B2(new_n279), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G190gat), .B(G218gat), .Z(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(G162gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT96), .B(G134gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n283), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n289), .B(new_n275), .C1(new_n280), .C2(new_n281), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n284), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n288), .B1(new_n284), .B2(new_n290), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n242), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n226), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n276), .A2(new_n227), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT10), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n276), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G230gat), .ZN(new_n302));
  INV_X1    g101(.A(G233gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n296), .A2(new_n297), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n304), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G176gat), .B(G204gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT100), .ZN(new_n311));
  XNOR2_X1  g110(.A(G120gat), .B(G148gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n314), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n295), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT80), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n322), .B(G57gat), .Z(new_n323));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324));
  INV_X1    g123(.A(G85gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n323), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  INV_X1    g128(.A(G141gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT74), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G141gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT75), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT74), .B(G141gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n329), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(G141gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G155gat), .ZN(new_n341));
  INV_X1    g140(.A(G162gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n349));
  INV_X1    g148(.A(G120gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(G113gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(G113gat), .ZN(new_n352));
  INV_X1    g151(.A(G113gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  OR2_X1    g154(.A1(G127gat), .A2(G134gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(G127gat), .A2(G134gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT1), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n353), .A2(G120gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n352), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n330), .A2(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n339), .A2(new_n366), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n345), .B(new_n343), .C1(new_n367), .C2(new_n344), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT69), .B1(new_n359), .B2(new_n364), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(new_n361), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(new_n356), .A3(new_n357), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n358), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT69), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n368), .B1(new_n340), .B2(new_n347), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n376), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n380), .A2(new_n385), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n348), .A2(new_n369), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT3), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n365), .B1(new_n380), .B2(new_n385), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT76), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n383), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n339), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n332), .A2(G141gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n330), .A2(KEYINPUT74), .ZN(new_n398));
  OAI21_X1  g197(.A(G148gat), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n396), .B1(new_n399), .B2(new_n336), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n346), .B1(new_n400), .B2(new_n335), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n387), .B1(new_n401), .B2(new_n368), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(KEYINPUT77), .A3(new_n370), .ZN(new_n403));
  INV_X1    g202(.A(new_n382), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n391), .A2(new_n405), .A3(new_n387), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n395), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n394), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n379), .A2(new_n380), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n371), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n413), .A2(new_n414), .A3(new_n382), .A4(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n328), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT38), .ZN(new_n425));
  INV_X1    g224(.A(G211gat), .ZN(new_n426));
  INV_X1    g225(.A(G218gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(KEYINPUT22), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT73), .B(G197gat), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(G204gat), .B2(new_n430), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n430), .A2(G204gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G211gat), .B(G218gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n434), .A3(new_n432), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT28), .ZN(new_n443));
  INV_X1    g242(.A(G190gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n444), .B1(new_n440), .B2(new_n441), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(KEYINPUT28), .ZN(new_n449));
  NAND2_X1  g248(.A1(G169gat), .A2(G176gat), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT64), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455));
  NOR2_X1   g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT26), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n457), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n454), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n449), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT23), .ZN(new_n463));
  INV_X1    g262(.A(G169gat), .ZN(new_n464));
  INV_X1    g263(.A(G176gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT25), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n468), .A2(new_n454), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(G183gat), .A2(G190gat), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n447), .B2(KEYINPUT24), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(KEYINPUT24), .B2(new_n447), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n468), .A2(new_n454), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n446), .A2(KEYINPUT65), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(G183gat), .A3(G190gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT24), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT66), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT24), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n476), .A2(new_n478), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n475), .B1(new_n472), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n462), .B(new_n474), .C1(new_n484), .C2(new_n469), .ZN(new_n485));
  AND2_X1   g284(.A1(G226gat), .A2(G233gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT29), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n486), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n439), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n468), .A2(new_n454), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(new_n472), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n494), .A2(KEYINPUT25), .B1(new_n473), .B2(new_n470), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT29), .B1(new_n495), .B2(new_n462), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n438), .B(new_n487), .C1(new_n496), .C2(new_n486), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(G8gat), .B(G36gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(G64gat), .B(G92gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n498), .A2(KEYINPUT37), .ZN(new_n504));
  INV_X1    g303(.A(new_n501), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n498), .B2(KEYINPUT37), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n425), .A2(new_n503), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n504), .A2(new_n506), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n425), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT84), .ZN(new_n510));
  INV_X1    g309(.A(new_n383), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n413), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n407), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT78), .B1(new_n407), .B2(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n419), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n510), .B1(new_n516), .B2(new_n328), .ZN(new_n517));
  AOI211_X1 g316(.A(KEYINPUT84), .B(new_n327), .C1(new_n515), .C2(new_n419), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n327), .A3(new_n419), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT81), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n515), .A2(KEYINPUT81), .A3(new_n327), .A4(new_n419), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n422), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n424), .B(new_n509), .C1(new_n519), .C2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT39), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n403), .A2(new_n406), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n382), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n417), .A2(new_n371), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n415), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(new_n390), .B2(new_n394), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n528), .B1(new_n531), .B2(new_n382), .ZN(new_n532));
  INV_X1    g331(.A(new_n394), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT76), .B1(new_n392), .B2(new_n393), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n418), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(new_n526), .A3(new_n404), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(new_n536), .A3(new_n327), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT83), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT40), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n505), .B1(new_n491), .B2(new_n497), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n502), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n498), .A2(KEYINPUT30), .A3(new_n501), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n538), .A2(new_n539), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n532), .A2(new_n536), .A3(new_n327), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT85), .B1(new_n519), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G78gat), .B(G106gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n386), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n439), .B1(new_n552), .B2(KEYINPUT29), .ZN(new_n553));
  INV_X1    g352(.A(G50gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT29), .B1(new_n436), .B2(new_n437), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n391), .B1(new_n555), .B2(KEYINPUT3), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n437), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n434), .B1(new_n431), .B2(new_n432), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n489), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n380), .B1(new_n560), .B2(new_n385), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n438), .B1(new_n386), .B2(new_n489), .ZN(new_n562));
  OAI21_X1  g361(.A(G50gat), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT31), .B(G22gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(G228gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n557), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n557), .B2(new_n563), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n551), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n557), .A2(new_n563), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n566), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n550), .A3(new_n568), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n421), .A2(KEYINPUT84), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n516), .A2(new_n510), .A3(new_n328), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OR3_X1    g377(.A1(new_n502), .A2(new_n542), .A3(new_n541), .ZN(new_n579));
  INV_X1    g378(.A(new_n544), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n579), .A2(new_n547), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT85), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n578), .A2(new_n581), .A3(new_n582), .A4(new_n540), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n525), .A2(new_n549), .A3(new_n575), .A4(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n495), .A2(new_n373), .A3(new_n378), .A4(new_n462), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n485), .A2(new_n379), .ZN(new_n586));
  INV_X1    g385(.A(G227gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(new_n303), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n589), .A2(KEYINPUT32), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(new_n586), .ZN(new_n592));
  INV_X1    g391(.A(new_n588), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI211_X1 g393(.A(KEYINPUT34), .B(new_n588), .C1(new_n585), .C2(new_n586), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n590), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n485), .A2(new_n379), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n485), .A2(new_n379), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT34), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n592), .A2(new_n591), .A3(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n589), .A2(KEYINPUT32), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n589), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT70), .B(G71gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n266), .ZN(new_n607));
  XNOR2_X1  g406(.A(G15gat), .B(G43gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n596), .A2(new_n603), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n610), .B1(new_n596), .B2(new_n603), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT71), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n611), .B2(new_n612), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n602), .B1(new_n600), .B2(new_n601), .ZN(new_n621));
  OAI22_X1  g420(.A1(new_n620), .A2(new_n621), .B1(new_n605), .B2(new_n609), .ZN(new_n622));
  INV_X1    g421(.A(new_n618), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n596), .A2(new_n603), .A3(new_n610), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n625), .A3(KEYINPUT36), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n616), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT82), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n421), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n516), .A2(KEYINPUT82), .A3(new_n328), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n424), .B1(new_n632), .B2(new_n524), .ZN(new_n633));
  INV_X1    g432(.A(new_n545), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n575), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n628), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n619), .A2(new_n625), .A3(new_n575), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n633), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT35), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n424), .B1(new_n519), .B2(new_n524), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT35), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n575), .A3(new_n613), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n584), .A2(new_n637), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n206), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n261), .A2(new_n648), .A3(new_n262), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n257), .A2(new_n206), .A3(new_n259), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT88), .ZN(new_n651));
  NAND2_X1  g450(.A1(G229gat), .A2(G233gat), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT89), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT18), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT18), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n260), .A2(new_n648), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n651), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n652), .B(KEYINPUT13), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664));
  INV_X1    g463(.A(G197gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT11), .B(G169gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT12), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n656), .A2(new_n658), .A3(new_n662), .A4(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n320), .B1(new_n647), .B2(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n522), .A2(new_n422), .A3(new_n523), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT82), .B1(new_n516), .B2(new_n328), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n629), .B(new_n327), .C1(new_n515), .C2(new_n419), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n423), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n636), .B1(new_n680), .B2(new_n545), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n584), .A3(new_n627), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT6), .B1(new_n520), .B2(new_n521), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n683), .A2(new_n630), .A3(new_n523), .A4(new_n631), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n545), .B(new_n638), .C1(new_n684), .C2(new_n424), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n646), .B1(new_n685), .B2(new_n643), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(KEYINPUT90), .A3(new_n673), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n319), .B1(new_n675), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n680), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g490(.A(KEYINPUT16), .B(G8gat), .Z(new_n692));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n545), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(KEYINPUT42), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n545), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(G8gat), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n694), .B1(new_n693), .B2(new_n697), .ZN(G1325gat));
  AOI21_X1  g497(.A(G15gat), .B1(new_n689), .B2(new_n613), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(KEYINPUT101), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(KEYINPUT101), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n627), .B(KEYINPUT102), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n689), .A2(G15gat), .A3(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n700), .A2(new_n701), .A3(new_n704), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n636), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(new_n318), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n241), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n294), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n675), .B2(new_n688), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n254), .A3(new_n680), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT45), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n673), .ZN(new_n715));
  INV_X1    g514(.A(new_n294), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n682), .B2(new_n686), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT103), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n720), .B(KEYINPUT44), .C1(new_n647), .C2(new_n716), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n641), .A2(KEYINPUT104), .A3(new_n646), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT104), .B1(new_n641), .B2(new_n646), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n682), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n293), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n726), .A2(KEYINPUT105), .A3(new_n291), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT105), .B1(new_n726), .B2(new_n291), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n715), .B1(new_n722), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n633), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n714), .A2(new_n735), .ZN(G1328gat));
  OAI21_X1  g535(.A(G36gat), .B1(new_n734), .B2(new_n634), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n712), .A2(new_n255), .A3(new_n545), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(G1329gat));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n613), .A2(new_n247), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n712), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n247), .B1(new_n733), .B2(new_n703), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI211_X1 g547(.A(KEYINPUT106), .B(new_n247), .C1(new_n733), .C2(new_n703), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n743), .B1(new_n712), .B2(new_n744), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n719), .A2(new_n721), .B1(new_n725), .B2(new_n731), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n627), .A3(new_n715), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n753), .B2(new_n247), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT107), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n756), .B(new_n751), .C1(new_n753), .C2(new_n247), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n750), .A2(new_n758), .ZN(G1330gat));
  INV_X1    g558(.A(new_n248), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n712), .B2(new_n636), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(KEYINPUT48), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n733), .A2(new_n636), .A3(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n762), .A2(KEYINPUT48), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1331gat));
  AND4_X1   g566(.A1(new_n674), .A2(new_n725), .A3(new_n295), .A4(new_n709), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n680), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(new_n222), .ZN(G1332gat));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n545), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT49), .B(G64gat), .Z(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(G1333gat));
  NAND2_X1  g573(.A1(new_n768), .A2(new_n703), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n614), .A2(G71gat), .ZN(new_n776));
  AOI22_X1  g575(.A1(new_n775), .A2(G71gat), .B1(new_n768), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n768), .A2(new_n636), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g580(.A1(new_n716), .A2(new_n673), .A3(new_n241), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n725), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT51), .Z(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(new_n325), .A3(new_n680), .A4(new_n709), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n674), .A2(new_n242), .A3(new_n709), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT110), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n752), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n789), .A3(new_n680), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G85gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n788), .B2(new_n680), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n785), .B1(new_n791), .B2(new_n792), .ZN(G1336gat));
  NOR3_X1   g592(.A1(new_n318), .A2(G92gat), .A3(new_n634), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n788), .A2(new_n545), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G92gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n725), .A2(KEYINPUT112), .A3(new_n782), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n799), .B2(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g599(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n725), .A2(new_n782), .B1(KEYINPUT112), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n796), .A2(G92gat), .B1(new_n803), .B2(new_n794), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n798), .B1(new_n804), .B2(new_n805), .ZN(G1337gat));
  INV_X1    g605(.A(new_n784), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n709), .A2(new_n266), .A3(new_n613), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n752), .A2(new_n702), .A3(new_n787), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n807), .A2(new_n808), .B1(new_n266), .B2(new_n809), .ZN(G1338gat));
  XOR2_X1   g609(.A(KEYINPUT114), .B(G106gat), .Z(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n788), .B2(new_n636), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n709), .A2(new_n267), .A3(new_n636), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n800), .A2(new_n802), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT53), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n788), .B2(new_n636), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n752), .A2(KEYINPUT115), .A3(new_n575), .A4(new_n787), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n807), .B2(new_n813), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n815), .B1(new_n819), .B2(new_n821), .ZN(G1339gat));
  NOR2_X1   g621(.A1(new_n319), .A2(new_n673), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n301), .A2(new_n305), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n304), .B1(new_n299), .B2(new_n300), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n314), .B1(new_n306), .B2(KEYINPUT54), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n313), .B1(new_n826), .B2(new_n825), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT116), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n827), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n315), .B1(new_n833), .B2(KEYINPUT55), .ZN(new_n834));
  INV_X1    g633(.A(new_n827), .ZN(new_n835));
  INV_X1    g634(.A(new_n832), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n831), .A2(KEYINPUT116), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n673), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n660), .A2(new_n661), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n652), .B1(new_n649), .B2(new_n651), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n668), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n672), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(new_n318), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n730), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n834), .A2(new_n840), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n672), .A2(KEYINPUT117), .A3(new_n844), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n849), .A2(new_n729), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n823), .B1(new_n854), .B2(new_n242), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n633), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n645), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n674), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n855), .A2(new_n633), .A3(new_n638), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n634), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n673), .A2(new_n353), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(G1340gat));
  OAI21_X1  g661(.A(G120gat), .B1(new_n857), .B2(new_n318), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n709), .A2(new_n350), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n860), .B2(new_n864), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n857), .B2(new_n242), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n242), .A2(G127gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT118), .ZN(G1342gat));
  NAND2_X1  g668(.A1(new_n294), .A2(new_n634), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT119), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(G134gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n859), .A2(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n873), .A2(KEYINPUT120), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n857), .B2(new_n716), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT121), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n874), .A2(KEYINPUT56), .A3(new_n875), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  OR3_X1    g681(.A1(new_n855), .A2(KEYINPUT57), .A3(new_n575), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n834), .A2(new_n852), .A3(new_n840), .A4(new_n850), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n730), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n294), .B1(new_n841), .B2(new_n846), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n823), .B1(new_n887), .B2(new_n242), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT57), .B1(new_n888), .B2(new_n575), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n628), .A2(new_n633), .A3(new_n545), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n337), .B1(new_n891), .B2(new_n674), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n703), .A2(new_n575), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n856), .A2(new_n634), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n330), .A3(new_n673), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n896), .B(new_n897), .ZN(G1344gat));
  NAND3_X1  g697(.A1(new_n894), .A2(new_n329), .A3(new_n709), .ZN(new_n899));
  INV_X1    g698(.A(new_n891), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT59), .B(new_n329), .C1(new_n900), .C2(new_n709), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n884), .A2(new_n716), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n242), .B1(new_n903), .B2(new_n886), .ZN(new_n904));
  INV_X1    g703(.A(new_n823), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n575), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n906), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT123), .B1(new_n906), .B2(KEYINPUT57), .ZN(new_n908));
  INV_X1    g707(.A(new_n855), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(KEYINPUT57), .A3(new_n636), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n709), .A3(new_n890), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n902), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n899), .B1(new_n901), .B2(new_n913), .ZN(G1345gat));
  AOI21_X1  g713(.A(G155gat), .B1(new_n894), .B2(new_n241), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n242), .A2(new_n341), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n900), .B2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n891), .B2(new_n730), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n871), .A2(G162gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n856), .A2(new_n893), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1347gat));
  AOI21_X1  g720(.A(new_n729), .B1(new_n841), .B2(new_n846), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n242), .B1(new_n885), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n680), .B1(new_n923), .B2(new_n905), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n545), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT124), .B(new_n680), .C1(new_n923), .C2(new_n905), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n926), .A2(new_n638), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n464), .A3(new_n673), .ZN(new_n929));
  AND4_X1   g728(.A1(new_n545), .A2(new_n924), .A3(new_n575), .A4(new_n613), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(new_n673), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n929), .B1(new_n464), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT125), .ZN(G1348gat));
  AOI21_X1  g732(.A(G176gat), .B1(new_n928), .B2(new_n709), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n318), .A2(new_n465), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n930), .B2(new_n935), .ZN(G1349gat));
  NAND2_X1  g735(.A1(new_n930), .A2(new_n241), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(G183gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n241), .A2(new_n442), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT126), .B1(new_n928), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT124), .B1(new_n855), .B2(new_n680), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n925), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n942), .A2(new_n943), .A3(new_n545), .A4(new_n639), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n939), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n938), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n949), .B(new_n938), .C1(new_n941), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n928), .A2(new_n444), .A3(new_n729), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n930), .A2(new_n294), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G190gat), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n943), .A3(new_n545), .A4(new_n893), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT127), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n665), .A3(new_n673), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n703), .A2(new_n680), .A3(new_n634), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n911), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(G197gat), .B1(new_n962), .B2(new_n674), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(G1352gat));
  NAND3_X1  g763(.A1(new_n911), .A2(new_n709), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n318), .A2(G204gat), .ZN(new_n967));
  OR3_X1    g766(.A1(new_n958), .A2(KEYINPUT62), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT62), .B1(new_n958), .B2(new_n967), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n959), .A2(new_n426), .A3(new_n241), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n911), .A2(new_n241), .A3(new_n961), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n972), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(G211gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(G1354gat));
  NOR3_X1   g774(.A1(new_n962), .A2(new_n427), .A3(new_n716), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n729), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(new_n427), .ZN(G1355gat));
endmodule


