//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n445, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n471), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n475), .A2(new_n474), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n483));
  INV_X1    g058(.A(new_n470), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n472), .A3(new_n485), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n470), .C2(G112), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  AND3_X1   g069(.A1(new_n472), .A2(G102), .A3(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(G126), .B1(new_n475), .B2(new_n474), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n464), .A2(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G138), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n478), .A2(KEYINPUT4), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT71), .B1(new_n515), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT5), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n516), .A2(new_n519), .B1(new_n515), .B2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(new_n511), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(G62), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(KEYINPUT72), .A3(G62), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n528), .A2(KEYINPUT73), .A3(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT73), .B1(new_n528), .B2(G651), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n514), .B(new_n522), .C1(new_n529), .C2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND2_X1  g107(.A1(new_n521), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n513), .A2(G51), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n533), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AOI22_X1  g114(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n507), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n520), .A2(new_n511), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n542), .A2(new_n543), .B1(new_n544), .B2(new_n512), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n541), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n507), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n542), .A2(new_n549), .B1(new_n550), .B2(new_n512), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT75), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n557), .B(new_n548), .C1(new_n553), .C2(new_n554), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT76), .Z(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND3_X1  g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT8), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n564), .A2(KEYINPUT8), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT77), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n520), .B2(G65), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n507), .B1(new_n542), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n508), .A2(new_n510), .A3(G53), .A4(G543), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n574), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  NAND2_X1  g161(.A1(new_n521), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n513), .A2(G49), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n507), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  INV_X1    g168(.A(G48), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n542), .A2(new_n593), .B1(new_n594), .B2(new_n512), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n507), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(KEYINPUT80), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(KEYINPUT80), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n600), .A2(new_n601), .B1(G47), .B2(new_n513), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT81), .B(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n521), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT84), .Z(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n521), .A2(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT10), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n611), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n513), .A2(G54), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n584), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n584), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n490), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n487), .A2(G123), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n631));
  OR3_X1    g206(.A1(new_n470), .A2(new_n631), .A3(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n470), .B2(G111), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n632), .A2(new_n633), .A3(G2104), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n629), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT86), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2100), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n650), .A2(KEYINPUT88), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(KEYINPUT88), .ZN(new_n652));
  OAI22_X1  g227(.A1(new_n651), .A2(new_n652), .B1(new_n645), .B2(new_n648), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2443), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n661), .A3(new_n659), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT89), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n671), .A3(KEYINPUT17), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT91), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n680), .A2(new_n681), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n683), .A2(new_n685), .A3(new_n688), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n687), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT93), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT92), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n693), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  INV_X1    g274(.A(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(G229));
  XNOR2_X1  g277(.A(KEYINPUT95), .B(G16), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G24), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n605), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT98), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G23), .ZN(new_n712));
  INV_X1    g287(.A(G288), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT33), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1976), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(G6), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n596), .B2(new_n711), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(KEYINPUT96), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(KEYINPUT96), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT32), .B(G1981), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n703), .A2(G22), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G303), .B2(new_n704), .ZN(new_n726));
  INV_X1    g301(.A(G1971), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n716), .A2(new_n724), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT97), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n710), .B1(new_n734), .B2(KEYINPUT34), .ZN(new_n735));
  AND2_X1   g310(.A1(KEYINPUT94), .A2(G29), .ZN(new_n736));
  NOR2_X1   g311(.A1(KEYINPUT94), .A2(G29), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n487), .A2(G119), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n490), .A2(G131), .ZN(new_n742));
  OAI221_X1 g317(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n470), .C2(G107), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(new_n739), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT35), .B(G1991), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n746), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n732), .B2(new_n733), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n735), .A2(KEYINPUT36), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n730), .A2(new_n731), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n730), .A2(new_n731), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n753), .A2(KEYINPUT34), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n751), .A2(new_n755), .A3(new_n749), .A4(new_n709), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT31), .B(G11), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT100), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(new_n484), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n490), .A2(G139), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G29), .B2(G33), .ZN(new_n769));
  INV_X1    g344(.A(G2072), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT101), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n704), .A2(KEYINPUT23), .A3(G20), .ZN(new_n773));
  AOI21_X1  g348(.A(KEYINPUT23), .B1(new_n704), .B2(G20), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n773), .B(new_n774), .C1(G299), .C2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n769), .A2(new_n770), .ZN(new_n778));
  NOR2_X1   g353(.A1(G5), .A2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G171), .B2(G16), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n490), .A2(G141), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n487), .A2(G129), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT102), .Z(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT26), .Z(new_n786));
  NAND4_X1  g361(.A1(new_n781), .A2(new_n782), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G29), .B2(G32), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT27), .B(G1996), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n778), .B1(G1961), .B2(new_n780), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n772), .A2(new_n777), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n739), .A2(G35), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G162), .B2(new_n739), .ZN(new_n795));
  MUX2_X1   g370(.A(new_n794), .B(new_n795), .S(KEYINPUT103), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT29), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n797), .A2(KEYINPUT104), .A3(G2090), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G4), .B2(G16), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n800), .A2(G4), .A3(G16), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n801), .B(new_n802), .C1(new_n616), .C2(new_n711), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1348), .ZN(new_n804));
  OAI221_X1 g379(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n470), .C2(G116), .ZN(new_n805));
  INV_X1    g380(.A(G128), .ZN(new_n806));
  INV_X1    g381(.A(G140), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n805), .B1(new_n486), .B2(new_n806), .C1(new_n807), .C2(new_n489), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n739), .A2(G26), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n808), .A2(G29), .B1(KEYINPUT28), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(KEYINPUT28), .B2(new_n809), .ZN(new_n811));
  INV_X1    g386(.A(G2067), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT24), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(G34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(G34), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n739), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G160), .ZN(new_n818));
  INV_X1    g393(.A(G29), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2084), .ZN(new_n821));
  INV_X1    g396(.A(new_n636), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT30), .B(G28), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n822), .A2(new_n738), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n780), .A2(G1961), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n711), .A2(G21), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G168), .B2(new_n711), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1966), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n739), .A2(G27), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G164), .B2(new_n739), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2078), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n826), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n804), .A2(new_n813), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n703), .A2(G19), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n559), .B2(new_n703), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(G1341), .Z(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n837), .C1(G2090), .C2(new_n797), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n790), .A2(new_n791), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT104), .B1(new_n797), .B2(G2090), .ZN(new_n840));
  NOR4_X1   g415(.A1(new_n799), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n752), .A2(new_n758), .A3(new_n759), .A4(new_n841), .ZN(G150));
  INV_X1    g417(.A(G150), .ZN(G311));
  AOI22_X1  g418(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n507), .ZN(new_n845));
  INV_X1    g420(.A(G93), .ZN(new_n846));
  INV_X1    g421(.A(G55), .ZN(new_n847));
  OAI22_X1  g422(.A1(new_n542), .A2(new_n846), .B1(new_n847), .B2(new_n512), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NOR2_X1   g427(.A1(new_n616), .A2(new_n623), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n559), .A2(new_n850), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n555), .A2(new_n849), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n855), .B(new_n858), .Z(new_n859));
  OAI21_X1  g434(.A(new_n852), .B1(new_n859), .B2(G860), .ZN(G145));
  OAI221_X1 g435(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n470), .C2(G118), .ZN(new_n861));
  INV_X1    g436(.A(G142), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n489), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G130), .B2(new_n487), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(new_n493), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n822), .ZN(new_n866));
  INV_X1    g441(.A(new_n640), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n808), .A2(G164), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n808), .A2(G164), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n787), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n808), .A2(G164), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n808), .A2(G164), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n788), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n867), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n873), .A3(new_n867), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n745), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n744), .B1(new_n878), .B2(new_n874), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n766), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n879), .A3(new_n766), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n866), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(new_n866), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n884), .A2(new_n880), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(G160), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n882), .A3(new_n866), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n884), .B2(new_n880), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n818), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g468(.A1(new_n849), .A2(G868), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n713), .B(new_n596), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(G303), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n605), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT42), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n858), .B(new_n625), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n616), .B(new_n584), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n899), .A2(new_n905), .A3(new_n907), .A4(new_n901), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI211_X1 g486(.A(KEYINPUT105), .B(new_n894), .C1(new_n911), .C2(G868), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n913));
  INV_X1    g488(.A(new_n910), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n899), .A2(new_n901), .B1(new_n905), .B2(new_n907), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n894), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n912), .A2(new_n918), .ZN(G295));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n917), .ZN(G331));
  XNOR2_X1  g495(.A(new_n616), .B(G299), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT41), .ZN(new_n922));
  OAI21_X1  g497(.A(G286), .B1(G171), .B2(KEYINPUT106), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n856), .B2(new_n857), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n849), .B1(new_n556), .B2(new_n558), .ZN(new_n925));
  INV_X1    g500(.A(new_n857), .ZN(new_n926));
  INV_X1    g501(.A(new_n923), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n929));
  NOR2_X1   g504(.A1(G301), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n924), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n856), .A2(new_n857), .A3(new_n923), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n925), .B2(new_n926), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n922), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n930), .A3(new_n934), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n904), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n898), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n906), .A2(new_n937), .A3(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n921), .B1(new_n932), .B2(new_n935), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n897), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n888), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n940), .A2(new_n946), .A3(new_n888), .A4(new_n943), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(G397));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n505), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G160), .A2(G40), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n808), .B(G2067), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n959), .B2(new_n787), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n961));
  INV_X1    g536(.A(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(G1996), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n958), .A2(KEYINPUT46), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT127), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT47), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n787), .B(new_n964), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(new_n959), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n744), .A2(new_n747), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(G2067), .B2(new_n808), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n958), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n605), .A2(new_n700), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(new_n962), .ZN(new_n977));
  XOR2_X1   g552(.A(new_n977), .B(KEYINPUT48), .Z(new_n978));
  INV_X1    g553(.A(new_n971), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n745), .A2(new_n748), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n979), .A2(new_n980), .A3(new_n972), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n978), .B1(new_n962), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n968), .A2(new_n975), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT63), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(KEYINPUT63), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n988));
  INV_X1    g563(.A(G40), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n471), .A2(new_n480), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT4), .B1(new_n478), .B2(new_n503), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n466), .A2(new_n470), .A3(new_n500), .A4(G138), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1384), .B1(new_n993), .B2(new_n499), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n988), .A2(new_n990), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(G2084), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n955), .B(G1384), .C1(new_n993), .C2(new_n499), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n990), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1002));
  OR3_X1    g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1966), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n998), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n957), .B1(new_n955), .B2(new_n954), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n727), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n994), .A2(new_n995), .ZN(new_n1012));
  AOI211_X1 g587(.A(KEYINPUT50), .B(G1384), .C1(new_n993), .C2(new_n499), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n957), .ZN(new_n1014));
  INV_X1    g589(.A(G2090), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1006), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1002), .A2(new_n999), .ZN(new_n1022));
  OAI22_X1  g597(.A1(G1971), .A2(new_n1022), .B1(new_n997), .B2(G2090), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(G8), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1020), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n1018), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n596), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT108), .B(G1981), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n592), .A2(new_n595), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1030), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n596), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(KEYINPUT49), .C1(new_n1028), .C2(new_n596), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n994), .A2(new_n990), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1032), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G288), .A2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1037), .A2(KEYINPUT107), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G288), .A2(new_n1040), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1039), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1007), .A2(new_n1021), .A3(new_n1026), .A4(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n985), .B(new_n987), .C1(new_n1049), .C2(G286), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1021), .A2(new_n1048), .A3(new_n1026), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(G168), .A3(new_n1007), .A4(new_n986), .ZN(new_n1052));
  XOR2_X1   g627(.A(new_n1037), .B(KEYINPUT109), .Z(new_n1053));
  NOR3_X1   g628(.A1(new_n1039), .A2(G1976), .A3(G288), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1031), .B(KEYINPUT110), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1050), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1048), .B(new_n1017), .C1(new_n1020), .C2(new_n1019), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1059), .A2(G2078), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1003), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1059), .B1(new_n1010), .B2(G2078), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT123), .B(G1961), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n997), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G301), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G168), .A2(new_n1006), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1067), .B(new_n1069), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n1071), .A2(G1966), .B1(G2084), .B2(new_n997), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT51), .B(G8), .C1(new_n1072), .C2(G286), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1070), .A2(new_n1073), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1074), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1051), .B1(new_n1077), .B2(KEYINPUT62), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1057), .B(new_n1058), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n956), .A2(new_n990), .A3(new_n1009), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT116), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1008), .A2(new_n1083), .A3(new_n1009), .A4(new_n1080), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n574), .A2(new_n577), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n584), .B2(KEYINPUT57), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n582), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n1093));
  NOR4_X1   g668(.A1(new_n1092), .A2(KEYINPUT115), .A3(new_n1093), .A4(new_n574), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1088), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT113), .B1(new_n997), .B2(new_n776), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n997), .A2(KEYINPUT113), .A3(new_n776), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1085), .B(new_n1095), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1085), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1095), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1014), .B2(G1956), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n997), .A2(KEYINPUT113), .A3(new_n776), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1105), .A2(new_n1106), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT117), .A3(new_n1095), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1100), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1002), .A2(G1996), .A3(new_n999), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT118), .B(G1341), .Z(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT58), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1036), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1112), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n956), .A2(new_n964), .A3(new_n990), .A4(new_n1009), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(KEYINPUT119), .A3(new_n1116), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n559), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1123), .A2(KEYINPUT59), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1118), .A2(KEYINPUT120), .A3(new_n559), .A4(new_n1120), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(KEYINPUT59), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1110), .B1(new_n1107), .B2(new_n1095), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1123), .A2(new_n1126), .B1(new_n1127), .B2(new_n1103), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1111), .A2(new_n1124), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1111), .A2(new_n1128), .A3(new_n1131), .A4(new_n1124), .ZN(new_n1132));
  INV_X1    g707(.A(G1348), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1036), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n997), .A2(new_n1133), .B1(new_n812), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n617), .B1(new_n1135), .B2(KEYINPUT60), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT122), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(KEYINPUT60), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1137), .B(new_n1138), .Z(new_n1139));
  NAND3_X1  g714(.A1(new_n1130), .A2(new_n1132), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1103), .B1(new_n616), .B2(new_n1135), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n1100), .A3(new_n1108), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1061), .A2(new_n1065), .A3(G301), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n1145));
  OAI21_X1  g720(.A(G40), .B1(new_n480), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n999), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n471), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1060), .B1(new_n480), .B2(new_n1145), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n956), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1062), .A2(new_n1064), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(G171), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1152), .B1(new_n1151), .B2(G171), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1144), .B(KEYINPUT54), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1151), .A2(G171), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT125), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1161), .B2(new_n1153), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(KEYINPUT126), .A3(new_n1144), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1151), .A2(G171), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1159), .B1(new_n1066), .B2(new_n1165), .ZN(new_n1166));
  AND4_X1   g741(.A1(new_n1077), .A2(new_n1164), .A3(new_n1051), .A4(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1079), .B1(new_n1143), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n981), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(G1986), .B2(G290), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n962), .B1(new_n1170), .B2(new_n976), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n983), .B1(new_n1168), .B2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g747(.A1(G401), .A2(new_n462), .ZN(new_n1174));
  NOR2_X1   g748(.A1(G229), .A2(G227), .ZN(new_n1175));
  NAND4_X1  g749(.A1(new_n948), .A2(new_n1174), .A3(new_n892), .A4(new_n1175), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


