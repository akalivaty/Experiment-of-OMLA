

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740;

  INV_X1 U375 ( .A(G953), .ZN(n731) );
  NOR2_X1 U376 ( .A1(n574), .A2(n573), .ZN(n668) );
  XNOR2_X1 U377 ( .A(n517), .B(n516), .ZN(n737) );
  NAND2_X2 U378 ( .A1(n595), .A2(n609), .ZN(n428) );
  INV_X2 U379 ( .A(n539), .ZN(n617) );
  AND2_X1 U380 ( .A1(n383), .A2(n414), .ZN(n727) );
  NOR2_X4 U381 ( .A1(n617), .A2(n618), .ZN(n615) );
  NOR2_X1 U382 ( .A1(n355), .A2(n359), .ZN(n365) );
  INV_X1 U383 ( .A(G116), .ZN(n389) );
  XNOR2_X1 U384 ( .A(n429), .B(n489), .ZN(n514) );
  NOR2_X1 U385 ( .A1(n426), .A2(n584), .ZN(n520) );
  XNOR2_X1 U386 ( .A(n560), .B(n398), .ZN(n584) );
  NAND2_X2 U387 ( .A1(n365), .A2(n419), .ZN(n560) );
  XNOR2_X1 U388 ( .A(n397), .B(n510), .ZN(n647) );
  XNOR2_X1 U389 ( .A(n370), .B(n500), .ZN(n711) );
  XNOR2_X1 U390 ( .A(n725), .B(G146), .ZN(n397) );
  XNOR2_X1 U391 ( .A(n380), .B(n466), .ZN(n725) );
  XNOR2_X1 U392 ( .A(n435), .B(n364), .ZN(n454) );
  XNOR2_X1 U393 ( .A(n396), .B(G128), .ZN(n447) );
  XNOR2_X1 U394 ( .A(n389), .B(G107), .ZN(n472) );
  XNOR2_X1 U395 ( .A(KEYINPUT71), .B(G110), .ZN(n473) );
  XNOR2_X1 U396 ( .A(G131), .B(KEYINPUT68), .ZN(n435) );
  BUF_X1 U397 ( .A(n596), .Z(n354) );
  XNOR2_X1 U398 ( .A(n363), .B(n544), .ZN(n596) );
  XNOR2_X2 U399 ( .A(n400), .B(n361), .ZN(n527) );
  NOR2_X1 U400 ( .A1(n706), .A2(n713), .ZN(n707) );
  NOR2_X1 U401 ( .A1(n700), .A2(n713), .ZN(n703) );
  XOR2_X1 U402 ( .A(G137), .B(G140), .Z(n491) );
  XNOR2_X1 U403 ( .A(n447), .B(n434), .ZN(n466) );
  INV_X1 U404 ( .A(KEYINPUT4), .ZN(n434) );
  NOR2_X1 U405 ( .A1(n560), .A2(n581), .ZN(n555) );
  OR2_X1 U406 ( .A1(G902), .A2(G237), .ZN(n485) );
  XNOR2_X1 U407 ( .A(G116), .B(G137), .ZN(n507) );
  XNOR2_X1 U408 ( .A(n506), .B(n418), .ZN(n417) );
  AND2_X1 U409 ( .A1(n505), .A2(G210), .ZN(n418) );
  XNOR2_X1 U410 ( .A(n454), .B(G134), .ZN(n380) );
  XNOR2_X1 U411 ( .A(G128), .B(KEYINPUT23), .ZN(n493) );
  XOR2_X1 U412 ( .A(G101), .B(G107), .Z(n433) );
  NOR2_X1 U413 ( .A1(n623), .A2(n399), .ZN(n624) );
  NOR2_X1 U414 ( .A1(n727), .A2(KEYINPUT2), .ZN(n413) );
  NOR2_X1 U415 ( .A1(n691), .A2(G902), .ZN(n442) );
  NOR2_X1 U416 ( .A1(n682), .A2(n415), .ZN(n414) );
  XNOR2_X1 U417 ( .A(n385), .B(n384), .ZN(n383) );
  INV_X1 U418 ( .A(n681), .ZN(n415) );
  INV_X1 U419 ( .A(KEYINPUT16), .ZN(n368) );
  XNOR2_X1 U420 ( .A(KEYINPUT3), .B(G119), .ZN(n469) );
  XOR2_X1 U421 ( .A(G101), .B(G113), .Z(n470) );
  XOR2_X1 U422 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n448) );
  XNOR2_X1 U423 ( .A(n449), .B(n391), .ZN(n390) );
  INV_X1 U424 ( .A(n447), .ZN(n391) );
  XNOR2_X1 U425 ( .A(G122), .B(G134), .ZN(n445) );
  XNOR2_X1 U426 ( .A(n382), .B(n381), .ZN(n589) );
  INV_X1 U427 ( .A(KEYINPUT39), .ZN(n381) );
  NOR2_X1 U428 ( .A1(n567), .A2(n605), .ZN(n382) );
  NAND2_X1 U429 ( .A1(n392), .A2(n431), .ZN(n430) );
  OR2_X1 U430 ( .A1(n647), .A2(n420), .ZN(n419) );
  NAND2_X1 U431 ( .A1(G472), .A2(n421), .ZN(n420) );
  XNOR2_X1 U432 ( .A(n453), .B(n394), .ZN(n530) );
  XNOR2_X1 U433 ( .A(n498), .B(n371), .ZN(n370) );
  INV_X1 U434 ( .A(KEYINPUT100), .ZN(n408) );
  NAND2_X1 U435 ( .A1(n576), .A2(n408), .ZN(n406) );
  INV_X1 U436 ( .A(KEYINPUT67), .ZN(n364) );
  XNOR2_X1 U437 ( .A(n465), .B(n379), .ZN(n490) );
  INV_X1 U438 ( .A(KEYINPUT10), .ZN(n379) );
  NOR2_X1 U439 ( .A1(n588), .A2(n587), .ZN(n387) );
  INV_X1 U440 ( .A(KEYINPUT48), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n490), .B(n491), .ZN(n724) );
  INV_X1 U442 ( .A(G143), .ZN(n396) );
  XOR2_X1 U443 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n446) );
  XNOR2_X1 U444 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U445 ( .A(KEYINPUT73), .B(KEYINPUT18), .Z(n478) );
  INV_X1 U446 ( .A(n618), .ZN(n431) );
  XNOR2_X1 U447 ( .A(n483), .B(KEYINPUT87), .ZN(n484) );
  INV_X1 U448 ( .A(G902), .ZN(n421) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n488) );
  XNOR2_X1 U450 ( .A(n417), .B(n416), .ZN(n509) );
  XNOR2_X1 U451 ( .A(n507), .B(KEYINPUT95), .ZN(n416) );
  XOR2_X1 U452 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n494) );
  XNOR2_X1 U453 ( .A(G119), .B(G110), .ZN(n496) );
  XNOR2_X1 U454 ( .A(n437), .B(n440), .ZN(n427) );
  XNOR2_X1 U455 ( .A(n439), .B(n438), .ZN(n440) );
  NOR2_X1 U456 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X1 U457 ( .A(n413), .B(n412), .ZN(n598) );
  INV_X1 U458 ( .A(KEYINPUT81), .ZN(n412) );
  AND2_X1 U459 ( .A1(n519), .A2(n424), .ZN(n625) );
  NOR2_X1 U460 ( .A1(n425), .A2(n560), .ZN(n424) );
  NOR2_X1 U461 ( .A1(n560), .A2(n559), .ZN(n561) );
  BUF_X1 U462 ( .A(n595), .Z(n375) );
  XNOR2_X1 U463 ( .A(n504), .B(n503), .ZN(n539) );
  NOR2_X1 U464 ( .A1(G902), .A2(n711), .ZN(n504) );
  INV_X1 U465 ( .A(KEYINPUT6), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n474), .B(n368), .ZN(n367) );
  XNOR2_X1 U467 ( .A(n390), .B(n388), .ZN(n452) );
  XNOR2_X1 U468 ( .A(n472), .B(n448), .ZN(n388) );
  NOR2_X1 U469 ( .A1(n604), .A2(n574), .ZN(n558) );
  AND2_X1 U470 ( .A1(n589), .A2(n669), .ZN(n565) );
  INV_X1 U471 ( .A(KEYINPUT32), .ZN(n516) );
  XNOR2_X1 U472 ( .A(n709), .B(n372), .ZN(n712) );
  AND2_X1 U473 ( .A1(n647), .A2(n422), .ZN(n355) );
  AND2_X1 U474 ( .A1(n487), .A2(n547), .ZN(n356) );
  XNOR2_X1 U475 ( .A(n568), .B(KEYINPUT75), .ZN(n357) );
  XOR2_X1 U476 ( .A(n454), .B(n490), .Z(n358) );
  XNOR2_X1 U477 ( .A(n393), .B(KEYINPUT101), .ZN(n607) );
  INV_X1 U478 ( .A(n607), .ZN(n392) );
  AND2_X1 U479 ( .A1(n422), .A2(G902), .ZN(n359) );
  AND2_X1 U480 ( .A1(n538), .A2(KEYINPUT100), .ZN(n360) );
  XOR2_X1 U481 ( .A(n523), .B(KEYINPUT74), .Z(n361) );
  INV_X1 U482 ( .A(G472), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n397), .B(n427), .ZN(n691) );
  XNOR2_X1 U484 ( .A(KEYINPUT106), .B(KEYINPUT62), .ZN(n362) );
  NOR2_X1 U485 ( .A1(n405), .A2(n403), .ZN(n410) );
  NAND2_X1 U486 ( .A1(n542), .A2(n543), .ZN(n363) );
  NAND2_X1 U487 ( .A1(n410), .A2(n423), .ZN(n374) );
  NAND2_X1 U488 ( .A1(n564), .A2(n366), .ZN(n567) );
  XNOR2_X1 U489 ( .A(n561), .B(KEYINPUT30), .ZN(n366) );
  NAND2_X1 U490 ( .A1(n667), .A2(n570), .ZN(n571) );
  NAND2_X1 U491 ( .A1(n569), .A2(n375), .ZN(n667) );
  AND2_X2 U492 ( .A1(n596), .A2(n727), .ZN(n643) );
  XNOR2_X1 U493 ( .A(n374), .B(KEYINPUT85), .ZN(n542) );
  XNOR2_X1 U494 ( .A(n475), .B(n367), .ZN(n476) );
  XNOR2_X1 U495 ( .A(n476), .B(n508), .ZN(n714) );
  NAND2_X1 U496 ( .A1(n369), .A2(n601), .ZN(n602) );
  XNOR2_X1 U497 ( .A(n600), .B(n599), .ZN(n369) );
  INV_X1 U498 ( .A(n605), .ZN(n395) );
  INV_X1 U499 ( .A(n724), .ZN(n371) );
  NOR2_X1 U500 ( .A1(n689), .A2(n713), .ZN(n690) );
  XNOR2_X1 U501 ( .A(n493), .B(n492), .ZN(n495) );
  INV_X1 U502 ( .A(n615), .ZN(n425) );
  XNOR2_X1 U503 ( .A(n711), .B(n710), .ZN(n372) );
  NAND2_X1 U504 ( .A1(n708), .A2(G478), .ZN(n704) );
  NOR2_X4 U505 ( .A1(n686), .A2(n644), .ZN(n708) );
  XNOR2_X1 U506 ( .A(n373), .B(n482), .ZN(n683) );
  XNOR2_X1 U507 ( .A(n714), .B(n481), .ZN(n373) );
  NAND2_X1 U508 ( .A1(n657), .A2(n674), .ZN(n537) );
  XNOR2_X2 U509 ( .A(n536), .B(KEYINPUT96), .ZN(n657) );
  NAND2_X1 U510 ( .A1(n404), .A2(n376), .ZN(n403) );
  INV_X1 U511 ( .A(n653), .ZN(n376) );
  NOR2_X2 U512 ( .A1(n541), .A2(n540), .ZN(n653) );
  XNOR2_X2 U513 ( .A(n377), .B(n484), .ZN(n595) );
  NAND2_X1 U514 ( .A1(n683), .A2(n644), .ZN(n377) );
  NAND2_X1 U515 ( .A1(n378), .A2(n579), .ZN(n580) );
  NAND2_X1 U516 ( .A1(n578), .A2(n577), .ZN(n378) );
  XNOR2_X2 U517 ( .A(n643), .B(KEYINPUT2), .ZN(n686) );
  XNOR2_X1 U518 ( .A(n402), .B(n688), .ZN(n689) );
  NAND2_X1 U519 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U520 ( .A(n566), .B(KEYINPUT46), .ZN(n386) );
  NAND2_X1 U521 ( .A1(n395), .A2(n392), .ZN(n611) );
  NOR2_X1 U522 ( .A1(n528), .A2(n530), .ZN(n393) );
  INV_X1 U523 ( .A(G478), .ZN(n394) );
  NOR2_X1 U524 ( .A1(n533), .A2(n399), .ZN(n535) );
  INV_X1 U525 ( .A(n560), .ZN(n399) );
  NAND2_X1 U526 ( .A1(n527), .A2(KEYINPUT44), .ZN(n423) );
  NAND2_X1 U527 ( .A1(n401), .A2(n357), .ZN(n400) );
  XNOR2_X1 U528 ( .A(n521), .B(KEYINPUT34), .ZN(n401) );
  NAND2_X1 U529 ( .A1(n708), .A2(G210), .ZN(n402) );
  NAND2_X1 U530 ( .A1(n537), .A2(n360), .ZN(n404) );
  NAND2_X1 U531 ( .A1(n407), .A2(n406), .ZN(n405) );
  NAND2_X1 U532 ( .A1(n409), .A2(n408), .ZN(n407) );
  INV_X1 U533 ( .A(n537), .ZN(n409) );
  XNOR2_X2 U534 ( .A(n411), .B(KEYINPUT0), .ZN(n533) );
  NAND2_X1 U535 ( .A1(n572), .A2(n356), .ZN(n411) );
  NAND2_X1 U536 ( .A1(n519), .A2(n615), .ZN(n426) );
  XNOR2_X2 U537 ( .A(n428), .B(KEYINPUT19), .ZN(n572) );
  NOR2_X2 U538 ( .A1(n533), .A2(n430), .ZN(n429) );
  XOR2_X2 U539 ( .A(G122), .B(G104), .Z(n471) );
  XOR2_X1 U540 ( .A(n457), .B(n456), .Z(n432) );
  INV_X1 U541 ( .A(n679), .ZN(n587) );
  INV_X1 U542 ( .A(KEYINPUT44), .ZN(n518) );
  INV_X1 U543 ( .A(KEYINPUT93), .ZN(n492) );
  XNOR2_X1 U544 ( .A(n436), .B(n473), .ZN(n437) );
  INV_X1 U545 ( .A(KEYINPUT86), .ZN(n479) );
  XNOR2_X1 U546 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U547 ( .A(n495), .B(n494), .ZN(n497) );
  XNOR2_X1 U548 ( .A(n432), .B(n458), .ZN(n459) );
  XNOR2_X1 U549 ( .A(n460), .B(n459), .ZN(n697) );
  XNOR2_X1 U550 ( .A(n502), .B(KEYINPUT25), .ZN(n503) );
  XNOR2_X1 U551 ( .A(n647), .B(n362), .ZN(n648) );
  XNOR2_X1 U552 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X1 U553 ( .A1(G952), .A2(n731), .ZN(n713) );
  XNOR2_X1 U554 ( .A(n491), .B(n433), .ZN(n436) );
  XOR2_X1 U555 ( .A(G104), .B(KEYINPUT91), .Z(n439) );
  NAND2_X1 U556 ( .A1(G227), .A2(n731), .ZN(n438) );
  XNOR2_X1 U557 ( .A(KEYINPUT69), .B(G469), .ZN(n441) );
  XNOR2_X2 U558 ( .A(n442), .B(n441), .ZN(n556) );
  XNOR2_X2 U559 ( .A(n556), .B(KEYINPUT1), .ZN(n519) );
  INV_X1 U560 ( .A(n519), .ZN(n590) );
  XNOR2_X1 U561 ( .A(KEYINPUT15), .B(G902), .ZN(n644) );
  NAND2_X1 U562 ( .A1(G234), .A2(n644), .ZN(n443) );
  XNOR2_X1 U563 ( .A(KEYINPUT20), .B(n443), .ZN(n501) );
  NAND2_X1 U564 ( .A1(n501), .A2(G221), .ZN(n444) );
  XNOR2_X1 U565 ( .A(KEYINPUT21), .B(n444), .ZN(n618) );
  XNOR2_X1 U566 ( .A(n446), .B(n445), .ZN(n449) );
  NAND2_X1 U567 ( .A1(G234), .A2(n731), .ZN(n450) );
  XOR2_X1 U568 ( .A(KEYINPUT8), .B(n450), .Z(n499) );
  NAND2_X1 U569 ( .A1(G217), .A2(n499), .ZN(n451) );
  XNOR2_X1 U570 ( .A(n452), .B(n451), .ZN(n705) );
  NOR2_X1 U571 ( .A1(G902), .A2(n705), .ZN(n453) );
  XNOR2_X1 U572 ( .A(KEYINPUT13), .B(G475), .ZN(n462) );
  XNOR2_X2 U573 ( .A(G125), .B(G146), .ZN(n465) );
  NOR2_X1 U574 ( .A1(G953), .A2(G237), .ZN(n505) );
  NAND2_X1 U575 ( .A1(G214), .A2(n505), .ZN(n455) );
  XNOR2_X1 U576 ( .A(n358), .B(n455), .ZN(n460) );
  XOR2_X1 U577 ( .A(KEYINPUT11), .B(G140), .Z(n457) );
  XNOR2_X1 U578 ( .A(G113), .B(G143), .ZN(n456) );
  XNOR2_X1 U579 ( .A(n471), .B(KEYINPUT12), .ZN(n458) );
  NOR2_X1 U580 ( .A1(G902), .A2(n697), .ZN(n461) );
  XNOR2_X1 U581 ( .A(n462), .B(n461), .ZN(n528) );
  XNOR2_X1 U582 ( .A(KEYINPUT89), .B(G898), .ZN(n718) );
  NAND2_X1 U583 ( .A1(n718), .A2(G953), .ZN(n463) );
  XOR2_X1 U584 ( .A(KEYINPUT90), .B(n463), .Z(n715) );
  NAND2_X1 U585 ( .A1(n715), .A2(G902), .ZN(n464) );
  NAND2_X1 U586 ( .A1(G952), .A2(n731), .ZN(n551) );
  NAND2_X1 U587 ( .A1(n464), .A2(n551), .ZN(n487) );
  XNOR2_X1 U588 ( .A(n465), .B(KEYINPUT72), .ZN(n468) );
  XNOR2_X1 U589 ( .A(n466), .B(KEYINPUT17), .ZN(n467) );
  XNOR2_X1 U590 ( .A(n468), .B(n467), .ZN(n482) );
  XNOR2_X1 U591 ( .A(n470), .B(n469), .ZN(n508) );
  XNOR2_X1 U592 ( .A(n472), .B(n471), .ZN(n475) );
  INV_X1 U593 ( .A(n473), .ZN(n474) );
  NAND2_X1 U594 ( .A1(G224), .A2(n731), .ZN(n477) );
  XNOR2_X1 U595 ( .A(n478), .B(n477), .ZN(n480) );
  NAND2_X1 U596 ( .A1(G210), .A2(n485), .ZN(n483) );
  NAND2_X1 U597 ( .A1(n485), .A2(G214), .ZN(n486) );
  XNOR2_X1 U598 ( .A(KEYINPUT88), .B(n486), .ZN(n609) );
  XNOR2_X1 U599 ( .A(KEYINPUT14), .B(n488), .ZN(n547) );
  INV_X1 U600 ( .A(n547), .ZN(n634) );
  XNOR2_X1 U601 ( .A(KEYINPUT64), .B(KEYINPUT22), .ZN(n489) );
  NAND2_X1 U602 ( .A1(n590), .A2(n514), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U604 ( .A1(G221), .A2(n499), .ZN(n500) );
  NAND2_X1 U605 ( .A1(n501), .A2(G217), .ZN(n502) );
  XOR2_X1 U606 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n506) );
  NAND2_X1 U607 ( .A1(n617), .A2(n560), .ZN(n511) );
  NOR2_X1 U608 ( .A1(n541), .A2(n511), .ZN(n661) );
  NAND2_X1 U609 ( .A1(n617), .A2(n584), .ZN(n512) );
  NOR2_X1 U610 ( .A1(n590), .A2(n512), .ZN(n513) );
  XNOR2_X1 U611 ( .A(KEYINPUT76), .B(n513), .ZN(n515) );
  NAND2_X1 U612 ( .A1(n515), .A2(n514), .ZN(n517) );
  NOR2_X2 U613 ( .A1(n661), .A2(n737), .ZN(n524) );
  XNOR2_X1 U614 ( .A(n524), .B(n518), .ZN(n526) );
  XNOR2_X1 U615 ( .A(n520), .B(KEYINPUT33), .ZN(n603) );
  NOR2_X1 U616 ( .A1(n533), .A2(n603), .ZN(n521) );
  NAND2_X1 U617 ( .A1(n528), .A2(n530), .ZN(n522) );
  XNOR2_X1 U618 ( .A(n522), .B(KEYINPUT102), .ZN(n568) );
  XOR2_X1 U619 ( .A(KEYINPUT84), .B(KEYINPUT35), .Z(n523) );
  NAND2_X1 U620 ( .A1(n524), .A2(n527), .ZN(n525) );
  NAND2_X1 U621 ( .A1(n526), .A2(n525), .ZN(n543) );
  XNOR2_X1 U622 ( .A(n528), .B(KEYINPUT97), .ZN(n529) );
  NOR2_X1 U623 ( .A1(n529), .A2(n530), .ZN(n669) );
  NAND2_X1 U624 ( .A1(n530), .A2(n529), .ZN(n675) );
  INV_X1 U625 ( .A(n675), .ZN(n662) );
  NOR2_X1 U626 ( .A1(n669), .A2(n662), .ZN(n606) );
  XNOR2_X1 U627 ( .A(n606), .B(KEYINPUT80), .ZN(n576) );
  INV_X1 U628 ( .A(n576), .ZN(n538) );
  INV_X1 U629 ( .A(n625), .ZN(n531) );
  NOR2_X1 U630 ( .A1(n533), .A2(n531), .ZN(n532) );
  XNOR2_X1 U631 ( .A(n532), .B(KEYINPUT31), .ZN(n674) );
  NAND2_X1 U632 ( .A1(n556), .A2(n615), .ZN(n562) );
  INV_X1 U633 ( .A(n562), .ZN(n534) );
  NAND2_X1 U634 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U635 ( .A1(n584), .A2(n539), .ZN(n540) );
  XOR2_X1 U636 ( .A(KEYINPUT83), .B(KEYINPUT45), .Z(n544) );
  INV_X1 U637 ( .A(n609), .ZN(n559) );
  XNOR2_X1 U638 ( .A(KEYINPUT38), .B(n595), .ZN(n605) );
  NOR2_X1 U639 ( .A1(n559), .A2(n611), .ZN(n546) );
  XNOR2_X1 U640 ( .A(KEYINPUT105), .B(KEYINPUT41), .ZN(n545) );
  XOR2_X1 U641 ( .A(n546), .B(n545), .Z(n604) );
  NAND2_X1 U642 ( .A1(G902), .A2(n547), .ZN(n548) );
  NOR2_X1 U643 ( .A1(G900), .A2(n548), .ZN(n549) );
  NAND2_X1 U644 ( .A1(G953), .A2(n549), .ZN(n550) );
  XNOR2_X1 U645 ( .A(n550), .B(KEYINPUT103), .ZN(n553) );
  NOR2_X1 U646 ( .A1(n634), .A2(n551), .ZN(n552) );
  NOR2_X1 U647 ( .A1(n553), .A2(n552), .ZN(n563) );
  NOR2_X1 U648 ( .A1(n563), .A2(n618), .ZN(n554) );
  NAND2_X1 U649 ( .A1(n617), .A2(n554), .ZN(n581) );
  XNOR2_X1 U650 ( .A(KEYINPUT28), .B(n555), .ZN(n557) );
  NAND2_X1 U651 ( .A1(n557), .A2(n556), .ZN(n574) );
  XNOR2_X1 U652 ( .A(n558), .B(KEYINPUT42), .ZN(n739) );
  NOR2_X1 U653 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U654 ( .A(n565), .B(KEYINPUT40), .ZN(n738) );
  NOR2_X1 U655 ( .A1(n739), .A2(n738), .ZN(n566) );
  NAND2_X1 U656 ( .A1(n606), .A2(KEYINPUT47), .ZN(n570) );
  NOR2_X1 U657 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U658 ( .A(KEYINPUT78), .B(n571), .Z(n579) );
  INV_X1 U659 ( .A(n572), .ZN(n573) );
  NAND2_X1 U660 ( .A1(KEYINPUT66), .A2(n668), .ZN(n575) );
  XNOR2_X1 U661 ( .A(n575), .B(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U662 ( .A1(n576), .A2(n668), .ZN(n577) );
  XNOR2_X1 U663 ( .A(KEYINPUT70), .B(n580), .ZN(n588) );
  INV_X1 U664 ( .A(n669), .ZN(n671) );
  NOR2_X1 U665 ( .A1(n581), .A2(n671), .ZN(n582) );
  NAND2_X1 U666 ( .A1(n609), .A2(n582), .ZN(n583) );
  NOR2_X1 U667 ( .A1(n584), .A2(n583), .ZN(n591) );
  AND2_X1 U668 ( .A1(n375), .A2(n591), .ZN(n585) );
  XNOR2_X1 U669 ( .A(n585), .B(KEYINPUT36), .ZN(n586) );
  NAND2_X1 U670 ( .A1(n586), .A2(n519), .ZN(n679) );
  NAND2_X1 U671 ( .A1(n589), .A2(n662), .ZN(n681) );
  XOR2_X1 U672 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n593) );
  NAND2_X1 U673 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U674 ( .A(n593), .B(n592), .ZN(n594) );
  NOR2_X1 U675 ( .A1(n375), .A2(n594), .ZN(n682) );
  NAND2_X1 U676 ( .A1(n643), .A2(KEYINPUT2), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n354), .A2(KEYINPUT2), .ZN(n597) );
  INV_X1 U678 ( .A(KEYINPUT77), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n602), .B(KEYINPUT82), .ZN(n640) );
  INV_X1 U680 ( .A(n603), .ZN(n613) );
  INV_X1 U681 ( .A(n604), .ZN(n627) );
  NAND2_X1 U682 ( .A1(n613), .A2(n627), .ZN(n637) );
  OR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n631) );
  NOR2_X1 U688 ( .A1(n615), .A2(n519), .ZN(n616) );
  XOR2_X1 U689 ( .A(KEYINPUT50), .B(n616), .Z(n622) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U691 ( .A(n619), .B(KEYINPUT115), .ZN(n620) );
  XNOR2_X1 U692 ( .A(KEYINPUT49), .B(n620), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U695 ( .A(KEYINPUT51), .B(n626), .ZN(n628) );
  NAND2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U697 ( .A(KEYINPUT116), .B(n629), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U699 ( .A(KEYINPUT52), .B(n632), .Z(n633) );
  NOR2_X1 U700 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U701 ( .A1(n635), .A2(G952), .ZN(n636) );
  NAND2_X1 U702 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U703 ( .A1(G953), .A2(n638), .ZN(n639) );
  NAND2_X1 U704 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U705 ( .A(KEYINPUT53), .B(KEYINPUT117), .ZN(n641) );
  XNOR2_X1 U706 ( .A(n642), .B(n641), .ZN(G75) );
  INV_X1 U707 ( .A(n686), .ZN(n646) );
  INV_X1 U708 ( .A(n644), .ZN(n687) );
  AND2_X1 U709 ( .A1(n687), .A2(G472), .ZN(n645) );
  NAND2_X1 U710 ( .A1(n646), .A2(n645), .ZN(n649) );
  NOR2_X1 U711 ( .A1(n713), .A2(n650), .ZN(n652) );
  XNOR2_X1 U712 ( .A(KEYINPUT63), .B(KEYINPUT107), .ZN(n651) );
  XNOR2_X1 U713 ( .A(n652), .B(n651), .ZN(G57) );
  XOR2_X1 U714 ( .A(n653), .B(G101), .Z(G3) );
  NOR2_X1 U715 ( .A1(n657), .A2(n671), .ZN(n655) );
  XNOR2_X1 U716 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n654) );
  XNOR2_X1 U717 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U718 ( .A(G104), .B(n656), .ZN(G6) );
  NOR2_X1 U719 ( .A1(n657), .A2(n675), .ZN(n659) );
  XNOR2_X1 U720 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n658) );
  XNOR2_X1 U721 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U722 ( .A(G107), .B(n660), .ZN(G9) );
  XOR2_X1 U723 ( .A(G110), .B(n661), .Z(G12) );
  XOR2_X1 U724 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n664) );
  NAND2_X1 U725 ( .A1(n668), .A2(n662), .ZN(n663) );
  XNOR2_X1 U726 ( .A(n664), .B(n663), .ZN(n666) );
  XOR2_X1 U727 ( .A(G128), .B(KEYINPUT110), .Z(n665) );
  XNOR2_X1 U728 ( .A(n666), .B(n665), .ZN(G30) );
  XNOR2_X1 U729 ( .A(G143), .B(n667), .ZN(G45) );
  NAND2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U731 ( .A(G146), .B(n670), .ZN(G48) );
  NOR2_X1 U732 ( .A1(n671), .A2(n674), .ZN(n672) );
  XOR2_X1 U733 ( .A(KEYINPUT112), .B(n672), .Z(n673) );
  XNOR2_X1 U734 ( .A(G113), .B(n673), .ZN(G15) );
  NOR2_X1 U735 ( .A1(n675), .A2(n674), .ZN(n677) );
  XNOR2_X1 U736 ( .A(G116), .B(KEYINPUT113), .ZN(n676) );
  XNOR2_X1 U737 ( .A(n677), .B(n676), .ZN(G18) );
  XOR2_X1 U738 ( .A(KEYINPUT37), .B(KEYINPUT114), .Z(n678) );
  XNOR2_X1 U739 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U740 ( .A(G125), .B(n680), .ZN(G27) );
  XNOR2_X1 U741 ( .A(G134), .B(n681), .ZN(G36) );
  XOR2_X1 U742 ( .A(G140), .B(n682), .Z(G42) );
  XNOR2_X1 U743 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n685) );
  XNOR2_X1 U744 ( .A(n683), .B(KEYINPUT79), .ZN(n684) );
  XOR2_X1 U745 ( .A(n685), .B(n684), .Z(n688) );
  XNOR2_X1 U746 ( .A(KEYINPUT56), .B(n690), .ZN(G51) );
  XNOR2_X1 U747 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n693) );
  XNOR2_X1 U748 ( .A(n691), .B(KEYINPUT57), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n708), .A2(G469), .ZN(n694) );
  XOR2_X1 U751 ( .A(n695), .B(n694), .Z(n696) );
  NOR2_X1 U752 ( .A1(n713), .A2(n696), .ZN(G54) );
  XOR2_X1 U753 ( .A(n697), .B(KEYINPUT59), .Z(n699) );
  NAND2_X1 U754 ( .A1(n708), .A2(G475), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U756 ( .A(KEYINPUT65), .B(KEYINPUT119), .ZN(n701) );
  XNOR2_X1 U757 ( .A(n701), .B(KEYINPUT60), .ZN(n702) );
  XNOR2_X1 U758 ( .A(n703), .B(n702), .ZN(G60) );
  XNOR2_X1 U759 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(KEYINPUT120), .ZN(G63) );
  XOR2_X1 U761 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n710) );
  NAND2_X1 U762 ( .A1(n708), .A2(G217), .ZN(n709) );
  NOR2_X1 U763 ( .A1(n713), .A2(n712), .ZN(G66) );
  NOR2_X1 U764 ( .A1(n715), .A2(n714), .ZN(n723) );
  NAND2_X1 U765 ( .A1(G953), .A2(G224), .ZN(n716) );
  XOR2_X1 U766 ( .A(KEYINPUT61), .B(n716), .Z(n717) );
  NOR2_X1 U767 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U768 ( .A(n719), .B(KEYINPUT123), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n354), .A2(n731), .ZN(n720) );
  NAND2_X1 U770 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U771 ( .A(n723), .B(n722), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n724), .B(KEYINPUT124), .ZN(n726) );
  XOR2_X1 U773 ( .A(n726), .B(n725), .Z(n729) );
  XNOR2_X1 U774 ( .A(n729), .B(n727), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(n731), .ZN(n734) );
  XOR2_X1 U776 ( .A(G227), .B(n729), .Z(n730) );
  NOR2_X1 U777 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U778 ( .A1(G900), .A2(n732), .ZN(n733) );
  NAND2_X1 U779 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U780 ( .A(KEYINPUT125), .B(n735), .ZN(G72) );
  XOR2_X1 U781 ( .A(G122), .B(n527), .Z(n736) );
  XNOR2_X1 U782 ( .A(KEYINPUT126), .B(n736), .ZN(G24) );
  XOR2_X1 U783 ( .A(G119), .B(n737), .Z(G21) );
  XOR2_X1 U784 ( .A(n738), .B(G131), .Z(G33) );
  XNOR2_X1 U785 ( .A(G137), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U786 ( .A(n740), .B(n739), .ZN(G39) );
endmodule

