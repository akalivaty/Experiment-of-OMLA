//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT68), .B1(new_n463), .B2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND4_X1   g043(.A1(KEYINPUT68), .A2(new_n466), .A3(new_n468), .A4(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  NOR3_X1   g047(.A1(new_n472), .A2(new_n465), .A3(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n466), .A2(new_n468), .A3(G137), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT69), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n463), .A2(new_n477), .A3(G137), .A4(new_n474), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n473), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n471), .A2(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n466), .A2(new_n468), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n481), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n474), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(new_n492), .A3(G138), .A4(new_n474), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n474), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n482), .A2(G126), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n511), .A3(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n507), .A2(G651), .B1(new_n513), .B2(G50), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n509), .A2(new_n511), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(new_n505), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n518), .A2(KEYINPUT70), .A3(new_n509), .A4(new_n511), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  AND2_X1   g098(.A1(new_n517), .A2(new_n519), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n512), .B(KEYINPUT71), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n525), .A2(new_n527), .A3(new_n528), .A4(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n524), .A2(G90), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n508), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT72), .B(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n505), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n524), .A2(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n526), .A2(G43), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND4_X1  g129(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT74), .A4(G543), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n555), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n508), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n517), .A2(G91), .A3(new_n519), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n559), .A2(new_n565), .A3(new_n561), .A4(new_n562), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n524), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n513), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n517), .A2(G86), .A3(new_n519), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n508), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n572), .A2(new_n573), .B1(KEYINPUT76), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n524), .A2(KEYINPUT77), .A3(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n575), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n580), .A2(new_n581), .B1(G48), .B2(new_n513), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n508), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n524), .B2(G85), .ZN(new_n586));
  INV_X1    g161(.A(new_n526), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT78), .B(G47), .Z(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OR3_X1    g166(.A1(new_n520), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT10), .B1(new_n520), .B2(new_n591), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  INV_X1    g169(.A(G79), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n505), .A2(new_n594), .B1(new_n595), .B2(new_n501), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n597), .A2(G651), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n526), .A2(G54), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n592), .A2(new_n593), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n590), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n590), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n564), .A2(new_n566), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  OAI21_X1  g185(.A(KEYINPUT80), .B1(new_n548), .B2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n609), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  MUX2_X1   g188(.A(KEYINPUT80), .B(new_n611), .S(new_n613), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g190(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2100), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n484), .A2(G135), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n622), .B(new_n623), .C1(G111), .C2(new_n474), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n482), .A2(G123), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n620), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT15), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2435), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G1341), .B(G1348), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n641), .A2(G14), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT17), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT82), .Z(new_n648));
  INV_X1    g223(.A(new_n645), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n646), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n649), .B(new_n650), .C1(new_n644), .C2(new_n646), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n649), .A2(new_n643), .A3(new_n646), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT18), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n648), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT83), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  AOI22_X1  g241(.A1(new_n664), .A2(new_n665), .B1(new_n660), .B2(new_n666), .ZN(new_n667));
  OR3_X1    g242(.A1(new_n660), .A2(new_n663), .A3(new_n666), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n667), .B(new_n668), .C1(new_n665), .C2(new_n664), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  INV_X1    g247(.A(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(KEYINPUT34), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT32), .B(G1981), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  OR2_X1    g254(.A1(G305), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(G6), .A2(G16), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n681), .A3(new_n678), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(G16), .A2(G23), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G288), .B2(new_n679), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT33), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT85), .B(G16), .ZN(new_n690));
  MUX2_X1   g265(.A(G22), .B(G303), .S(new_n690), .Z(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n677), .B1(new_n685), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n684), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(new_n682), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n697), .A2(KEYINPUT34), .A3(new_n693), .A4(new_n689), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  MUX2_X1   g274(.A(G24), .B(G290), .S(new_n690), .Z(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(G1986), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n482), .A2(G119), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n484), .A2(G131), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n474), .A2(G107), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n702), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G25), .B(new_n706), .S(G29), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT35), .B(G1991), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n707), .B(new_n708), .Z(new_n709));
  NAND3_X1  g284(.A1(new_n699), .A2(new_n701), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(KEYINPUT86), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n712), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n699), .A2(new_n714), .A3(new_n701), .A4(new_n709), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(KEYINPUT24), .A2(G34), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(KEYINPUT24), .A2(G34), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n718), .A2(new_n719), .A3(G29), .ZN(new_n720));
  INV_X1    g295(.A(G160), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G29), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT28), .ZN(new_n725));
  INV_X1    g300(.A(G26), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n482), .A2(G128), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n484), .A2(G140), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n474), .A2(G116), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n729), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n728), .B1(new_n733), .B2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(new_n725), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT89), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT88), .B(G2067), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(KEYINPUT89), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n737), .B1(new_n736), .B2(new_n738), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G4), .B2(G16), .ZN(new_n743));
  OR3_X1    g318(.A1(new_n742), .A2(G4), .A3(G16), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n743), .B(new_n744), .C1(new_n601), .C2(new_n679), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1348), .ZN(new_n746));
  INV_X1    g321(.A(G19), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n690), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n547), .B2(new_n690), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1341), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n741), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT90), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n722), .A2(new_n723), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n741), .A2(KEYINPUT90), .A3(new_n746), .A4(new_n750), .ZN(new_n755));
  NAND2_X1  g330(.A1(G171), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G5), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1961), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G27), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n760), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2078), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G11), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(G28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(G28), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n767), .A2(new_n768), .A3(new_n760), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n765), .B(new_n769), .C1(new_n626), .C2(new_n760), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT94), .Z(new_n771));
  NOR3_X1   g346(.A1(new_n759), .A2(new_n763), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n760), .A2(G35), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G162), .B2(new_n760), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT29), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G2090), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n484), .A2(G139), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n779), .B(new_n780), .C1(new_n474), .C2(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G33), .B(new_n782), .S(G29), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2072), .ZN(new_n784));
  OR2_X1    g359(.A1(G16), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G286), .B2(new_n679), .ZN(new_n786));
  INV_X1    g361(.A(G1966), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT92), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(KEYINPUT92), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n777), .B(new_n784), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G20), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n690), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT95), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT23), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1956), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n776), .A2(G2090), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(KEYINPUT96), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n786), .A2(new_n787), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n797), .A2(new_n802), .A3(new_n798), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n791), .A2(new_n800), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n773), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n716), .A2(new_n724), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n484), .A2(G141), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n482), .A2(G129), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n474), .A2(G105), .A3(G2104), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT26), .Z(new_n811));
  NAND4_X1  g386(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT91), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G32), .B(new_n814), .S(G29), .Z(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT27), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1996), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n757), .A2(new_n758), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n806), .A2(KEYINPUT97), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n716), .A2(new_n805), .A3(new_n819), .A4(new_n724), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n817), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n823), .ZN(G311));
  NAND3_X1  g399(.A1(new_n806), .A2(new_n818), .A3(new_n819), .ZN(G150));
  NAND2_X1  g400(.A1(new_n524), .A2(G93), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n508), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n526), .A2(G55), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT98), .B(G860), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND4_X1  g408(.A1(new_n547), .A2(new_n828), .A3(new_n826), .A4(new_n829), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n830), .A2(new_n545), .A3(new_n546), .A4(new_n544), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n602), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n833), .B1(new_n840), .B2(new_n831), .ZN(G145));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n484), .A2(G142), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n482), .A2(G130), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n847));
  OR3_X1    g422(.A1(new_n847), .A2(new_n474), .A3(G118), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n474), .B2(G118), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n846), .A2(new_n848), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n843), .A2(new_n844), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n782), .A2(new_n812), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n814), .B2(new_n782), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n617), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n617), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n856), .A3(new_n852), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n706), .B(new_n733), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n498), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n859), .A2(new_n861), .A3(new_n864), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G160), .B(new_n488), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n626), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n842), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n868), .B2(new_n871), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n866), .A2(new_n867), .A3(new_n870), .A4(KEYINPUT101), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g451(.A(G290), .B(G305), .ZN(new_n877));
  XNOR2_X1  g452(.A(G288), .B(G303), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT104), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(KEYINPUT104), .A3(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n882), .B1(new_n886), .B2(KEYINPUT42), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n836), .B(new_n612), .Z(new_n888));
  NAND3_X1  g463(.A1(new_n606), .A2(KEYINPUT102), .A3(new_n601), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n602), .B2(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n602), .A2(G299), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n889), .A2(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT103), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n889), .A2(new_n891), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n892), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n896), .B1(new_n901), .B2(new_n895), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n887), .B(new_n894), .C1(new_n888), .C2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n894), .B1(new_n902), .B2(new_n888), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n879), .A2(KEYINPUT104), .A3(new_n880), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n883), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(new_n908), .B2(new_n882), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n909), .A3(G868), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G868), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT105), .B1(new_n830), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n914), .B2(new_n910), .ZN(G295));
  AOI21_X1  g490(.A(new_n912), .B1(new_n914), .B2(new_n910), .ZN(G331));
  NAND2_X1  g491(.A1(G168), .A2(G301), .ZN(new_n917));
  NAND2_X1  g492(.A1(G171), .A2(G286), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n836), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n834), .A2(new_n917), .A3(new_n835), .A4(new_n918), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  INV_X1    g500(.A(new_n893), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n886), .C1(new_n902), .C2(new_n923), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n901), .A2(KEYINPUT41), .A3(new_n922), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n926), .B1(new_n923), .B2(new_n895), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n906), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n900), .A2(new_n892), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n899), .B1(new_n889), .B2(new_n891), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n895), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n896), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n922), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n886), .B1(new_n943), .B2(new_n928), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n933), .A4(new_n929), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n934), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n937), .A2(KEYINPUT44), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n929), .A2(new_n933), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n950), .B2(new_n944), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n929), .A2(new_n932), .A3(new_n946), .A4(new_n933), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n955), .ZN(G397));
  NAND3_X1  g531(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT68), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n463), .A2(KEYINPUT68), .A3(G125), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n959), .A2(new_n960), .B1(G113), .B2(G2104), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n479), .B(G40), .C1(new_n961), .C2(new_n474), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n471), .A2(KEYINPUT109), .A3(G40), .A4(new_n479), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n498), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G2067), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n733), .B(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n814), .B2(G1996), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(G1996), .B2(new_n812), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n706), .A2(new_n708), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n706), .A2(new_n708), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(G290), .B(G1986), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n971), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n498), .A2(new_n981), .A3(new_n968), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n498), .B2(new_n968), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n966), .ZN(new_n985));
  INV_X1    g560(.A(G1348), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n498), .A2(new_n968), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n964), .B2(new_n965), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n972), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n602), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n993));
  INV_X1    g568(.A(G1956), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n964), .A2(new_n965), .ZN(new_n995));
  INV_X1    g570(.A(new_n983), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n498), .A2(new_n981), .A3(new_n968), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n994), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n969), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT56), .B(G2072), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n966), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n563), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n563), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n993), .B1(new_n1004), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g588(.A(KEYINPUT117), .B(new_n1011), .C1(new_n999), .C2(new_n1003), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n992), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n999), .A2(new_n1011), .A3(new_n1003), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT61), .B(new_n1017), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1019));
  INV_X1    g594(.A(new_n988), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n966), .A2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT58), .B(G1341), .Z(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1996), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1001), .A2(new_n966), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1026), .A2(KEYINPUT59), .A3(new_n548), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT59), .B1(new_n1026), .B2(new_n548), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT60), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n991), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n601), .B(KEYINPUT119), .Z(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(new_n987), .A3(KEYINPUT60), .A4(new_n990), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n991), .A2(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n601), .A2(KEYINPUT119), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1031), .B(new_n1033), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1019), .A2(new_n1029), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1011), .B1(new_n999), .B2(new_n1003), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1016), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT118), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n1038), .C1(new_n1016), .C2(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1018), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT120), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G286), .A2(G8), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n984), .A2(new_n966), .A3(new_n723), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT113), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1020), .A2(new_n967), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n988), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n966), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n787), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n984), .A2(new_n966), .A3(new_n1055), .A4(new_n723), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1049), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1049), .A2(new_n1054), .A3(KEYINPUT121), .A4(new_n1056), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1047), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(G168), .A3(new_n1060), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1064), .A2(KEYINPUT122), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(KEYINPUT122), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1057), .A2(G8), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1061), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G2078), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1001), .A2(new_n966), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n985), .A2(new_n758), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1075), .A2(G2078), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n966), .A2(new_n1050), .A3(new_n1052), .A4(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(G301), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT125), .ZN(new_n1081));
  INV_X1    g656(.A(G40), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n474), .B1(new_n961), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n470), .A2(KEYINPUT124), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1001), .A2(new_n479), .A3(new_n1078), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1076), .A2(new_n1077), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1074), .A2(new_n1075), .B1(new_n985), .B2(new_n758), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT125), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(G301), .A4(new_n1079), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1081), .A2(new_n1089), .A3(new_n1092), .A4(KEYINPUT54), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G303), .A2(G8), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT55), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1001), .A2(new_n966), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n692), .ZN(new_n1098));
  INV_X1    g673(.A(G2090), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n984), .A2(new_n966), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1096), .B1(new_n1101), .B2(G8), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1063), .B(new_n1095), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT110), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1021), .A2(new_n1105), .A3(G8), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT110), .B1(new_n989), .B2(new_n1063), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G288), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G1976), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n513), .A2(G48), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n572), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT111), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT111), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n572), .A2(new_n1115), .A3(new_n1112), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n580), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G1981), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n578), .A2(new_n577), .A3(new_n582), .A4(new_n673), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(KEYINPUT49), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT49), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1111), .A2(KEYINPUT52), .B1(new_n1123), .B2(new_n1108), .ZN(new_n1124));
  INV_X1    g699(.A(G1976), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT52), .B1(G288), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1108), .A2(new_n1110), .A3(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1093), .A2(new_n1104), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1090), .A2(new_n1079), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G171), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1090), .A2(G301), .A3(new_n1087), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1072), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1135), .B(new_n1018), .C1(new_n1037), .C2(new_n1044), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1046), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1061), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1062), .A2(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT62), .B1(new_n1142), .B2(new_n1061), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1122), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1108), .A2(new_n1144), .A3(new_n1120), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT52), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1106), .A2(new_n1107), .B1(G1976), .B2(new_n1109), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1145), .B(new_n1127), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1148), .A2(new_n1103), .A3(new_n1102), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1131), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1141), .A2(new_n1143), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1103), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1108), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1145), .A2(new_n1125), .A3(new_n1109), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1119), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT112), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1124), .A2(new_n1103), .A3(new_n1127), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT112), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1119), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1976), .B1(new_n1123), .B2(new_n1108), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(new_n1109), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1158), .B(new_n1159), .C1(new_n1154), .C2(new_n1162), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1057), .A2(G8), .A3(G168), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1104), .A2(new_n1124), .A3(new_n1127), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT114), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(KEYINPUT63), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1148), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1167), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1169), .A2(new_n1104), .A3(new_n1170), .A4(new_n1164), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1157), .A2(new_n1163), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1151), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n980), .B1(new_n1137), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n733), .A2(G2067), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n706), .A2(new_n708), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n975), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n970), .ZN(new_n1178));
  INV_X1    g753(.A(new_n973), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n971), .B1(new_n812), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n971), .A2(KEYINPUT46), .A3(new_n1024), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT46), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n970), .B2(G1996), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT126), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT47), .Z(new_n1186));
  NAND2_X1  g761(.A1(new_n978), .A2(new_n971), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n970), .A2(G1986), .A3(G290), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT48), .Z(new_n1189));
  AOI211_X1 g764(.A(new_n1178), .B(new_n1186), .C1(new_n1187), .C2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1174), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g766(.A(G229), .ZN(new_n1193));
  AND2_X1   g767(.A1(new_n875), .A2(G319), .ZN(new_n1194));
  AOI21_X1  g768(.A(G227), .B1(new_n641), .B2(G14), .ZN(new_n1195));
  AND4_X1   g769(.A1(new_n1193), .A2(new_n953), .A3(new_n1194), .A4(new_n1195), .ZN(G308));
  NAND4_X1  g770(.A1(new_n953), .A2(new_n1194), .A3(new_n1193), .A4(new_n1195), .ZN(G225));
endmodule


