//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g0015(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(G58), .A2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n212), .B1(new_n218), .B2(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  INV_X1    g0041(.A(G107), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G97), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G107), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n223), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n248), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n215), .A2(new_n216), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n206), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n263), .B1(new_n206), .B2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n260), .A2(new_n261), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n262), .A2(new_n264), .B1(new_n266), .B2(new_n263), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT16), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n273), .B2(G20), .ZN(new_n274));
  AND2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n223), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT72), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G58), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n223), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n283), .B2(new_n219), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G159), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n279), .B2(KEYINPUT72), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n269), .B1(new_n281), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n257), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n279), .A2(new_n287), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(KEYINPUT16), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n268), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT74), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT17), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  INV_X1    g0097(.A(G226), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G1698), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n273), .B(new_n299), .C1(G223), .C2(G1698), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G87), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n217), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n303), .A2(G1), .A3(G13), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(G274), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n306), .ZN(new_n310));
  INV_X1    g0110(.A(G232), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n297), .B1(new_n305), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n217), .A2(new_n303), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n300), .B2(new_n301), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n316), .A2(new_n317), .A3(new_n312), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n295), .A2(KEYINPUT17), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n294), .A2(new_n296), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n274), .A2(new_n278), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G68), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n287), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT16), .B1(new_n326), .B2(new_n280), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n292), .A2(KEYINPUT16), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n257), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n319), .B(new_n267), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(KEYINPUT74), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n305), .A2(new_n313), .A3(G179), .ZN(new_n333));
  OAI21_X1  g0133(.A(G169), .B1(new_n316), .B2(new_n312), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(KEYINPUT73), .A3(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT18), .B1(new_n339), .B2(new_n294), .ZN(new_n340));
  INV_X1    g0140(.A(new_n338), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT73), .B1(new_n333), .B2(new_n334), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n267), .B1(new_n327), .B2(new_n329), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT18), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AND4_X1   g0146(.A1(new_n322), .A2(new_n332), .A3(new_n340), .A4(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT67), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n273), .A2(new_n349), .A3(G1698), .ZN(new_n350));
  OAI21_X1  g0150(.A(G1698), .B1(new_n275), .B2(new_n276), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT67), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n348), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G1698), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n275), .B2(new_n276), .ZN(new_n355));
  INV_X1    g0155(.A(G222), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n355), .A2(new_n356), .B1(new_n273), .B2(new_n202), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n304), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n308), .A2(G226), .A3(new_n306), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n309), .A2(new_n359), .A3(KEYINPUT66), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT66), .B1(new_n309), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n285), .A2(G150), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n207), .A2(G33), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n201), .B2(new_n207), .C1(new_n263), .C2(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n257), .B1(new_n266), .B2(new_n249), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n206), .A2(G20), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n291), .A2(new_n265), .A3(G50), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  INV_X1    g0174(.A(new_n363), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT70), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n358), .A2(new_n362), .A3(G190), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n368), .A2(new_n257), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n266), .A2(new_n249), .ZN(new_n381));
  AND4_X1   g0181(.A1(new_n379), .A2(new_n380), .A3(new_n371), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n379), .B1(new_n369), .B2(new_n371), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n377), .B(new_n378), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n363), .A2(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n372), .A2(KEYINPUT9), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n369), .A2(new_n379), .A3(new_n371), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n377), .B1(new_n389), .B2(new_n378), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT10), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT69), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT10), .B1(new_n375), .B2(G190), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n387), .A2(KEYINPUT69), .A3(new_n388), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n385), .A4(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n376), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT12), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n266), .A2(new_n398), .A3(new_n223), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT12), .B1(new_n265), .B2(G68), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n223), .B1(new_n206), .B2(G20), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n399), .A2(new_n400), .B1(new_n262), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n285), .A2(G50), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n223), .A2(G20), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n202), .C2(new_n367), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT11), .B1(new_n405), .B2(new_n257), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT71), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n408), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT71), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(new_n406), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n402), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g0214(.A(G232), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G97), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n415), .B(new_n416), .C1(new_n355), .C2(new_n298), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n304), .ZN(new_n418));
  INV_X1    g0218(.A(new_n310), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n308), .A2(G274), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n419), .A2(G238), .B1(new_n420), .B2(new_n307), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT13), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT13), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n418), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(G179), .A3(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n418), .A2(new_n421), .A3(new_n424), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n418), .B2(new_n421), .ZN(new_n428));
  OAI21_X1  g0228(.A(G169), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n426), .B1(new_n429), .B2(KEYINPUT14), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n423), .A2(new_n425), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(G169), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n414), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(G200), .B1(new_n427), .B2(new_n428), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n423), .A2(G190), .A3(new_n425), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n413), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n224), .B1(new_n350), .B2(new_n352), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n273), .A2(G232), .A3(new_n354), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n242), .B2(new_n273), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n304), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n419), .A2(G244), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n309), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(G179), .ZN(new_n444));
  INV_X1    g0244(.A(new_n263), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT15), .B(G87), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n367), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n257), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n262), .A2(G77), .A3(new_n370), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n266), .A2(new_n202), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n443), .A2(new_n364), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n444), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n443), .A2(G200), .ZN(new_n455));
  INV_X1    g0255(.A(new_n452), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n455), .B(new_n456), .C1(new_n317), .C2(new_n443), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n434), .A2(new_n437), .A3(new_n454), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n347), .A2(new_n397), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT75), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT75), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n347), .A2(new_n397), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n206), .A2(G33), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n291), .A2(new_n265), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n242), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT25), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n265), .B2(G107), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n273), .A2(new_n471), .A3(new_n207), .A4(G87), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n207), .B(G87), .C1(new_n275), .C2(new_n276), .ZN(new_n473));
  XOR2_X1   g0273(.A(KEYINPUT84), .B(KEYINPUT22), .Z(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT85), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT23), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(new_n242), .A3(G20), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT85), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n472), .A2(new_n475), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT86), .ZN(new_n485));
  AND4_X1   g0285(.A1(new_n483), .A2(new_n476), .A3(new_n477), .A4(new_n479), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT86), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n472), .A4(new_n475), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n485), .A2(KEYINPUT24), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT24), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n484), .A2(KEYINPUT86), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n257), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n470), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G41), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n206), .B(G45), .C1(new_n494), .C2(KEYINPUT5), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT78), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n500));
  AOI21_X1  g0300(.A(G41), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT79), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n496), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n504));
  NOR2_X1   g0304(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n502), .B(new_n494), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G264), .B(new_n308), .C1(new_n503), .C2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n494), .B1(new_n504), .B2(new_n505), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT79), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n506), .A3(new_n496), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n513), .A2(KEYINPUT87), .A3(G264), .A4(new_n308), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(G1698), .B1(new_n271), .B2(new_n272), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n273), .A2(G257), .A3(G1698), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n315), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n512), .A2(new_n420), .A3(new_n506), .A4(new_n496), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n297), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n508), .A3(new_n521), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n524), .A2(G190), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n493), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n519), .B1(new_n510), .B2(new_n514), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(G179), .A3(new_n521), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n524), .A2(G169), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n485), .A2(KEYINPUT24), .A3(new_n488), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n257), .A3(new_n491), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(new_n470), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n534));
  NOR2_X1   g0334(.A1(KEYINPUT81), .A2(KEYINPUT19), .ZN(new_n535));
  OAI211_X1 g0335(.A(G33), .B(G97), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  XNOR2_X1  g0337(.A(KEYINPUT82), .B(G87), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n536), .A2(new_n207), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n207), .B(G68), .C1(new_n275), .C2(new_n276), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n534), .A2(new_n535), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n367), .A2(new_n244), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n257), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n266), .A2(new_n447), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n262), .A2(G87), .A3(new_n464), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G45), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n226), .B1(new_n548), .B2(G1), .ZN(new_n549));
  INV_X1    g0349(.A(G274), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n206), .A2(new_n550), .A3(G45), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n308), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n554), .B(new_n555), .C1(new_n355), .C2(new_n224), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n553), .B1(new_n556), .B2(new_n304), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n297), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n317), .B(new_n553), .C1(new_n556), .C2(new_n304), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n547), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n447), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n262), .A2(new_n561), .A3(new_n464), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n544), .A2(new_n562), .A3(new_n545), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n304), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(G179), .A3(new_n552), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n364), .B2(new_n557), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT80), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n565), .B(KEYINPUT80), .C1(new_n364), .C2(new_n557), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n560), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n323), .A2(G107), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n285), .A2(G77), .ZN(new_n572));
  XNOR2_X1  g0372(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n573));
  MUX2_X1   g0373(.A(new_n243), .B(new_n246), .S(new_n573), .Z(new_n574));
  OAI211_X1 g0374(.A(new_n571), .B(new_n572), .C1(new_n207), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n257), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n266), .A2(new_n244), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n465), .B2(new_n244), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G244), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT77), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT77), .ZN(new_n583));
  OAI211_X1 g0383(.A(KEYINPUT4), .B(new_n582), .C1(new_n516), .C2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G250), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G283), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT4), .ZN(new_n588));
  OAI211_X1 g0388(.A(KEYINPUT77), .B(new_n588), .C1(new_n355), .C2(new_n581), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n304), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n513), .A2(G257), .A3(new_n308), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n521), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(new_n374), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n592), .A2(new_n521), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n364), .B1(new_n595), .B2(new_n591), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n580), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(G200), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n578), .B1(new_n575), .B2(new_n257), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(G190), .A3(new_n591), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n570), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G270), .ZN(new_n603));
  INV_X1    g0403(.A(new_n308), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n495), .B1(new_n511), .B2(KEYINPUT79), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n506), .ZN(new_n606));
  OAI211_X1 g0406(.A(G264), .B(G1698), .C1(new_n275), .C2(new_n276), .ZN(new_n607));
  OAI211_X1 g0407(.A(G257), .B(new_n354), .C1(new_n275), .C2(new_n276), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n271), .A2(G303), .A3(new_n272), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n304), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n521), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n262), .B2(new_n464), .ZN(new_n615));
  AOI21_X1  g0415(.A(G116), .B1(new_n260), .B2(new_n261), .ZN(new_n616));
  AOI21_X1  g0416(.A(G20), .B1(G33), .B2(G283), .ZN(new_n617));
  INV_X1    g0417(.A(G33), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G97), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n617), .A2(new_n619), .B1(G20), .B2(new_n614), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT20), .B1(new_n620), .B2(new_n257), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(new_n257), .A3(KEYINPUT20), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n615), .A2(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n613), .A2(new_n623), .A3(KEYINPUT83), .A4(G179), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT83), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n616), .B1(new_n465), .B2(G116), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n622), .A2(new_n621), .ZN(new_n627));
  OAI21_X1  g0427(.A(G179), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n513), .A2(G270), .A3(new_n308), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(new_n521), .A3(new_n611), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n623), .A2(new_n630), .A3(G169), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n623), .A2(new_n630), .A3(KEYINPUT21), .A4(G169), .ZN(new_n636));
  INV_X1    g0436(.A(new_n623), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n630), .A2(G200), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n637), .B(new_n638), .C1(new_n317), .C2(new_n630), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n632), .A2(new_n635), .A3(new_n636), .A4(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n602), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n463), .A2(new_n533), .A3(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n528), .A2(new_n529), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n493), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n635), .A2(new_n636), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n632), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n523), .A2(new_n525), .ZN(new_n647));
  INV_X1    g0447(.A(new_n493), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n593), .A2(G169), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n595), .A2(G179), .A3(new_n591), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n599), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n564), .A2(new_n552), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT88), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(G200), .ZN(new_n658));
  INV_X1    g0458(.A(new_n559), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT88), .B1(new_n557), .B2(new_n297), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n655), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n544), .A2(new_n545), .A3(new_n562), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n566), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n661), .A2(KEYINPUT89), .A3(new_n663), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n646), .A2(new_n649), .A3(new_n654), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n663), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n570), .A2(new_n653), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n651), .A2(new_n652), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n599), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT90), .ZN(new_n677));
  INV_X1    g0477(.A(new_n667), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT89), .B1(new_n661), .B2(new_n663), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n676), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n673), .B1(new_n672), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n463), .B1(new_n670), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n345), .B1(new_n344), .B2(new_n335), .ZN(new_n683));
  INV_X1    g0483(.A(new_n335), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n294), .A2(KEYINPUT18), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n454), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n429), .A2(KEYINPUT14), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n432), .A2(new_n431), .A3(G169), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n426), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n687), .A2(new_n437), .B1(new_n690), .B2(new_n414), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n332), .A2(new_n322), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n686), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n391), .A2(new_n396), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n376), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n682), .A2(new_n695), .ZN(G369));
  NAND2_X1  g0496(.A1(new_n645), .A2(new_n632), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n637), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n640), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n533), .B1(new_n648), .B2(new_n704), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n644), .B2(new_n704), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n697), .A2(new_n704), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n714), .A2(new_n533), .B1(new_n532), .B2(new_n704), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n210), .ZN(new_n717));
  OR3_X1    g0517(.A1(new_n717), .A2(KEYINPUT91), .A3(G41), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT91), .B1(new_n717), .B2(G41), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n538), .A2(new_n614), .A3(new_n537), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n221), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n671), .A2(new_n672), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n680), .B2(new_n672), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n669), .A3(new_n663), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .A3(new_n704), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n668), .A2(new_n649), .A3(new_n654), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n730), .A2(new_n646), .B1(new_n566), .B2(new_n662), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n680), .A2(new_n672), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n672), .B2(new_n671), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n703), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n729), .B1(new_n734), .B2(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n585), .A2(new_n586), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n583), .B1(new_n516), .B2(G244), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n736), .B1(new_n737), .B2(new_n588), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n315), .B1(new_n738), .B2(new_n584), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n592), .A2(new_n521), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n565), .A2(new_n606), .A3(new_n612), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n527), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n527), .A2(new_n742), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n595), .A2(KEYINPUT30), .A3(new_n591), .ZN(new_n747));
  INV_X1    g0547(.A(new_n521), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n519), .B(new_n748), .C1(new_n510), .C2(new_n514), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n557), .A2(G179), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n630), .B(new_n750), .C1(new_n739), .C2(new_n740), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n746), .A2(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n703), .B1(new_n745), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n743), .A2(new_n744), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n522), .A2(new_n630), .A3(new_n593), .A4(new_n750), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n741), .A2(new_n527), .A3(new_n742), .A4(KEYINPUT30), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT31), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(new_n759), .A3(new_n703), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n526), .A2(new_n532), .A3(new_n703), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n754), .A2(new_n760), .B1(new_n641), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G330), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n735), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n725), .B1(new_n766), .B2(G1), .ZN(G364));
  OAI21_X1  g0567(.A(new_n217), .B1(new_n207), .B2(G169), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT93), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(G20), .A2(G179), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G190), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n277), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n773), .A2(new_n317), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n207), .A2(G179), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n775), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n778), .B(new_n782), .C1(G329), .C2(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n773), .A2(new_n317), .A3(new_n297), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT94), .B(G326), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n774), .A2(new_n317), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT33), .B(G317), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G303), .A2(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n317), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n207), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n783), .A2(new_n317), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n798), .A2(G294), .B1(new_n800), .B2(G283), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n786), .A2(new_n789), .A3(new_n795), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n784), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT32), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n805), .B1(new_n223), .B2(new_n792), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n273), .B1(new_n780), .B2(new_n282), .ZN(new_n808));
  INV_X1    g0608(.A(new_n776), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(G77), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n538), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n798), .A2(G97), .B1(new_n791), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n800), .A2(G107), .B1(G50), .B2(new_n787), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n807), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n772), .B1(new_n802), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n720), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n207), .A2(G13), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n206), .B1(new_n817), .B2(G45), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(G13), .A2(G33), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(G20), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n771), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n717), .A2(new_n277), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(G355), .B1(new_n614), .B2(new_n717), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n717), .A2(new_n273), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(G45), .B2(new_n221), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n254), .A2(new_n548), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n815), .B(new_n821), .C1(new_n825), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n824), .B(KEYINPUT95), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n707), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n708), .A2(new_n821), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n707), .A2(G330), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(G396));
  INV_X1    g0637(.A(new_n787), .ZN(new_n838));
  INV_X1    g0638(.A(G303), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n838), .A2(new_n839), .B1(new_n799), .B2(new_n225), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G107), .B2(new_n791), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n273), .B1(new_n809), .B2(G116), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n785), .A2(G311), .B1(G294), .B2(new_n779), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n798), .A2(G97), .B1(new_n793), .B2(G283), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n809), .A2(G159), .B1(G143), .B2(new_n779), .ZN(new_n846));
  INV_X1    g0646(.A(G150), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n847), .B2(new_n792), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G137), .B2(new_n787), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT96), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT34), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n800), .A2(G68), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n277), .B1(new_n785), .B2(G132), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n798), .A2(G58), .B1(new_n791), .B2(G50), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n851), .A2(new_n852), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n850), .A2(KEYINPUT34), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n845), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n771), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n771), .A2(new_n822), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n820), .C1(G77), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n456), .A2(new_n704), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n454), .A2(new_n863), .A3(KEYINPUT97), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n863), .B1(new_n454), .B2(KEYINPUT97), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n457), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n861), .B1(new_n822), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n867), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n734), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n457), .B(new_n704), .C1(new_n865), .C2(new_n866), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n731), .B2(new_n733), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n764), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n821), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n875), .A2(KEYINPUT98), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(new_n764), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n875), .B2(KEYINPUT98), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n868), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT99), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n218), .A2(new_n614), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT35), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n882), .B1(new_n574), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n883), .B2(new_n574), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT36), .ZN(new_n886));
  OR3_X1    g0686(.A1(new_n221), .A2(new_n202), .A3(new_n283), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n206), .B(G13), .C1(new_n887), .C2(new_n250), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n293), .B1(KEYINPUT16), .B2(new_n292), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n701), .B1(new_n890), .B2(new_n267), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n340), .A2(new_n346), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n692), .ZN(new_n893));
  INV_X1    g0693(.A(new_n330), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n890), .A2(new_n267), .B1(new_n684), .B2(new_n701), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT37), .B1(new_n343), .B2(new_n344), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n701), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n344), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n330), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n896), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n893), .A2(new_n902), .A3(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n414), .A2(new_n703), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n434), .A2(new_n437), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n437), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n414), .B(new_n703), .C1(new_n690), .C2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n762), .A2(new_n867), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n906), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n332), .A2(new_n322), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n900), .B1(new_n917), .B2(new_n686), .ZN(new_n918));
  INV_X1    g0718(.A(new_n901), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n344), .A2(new_n335), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n900), .A3(new_n330), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n919), .A2(new_n897), .B1(new_n921), .B2(KEYINPUT37), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n916), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n905), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n913), .B1(new_n924), .B2(new_n912), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n915), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n760), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n759), .B1(new_n758), .B2(new_n703), .ZN(new_n929));
  AND4_X1   g0729(.A1(new_n632), .A2(new_n635), .A3(new_n636), .A4(new_n639), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n654), .A3(new_n570), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n649), .A2(new_n644), .A3(new_n704), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n928), .A2(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n463), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT100), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n927), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n936), .A2(new_n937), .A3(new_n763), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n924), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n690), .A2(new_n414), .A3(new_n704), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n904), .A2(KEYINPUT39), .A3(new_n905), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n871), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n670), .B2(new_n681), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n454), .A2(new_n703), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n911), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n906), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n701), .B1(new_n683), .B2(new_n685), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n729), .B(new_n463), .C1(new_n734), .C2(KEYINPUT29), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(new_n695), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n938), .A2(new_n955), .B1(new_n206), .B2(new_n817), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n938), .A2(new_n955), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n889), .B1(new_n956), .B2(new_n957), .ZN(G367));
  NAND2_X1  g0758(.A1(new_n547), .A2(new_n703), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n663), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(new_n668), .B2(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n654), .B1(new_n599), .B2(new_n704), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n676), .A2(new_n677), .A3(new_n703), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n714), .A2(new_n533), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT42), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n966), .A2(new_n532), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n703), .B1(new_n971), .B2(new_n597), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n963), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT101), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT102), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n975), .A2(KEYINPUT102), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n712), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n966), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n720), .B(KEYINPUT41), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n968), .B1(new_n711), .B2(new_n714), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(new_n709), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n766), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n715), .A2(new_n966), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n715), .A2(new_n966), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n715), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n989), .A2(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n987), .B1(new_n712), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT104), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n995), .A2(KEYINPUT103), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n980), .B1(new_n995), .B2(KEYINPUT103), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1001), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(KEYINPUT104), .A3(new_n999), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n997), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n766), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n984), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n818), .B(KEYINPUT105), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n982), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n825), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n828), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1012), .A2(new_n240), .B1(new_n210), .B2(new_n447), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n820), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n790), .A2(new_n614), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1015), .A2(KEYINPUT46), .B1(G294), .B2(new_n793), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1015), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT46), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(KEYINPUT106), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT106), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1016), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT107), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(KEYINPUT107), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n273), .B1(new_n785), .B2(G317), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n798), .A2(G107), .B1(new_n800), .B2(G97), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n809), .A2(G283), .B1(G303), .B2(new_n779), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n787), .A2(G311), .ZN(new_n1028));
  AND4_X1   g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1023), .A2(new_n1024), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT108), .Z(new_n1031));
  NAND2_X1  g0831(.A1(new_n800), .A2(G77), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n282), .B2(new_n790), .C1(new_n803), .C2(new_n792), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT109), .B(G137), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n785), .A2(new_n1034), .B1(new_n779), .B2(G150), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n273), .C1(new_n249), .C2(new_n776), .ZN(new_n1036));
  INV_X1    g0836(.A(G143), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1037), .A2(new_n838), .B1(new_n797), .B2(new_n223), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT47), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n772), .B1(new_n1040), .B2(KEYINPUT47), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1014), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n962), .A2(new_n833), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1010), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(G387));
  OAI21_X1  g0848(.A(new_n828), .B1(new_n237), .B2(new_n548), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n826), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n721), .B2(new_n1050), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n263), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1052));
  AOI21_X1  g0852(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1053));
  OAI21_X1  g0853(.A(KEYINPUT50), .B1(new_n263), .B2(G50), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1052), .A2(new_n721), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1051), .A2(new_n1055), .B1(new_n242), .B2(new_n717), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n820), .B1(new_n1056), .B2(new_n1011), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n277), .B1(new_n785), .B2(G150), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n202), .B2(new_n790), .C1(new_n244), .C2(new_n799), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT110), .Z(new_n1060));
  NOR2_X1   g0860(.A1(new_n797), .A2(new_n447), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n809), .A2(G68), .B1(G50), .B2(new_n779), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n263), .B2(new_n792), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(G159), .C2(new_n787), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n273), .B1(new_n785), .B2(new_n788), .ZN(new_n1066));
  INV_X1    g0866(.A(G283), .ZN(new_n1067));
  INV_X1    g0867(.A(G294), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n797), .A2(new_n1067), .B1(new_n790), .B2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n809), .A2(G303), .B1(G317), .B2(new_n779), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n777), .B2(new_n792), .C1(new_n781), .C2(new_n838), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1069), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1066), .B1(new_n614), .B2(new_n799), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1065), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT111), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1080), .A2(new_n771), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1057), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n711), .B2(new_n833), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT112), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n986), .B2(new_n1008), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n987), .A2(new_n816), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n766), .A2(new_n986), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(G393));
  XNOR2_X1  g0889(.A(new_n995), .B(new_n980), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n987), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n816), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1004), .A2(new_n1002), .ZN(new_n1094));
  OAI211_X1 g0894(.A(KEYINPUT114), .B(new_n1093), .C1(new_n1094), .C2(new_n997), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n1005), .B2(new_n1092), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1012), .A2(new_n248), .B1(new_n244), .B2(new_n210), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n820), .B1(new_n1011), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n798), .A2(G77), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n223), .B2(new_n790), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n273), .B1(new_n784), .B2(new_n1037), .C1(new_n263), .C2(new_n776), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n799), .A2(new_n225), .B1(new_n792), .B2(new_n249), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G150), .A2(new_n787), .B1(new_n779), .B2(G159), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT51), .Z(new_n1107));
  AOI22_X1  g0907(.A1(G317), .A2(new_n787), .B1(new_n779), .B2(G311), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT52), .Z(new_n1109));
  OAI221_X1 g0909(.A(new_n277), .B1(new_n776), .B2(new_n1068), .C1(new_n781), .C2(new_n784), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n797), .A2(new_n614), .B1(new_n790), .B2(new_n1067), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n799), .A2(new_n242), .B1(new_n792), .B2(new_n839), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1105), .A2(new_n1107), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT113), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n772), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1100), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n824), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1118), .B1(new_n966), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1090), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n1009), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1098), .A2(new_n1123), .ZN(G390));
  INV_X1    g0924(.A(KEYINPUT119), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n463), .A2(new_n764), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n953), .A2(new_n695), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT117), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n946), .A2(new_n948), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n911), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n754), .A2(new_n760), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n641), .A2(new_n761), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n867), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1133), .B2(G330), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n762), .A2(new_n763), .A3(new_n867), .A4(new_n911), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1128), .B(new_n1129), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n933), .A2(G330), .A3(new_n869), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n911), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(G330), .A3(new_n1130), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n728), .A2(new_n704), .A3(new_n869), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n948), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1128), .B1(new_n1143), .B2(new_n1129), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1127), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT118), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT118), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1127), .B(new_n1147), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n942), .B1(new_n923), .B2(new_n905), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1140), .A2(new_n948), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n911), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n905), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1152), .A2(new_n903), .A3(new_n939), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT39), .B1(new_n923), .B2(new_n905), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n949), .A2(new_n942), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1135), .A2(KEYINPUT116), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1151), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT116), .B1(new_n1135), .B2(KEYINPUT115), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1158), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1151), .A2(new_n1155), .A3(new_n1160), .A4(new_n1156), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1146), .A2(new_n1148), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1125), .B1(new_n1162), .B2(new_n720), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1148), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1129), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT117), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n1141), .A3(new_n1136), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1147), .B1(new_n1168), .B2(new_n1127), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1164), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(KEYINPUT119), .A3(new_n816), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1163), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n822), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n780), .A2(new_n614), .B1(new_n776), .B2(new_n244), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n273), .B(new_n1176), .C1(G294), .C2(new_n785), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n838), .A2(new_n1067), .B1(new_n242), .B2(new_n792), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G87), .B2(new_n791), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1177), .A2(new_n852), .A3(new_n1101), .A4(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT54), .B(G143), .ZN(new_n1181));
  INV_X1    g0981(.A(G125), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n776), .A2(new_n1181), .B1(new_n784), .B2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n277), .B(new_n1183), .C1(G132), .C2(new_n779), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n790), .A2(new_n847), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT53), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G50), .A2(new_n800), .B1(new_n793), .B2(new_n1034), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n798), .A2(G159), .B1(G128), .B2(new_n787), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n772), .B1(new_n1180), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n821), .B(new_n1190), .C1(new_n263), .C2(new_n859), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT120), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1164), .A2(new_n1008), .B1(new_n1175), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1174), .A2(new_n1193), .ZN(G378));
  AND3_X1   g0994(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n1195));
  OAI21_X1  g0995(.A(G330), .B1(new_n915), .B2(new_n925), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n925), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n763), .B1(new_n1198), .B2(new_n914), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n952), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n372), .A2(new_n899), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n397), .B(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT122), .ZN(new_n1203));
  XOR2_X1   g1003(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1204));
  XNOR2_X1  g1004(.A(new_n1203), .B(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1197), .A2(new_n1200), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1205), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(new_n823), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(G33), .A2(G41), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G50), .B(new_n1211), .C1(new_n277), .C2(new_n494), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n800), .A2(G58), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n244), .B2(new_n792), .C1(new_n614), .C2(new_n838), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n494), .B(new_n277), .C1(new_n784), .C2(new_n1067), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n780), .A2(new_n242), .B1(new_n447), .B2(new_n776), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n797), .A2(new_n223), .B1(new_n790), .B2(new_n202), .ZN(new_n1217));
  OR4_X1    g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT58), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1212), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1219), .B2(new_n1218), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n798), .A2(G150), .B1(G125), .B2(new_n787), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT121), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n809), .A2(G137), .B1(G128), .B2(new_n779), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n790), .B2(new_n1181), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G132), .B2(new_n793), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1228));
  INV_X1    g1028(.A(G124), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1211), .B1(new_n784), .B2(new_n1229), .C1(new_n803), .C2(new_n799), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1227), .B2(KEYINPUT59), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1221), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n820), .B1(G50), .B2(new_n860), .C1(new_n1232), .C2(new_n772), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1208), .A2(new_n1009), .B1(new_n1210), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1209), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1197), .A2(new_n1200), .A3(new_n1205), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1127), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(KEYINPUT57), .C1(new_n1240), .C2(new_n1162), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n816), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1170), .A2(new_n1127), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT57), .B1(new_n1243), .B2(new_n1239), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1235), .B1(new_n1242), .B2(new_n1244), .ZN(G375));
  NAND4_X1  g1045(.A1(new_n1240), .A2(new_n1167), .A3(new_n1141), .A4(new_n1136), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1172), .A2(new_n984), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n911), .A2(new_n822), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n820), .B1(new_n860), .B2(G68), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n780), .A2(new_n1067), .B1(new_n776), .B2(new_n242), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n273), .B(new_n1250), .C1(G303), .C2(new_n785), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1061), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n838), .A2(new_n1068), .B1(new_n614), .B2(new_n792), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G97), .B2(new_n791), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1251), .A2(new_n1032), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n273), .B1(new_n776), .B2(new_n847), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1213), .B1(new_n803), .B2(new_n790), .C1(new_n249), .C2(new_n797), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(G128), .C2(new_n785), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT123), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n787), .A2(G132), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1181), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n793), .A2(new_n1261), .B1(new_n779), .B2(new_n1034), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1258), .A2(KEYINPUT123), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1255), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1249), .B1(new_n1265), .B2(new_n771), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1168), .A2(new_n1008), .B1(new_n1248), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1247), .A2(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT124), .ZN(G381));
  AND3_X1   g1069(.A1(new_n1174), .A2(KEYINPUT125), .A3(new_n1193), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT125), .B1(new_n1174), .B2(new_n1193), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1244), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n816), .A3(new_n1241), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n1235), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1122), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1047), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  OR3_X1    g1078(.A1(new_n1275), .A2(new_n1278), .A3(G381), .ZN(G407));
  OAI211_X1 g1079(.A(G407), .B(G213), .C1(G343), .C2(new_n1275), .ZN(G409));
  NAND2_X1  g1080(.A1(new_n702), .A2(G213), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1246), .A2(KEYINPUT126), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n720), .B1(new_n1282), .B2(KEYINPUT60), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1246), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1283), .B1(KEYINPUT60), .B2(new_n1282), .C1(new_n1172), .C2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n880), .B1(new_n1285), .B2(new_n1267), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n880), .A3(new_n1267), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1162), .A2(new_n1240), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(new_n1208), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1234), .B1(new_n1291), .B2(new_n984), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1270), .A2(new_n1271), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(G378), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(G375), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1281), .B(new_n1289), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1281), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1281), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1288), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G2897), .B(new_n1299), .C1(new_n1300), .C2(new_n1286), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(G2897), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1287), .A2(new_n1288), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT125), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G378), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1291), .A2(new_n984), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1235), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1174), .A2(KEYINPUT125), .A3(new_n1193), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1274), .A2(G378), .A3(new_n1235), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT62), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1281), .A4(new_n1289), .ZN(new_n1315));
  XOR2_X1   g1115(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1316));
  NAND4_X1  g1116(.A1(new_n1297), .A2(new_n1305), .A3(new_n1315), .A4(new_n1316), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G390), .B(new_n1045), .C1(new_n1318), .C2(new_n982), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1276), .B1(new_n1010), .B2(new_n1046), .ZN(new_n1320));
  XOR2_X1   g1120(.A(G393), .B(G396), .Z(new_n1321));
  AND3_X1   g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1323));
  OR2_X1    g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1317), .A2(new_n1324), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1322), .A2(new_n1323), .A3(KEYINPUT61), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1296), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1281), .A4(new_n1289), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1326), .A2(new_n1305), .A3(new_n1328), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1325), .A2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(new_n1272), .A2(G375), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1332), .A2(new_n1312), .A3(new_n1289), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1289), .B1(new_n1332), .B2(new_n1312), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1335), .B(new_n1324), .ZN(G402));
endmodule


