

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754;

  XNOR2_X1 U378 ( .A(n358), .B(n357), .ZN(G51) );
  INV_X1 U379 ( .A(KEYINPUT56), .ZN(n357) );
  AND2_X1 U380 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U381 ( .A1(n360), .A2(n402), .ZN(n604) );
  AND2_X1 U382 ( .A1(n523), .A2(n524), .ZN(n526) );
  XNOR2_X1 U383 ( .A(n557), .B(n512), .ZN(n533) );
  XNOR2_X1 U384 ( .A(n511), .B(G472), .ZN(n557) );
  OR2_X1 U385 ( .A1(n630), .A2(G902), .ZN(n511) );
  XNOR2_X1 U386 ( .A(n515), .B(n514), .ZN(n743) );
  OR2_X2 U387 ( .A1(n718), .A2(G902), .ZN(n393) );
  NAND2_X1 U388 ( .A1(n709), .A2(G475), .ZN(n646) );
  AND2_X2 U389 ( .A1(n629), .A2(n367), .ZN(n709) );
  NAND2_X1 U390 ( .A1(n716), .A2(n715), .ZN(n358) );
  NAND2_X1 U391 ( .A1(n359), .A2(n366), .ZN(n567) );
  AND2_X2 U392 ( .A1(n559), .A2(n533), .ZN(n513) );
  NAND2_X2 U393 ( .A1(n605), .A2(n580), .ZN(n597) );
  XNOR2_X2 U394 ( .A(n604), .B(n372), .ZN(n614) );
  NOR2_X1 U395 ( .A1(n531), .A2(n532), .ZN(n381) );
  INV_X4 U396 ( .A(G953), .ZN(n496) );
  XNOR2_X1 U397 ( .A(n391), .B(n371), .ZN(n600) );
  AND2_X1 U398 ( .A1(n380), .A2(n535), .ZN(n547) );
  XNOR2_X1 U399 ( .A(n381), .B(KEYINPUT74), .ZN(n380) );
  XNOR2_X1 U400 ( .A(n400), .B(KEYINPUT19), .ZN(n586) );
  XNOR2_X1 U401 ( .A(n414), .B(KEYINPUT75), .ZN(n419) );
  NAND2_X1 U402 ( .A1(n496), .A2(G224), .ZN(n414) );
  XNOR2_X1 U403 ( .A(G113), .B(G104), .ZN(n463) );
  NOR2_X4 U404 ( .A1(n623), .A2(n622), .ZN(n744) );
  XNOR2_X2 U405 ( .A(n567), .B(KEYINPUT48), .ZN(n623) );
  NOR2_X1 U406 ( .A1(n591), .A2(n696), .ZN(n412) );
  AND2_X1 U407 ( .A1(n637), .A2(n754), .ZN(n615) );
  XNOR2_X1 U408 ( .A(n399), .B(n587), .ZN(n592) );
  NAND2_X1 U409 ( .A1(n638), .A2(KEYINPUT44), .ZN(n390) );
  XNOR2_X1 U410 ( .A(n409), .B(n408), .ZN(n389) );
  INV_X1 U411 ( .A(KEYINPUT108), .ZN(n408) );
  NAND2_X1 U412 ( .A1(n616), .A2(n615), .ZN(n384) );
  NAND2_X1 U413 ( .A1(n612), .A2(n415), .ZN(n385) );
  NOR2_X1 U414 ( .A1(n615), .A2(KEYINPUT44), .ZN(n415) );
  NOR2_X1 U415 ( .A1(n752), .A2(n753), .ZN(n382) );
  INV_X1 U416 ( .A(KEYINPUT110), .ZN(n417) );
  XNOR2_X1 U417 ( .A(n448), .B(n447), .ZN(n475) );
  NAND2_X1 U418 ( .A1(n496), .A2(G234), .ZN(n448) );
  XNOR2_X1 U419 ( .A(n436), .B(n435), .ZN(n539) );
  OR2_X1 U420 ( .A1(n640), .A2(G902), .ZN(n489) );
  NOR2_X1 U421 ( .A1(n597), .A2(n581), .ZN(n686) );
  XNOR2_X1 U422 ( .A(n594), .B(n416), .ZN(n606) );
  INV_X1 U423 ( .A(KEYINPUT22), .ZN(n416) );
  NAND2_X1 U424 ( .A1(n367), .A2(n377), .ZN(n376) );
  NAND2_X1 U425 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U426 ( .A(KEYINPUT2), .ZN(n378) );
  INV_X1 U427 ( .A(KEYINPUT84), .ZN(n674) );
  XNOR2_X1 U428 ( .A(n386), .B(KEYINPUT45), .ZN(n619) );
  NAND2_X1 U429 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U430 ( .A1(n392), .A2(n608), .ZN(n391) );
  XNOR2_X1 U431 ( .A(n597), .B(n417), .ZN(n392) );
  AND2_X1 U432 ( .A1(n405), .A2(n603), .ZN(n404) );
  NAND2_X1 U433 ( .A1(n598), .A2(KEYINPUT34), .ZN(n405) );
  NAND2_X1 U434 ( .A1(n403), .A2(KEYINPUT34), .ZN(n402) );
  XNOR2_X1 U435 ( .A(n446), .B(n445), .ZN(n450) );
  NAND2_X1 U436 ( .A1(n401), .A2(n691), .ZN(n400) );
  XNOR2_X1 U437 ( .A(n456), .B(n455), .ZN(n550) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n640) );
  XNOR2_X1 U439 ( .A(n741), .B(n477), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n483), .B(n368), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n383), .B(KEYINPUT40), .ZN(n752) );
  AND2_X1 U442 ( .A1(n576), .A2(n665), .ZN(n383) );
  NAND2_X1 U443 ( .A1(n686), .A2(n592), .ZN(n413) );
  NAND2_X1 U444 ( .A1(n396), .A2(n676), .ZN(n637) );
  XNOR2_X1 U445 ( .A(n398), .B(n397), .ZN(n396) );
  INV_X1 U446 ( .A(KEYINPUT64), .ZN(n397) );
  NOR2_X1 U447 ( .A1(n395), .A2(n394), .ZN(n708) );
  NAND2_X1 U448 ( .A1(n707), .A2(n496), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n376), .B(n674), .ZN(n395) );
  INV_X1 U450 ( .A(n598), .ZN(n599) );
  AND2_X1 U451 ( .A1(n566), .A2(n672), .ZN(n359) );
  AND2_X1 U452 ( .A1(n406), .A2(n404), .ZN(n360) );
  NOR2_X1 U453 ( .A1(n687), .A2(n686), .ZN(n361) );
  XOR2_X1 U454 ( .A(n443), .B(n442), .Z(n362) );
  NOR2_X1 U455 ( .A1(n605), .A2(n533), .ZN(n363) );
  XOR2_X1 U456 ( .A(n661), .B(KEYINPUT82), .Z(n364) );
  NOR2_X1 U457 ( .A1(n699), .A2(n403), .ZN(n365) );
  XOR2_X1 U458 ( .A(n382), .B(n538), .Z(n366) );
  NAND2_X1 U459 ( .A1(n617), .A2(n729), .ZN(n367) );
  BUF_X1 U460 ( .A(n539), .Z(n573) );
  INV_X1 U461 ( .A(n539), .ZN(n401) );
  AND2_X1 U462 ( .A1(n475), .A2(G221), .ZN(n368) );
  AND2_X1 U463 ( .A1(n610), .A2(n609), .ZN(n369) );
  AND2_X1 U464 ( .A1(n681), .A2(n595), .ZN(n370) );
  XOR2_X1 U465 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n371) );
  XOR2_X1 U466 ( .A(KEYINPUT86), .B(KEYINPUT35), .Z(n372) );
  XNOR2_X1 U467 ( .A(n743), .B(n522), .ZN(n718) );
  XNOR2_X1 U468 ( .A(n713), .B(n712), .ZN(n373) );
  NAND2_X1 U469 ( .A1(n744), .A2(n729), .ZN(n379) );
  NAND2_X1 U470 ( .A1(n547), .A2(n692), .ZN(n537) );
  NAND2_X1 U471 ( .A1(n385), .A2(n384), .ZN(n387) );
  XNOR2_X1 U472 ( .A(n523), .B(n564), .ZN(n568) );
  XNOR2_X2 U473 ( .A(n393), .B(G469), .ZN(n523) );
  NAND2_X1 U474 ( .A1(n606), .A2(n363), .ZN(n398) );
  NAND2_X1 U475 ( .A1(n589), .A2(n523), .ZN(n590) );
  NAND2_X1 U476 ( .A1(n586), .A2(n585), .ZN(n399) );
  INV_X1 U477 ( .A(n568), .ZN(n605) );
  INV_X1 U478 ( .A(n600), .ZN(n403) );
  NAND2_X1 U479 ( .A1(n600), .A2(n407), .ZN(n406) );
  AND2_X1 U480 ( .A1(n599), .A2(n601), .ZN(n407) );
  NAND2_X1 U481 ( .A1(n410), .A2(n596), .ZN(n409) );
  XNOR2_X1 U482 ( .A(n412), .B(n411), .ZN(n410) );
  INV_X1 U483 ( .A(KEYINPUT106), .ZN(n411) );
  XNOR2_X2 U484 ( .A(n413), .B(KEYINPUT31), .ZN(n669) );
  NAND2_X1 U485 ( .A1(n606), .A2(n369), .ZN(n611) );
  NAND2_X1 U486 ( .A1(n606), .A2(n370), .ZN(n596) );
  NOR2_X2 U487 ( .A1(n552), .A2(n551), .ZN(n661) );
  BUF_X1 U488 ( .A(n709), .Z(n724) );
  INV_X1 U489 ( .A(KEYINPUT8), .ZN(n447) );
  XNOR2_X1 U490 ( .A(n441), .B(n362), .ZN(n446) );
  BUF_X1 U491 ( .A(n557), .Z(n679) );
  BUF_X1 U492 ( .A(n619), .Z(n729) );
  XNOR2_X1 U493 ( .A(n454), .B(n453), .ZN(n455) );
  BUF_X1 U494 ( .A(n568), .Z(n681) );
  INV_X1 U495 ( .A(n728), .ZN(n715) );
  INV_X1 U496 ( .A(KEYINPUT63), .ZN(n635) );
  XOR2_X1 U497 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n418) );
  XNOR2_X1 U498 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U499 ( .A(G146), .B(G125), .ZN(n461) );
  XNOR2_X1 U500 ( .A(KEYINPUT70), .B(G110), .ZN(n519) );
  XNOR2_X1 U501 ( .A(n461), .B(n519), .ZN(n420) );
  XNOR2_X1 U502 ( .A(n421), .B(n420), .ZN(n423) );
  XNOR2_X2 U503 ( .A(G143), .B(KEYINPUT78), .ZN(n422) );
  XNOR2_X2 U504 ( .A(n422), .B(G128), .ZN(n441) );
  XNOR2_X2 U505 ( .A(n441), .B(KEYINPUT4), .ZN(n502) );
  XNOR2_X1 U506 ( .A(n502), .B(n423), .ZN(n429) );
  XNOR2_X1 U507 ( .A(G119), .B(G116), .ZN(n424) );
  XNOR2_X1 U508 ( .A(n424), .B(KEYINPUT3), .ZN(n426) );
  XNOR2_X1 U509 ( .A(G101), .B(KEYINPUT68), .ZN(n425) );
  XNOR2_X1 U510 ( .A(n426), .B(n425), .ZN(n508) );
  XNOR2_X1 U511 ( .A(n463), .B(KEYINPUT16), .ZN(n427) );
  INV_X1 U512 ( .A(G122), .ZN(n639) );
  XNOR2_X1 U513 ( .A(n639), .B(G107), .ZN(n444) );
  XNOR2_X1 U514 ( .A(n427), .B(n444), .ZN(n428) );
  XNOR2_X1 U515 ( .A(n508), .B(n428), .ZN(n734) );
  XNOR2_X1 U516 ( .A(n429), .B(n734), .ZN(n712) );
  XNOR2_X1 U517 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n430) );
  XNOR2_X1 U518 ( .A(n430), .B(G902), .ZN(n625) );
  NAND2_X1 U519 ( .A1(n712), .A2(n625), .ZN(n436) );
  NOR2_X1 U520 ( .A1(G902), .A2(G237), .ZN(n432) );
  INV_X1 U521 ( .A(KEYINPUT73), .ZN(n431) );
  XNOR2_X1 U522 ( .A(n432), .B(n431), .ZN(n438) );
  INV_X1 U523 ( .A(n438), .ZN(n433) );
  AND2_X1 U524 ( .A1(n433), .A2(G210), .ZN(n434) );
  XNOR2_X1 U525 ( .A(n434), .B(KEYINPUT93), .ZN(n435) );
  XNOR2_X1 U526 ( .A(n573), .B(KEYINPUT38), .ZN(n692) );
  INV_X1 U527 ( .A(G214), .ZN(n437) );
  OR2_X1 U528 ( .A1(n438), .A2(n437), .ZN(n691) );
  NAND2_X1 U529 ( .A1(n692), .A2(n691), .ZN(n695) );
  XOR2_X1 U530 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n440) );
  XNOR2_X1 U531 ( .A(G134), .B(G116), .ZN(n439) );
  XNOR2_X1 U532 ( .A(n440), .B(n439), .ZN(n452) );
  XOR2_X1 U533 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n443) );
  XNOR2_X1 U534 ( .A(KEYINPUT101), .B(KEYINPUT7), .ZN(n442) );
  XNOR2_X1 U535 ( .A(n444), .B(KEYINPUT100), .ZN(n445) );
  NAND2_X1 U536 ( .A1(G217), .A2(n475), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U538 ( .A(n452), .B(n451), .ZN(n725) );
  NOR2_X1 U539 ( .A1(G902), .A2(n725), .ZN(n456) );
  INV_X1 U540 ( .A(G478), .ZN(n454) );
  INV_X1 U541 ( .A(KEYINPUT105), .ZN(n453) );
  INV_X1 U542 ( .A(n550), .ZN(n473) );
  XOR2_X1 U543 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n458) );
  XNOR2_X1 U544 ( .A(G122), .B(KEYINPUT98), .ZN(n457) );
  XNOR2_X1 U545 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U546 ( .A(KEYINPUT67), .B(G131), .ZN(n500) );
  XNOR2_X1 U547 ( .A(n459), .B(n500), .ZN(n462) );
  INV_X1 U548 ( .A(KEYINPUT10), .ZN(n460) );
  XNOR2_X1 U549 ( .A(n461), .B(n460), .ZN(n741) );
  XNOR2_X1 U550 ( .A(n462), .B(n741), .ZN(n469) );
  NOR2_X1 U551 ( .A1(G953), .A2(G237), .ZN(n505) );
  NAND2_X1 U552 ( .A1(G214), .A2(n505), .ZN(n464) );
  XNOR2_X1 U553 ( .A(n464), .B(n463), .ZN(n467) );
  XNOR2_X1 U554 ( .A(G143), .B(G140), .ZN(n465) );
  XNOR2_X1 U555 ( .A(n465), .B(KEYINPUT12), .ZN(n466) );
  XNOR2_X1 U556 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U557 ( .A(n469), .B(n468), .ZN(n644) );
  INV_X1 U558 ( .A(G902), .ZN(n470) );
  NAND2_X1 U559 ( .A1(n644), .A2(n470), .ZN(n472) );
  XNOR2_X1 U560 ( .A(KEYINPUT13), .B(G475), .ZN(n471) );
  XNOR2_X1 U561 ( .A(n472), .B(n471), .ZN(n548) );
  NAND2_X1 U562 ( .A1(n473), .A2(n548), .ZN(n694) );
  NOR2_X1 U563 ( .A1(n695), .A2(n694), .ZN(n474) );
  XNOR2_X1 U564 ( .A(n474), .B(KEYINPUT41), .ZN(n704) );
  INV_X1 U565 ( .A(G140), .ZN(n476) );
  XNOR2_X1 U566 ( .A(n476), .B(G137), .ZN(n514) );
  INV_X1 U567 ( .A(n514), .ZN(n477) );
  XNOR2_X1 U568 ( .A(G119), .B(KEYINPUT24), .ZN(n479) );
  XNOR2_X1 U569 ( .A(KEYINPUT69), .B(KEYINPUT95), .ZN(n478) );
  XNOR2_X1 U570 ( .A(n479), .B(n478), .ZN(n482) );
  XNOR2_X1 U571 ( .A(G128), .B(G110), .ZN(n480) );
  XNOR2_X1 U572 ( .A(n480), .B(KEYINPUT23), .ZN(n481) );
  XNOR2_X1 U573 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U574 ( .A1(n625), .A2(G234), .ZN(n485) );
  XOR2_X1 U575 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n484) );
  XNOR2_X1 U576 ( .A(n485), .B(n484), .ZN(n490) );
  AND2_X1 U577 ( .A1(n490), .A2(G217), .ZN(n487) );
  XNOR2_X1 U578 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n486) );
  XNOR2_X1 U579 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X2 U580 ( .A(n489), .B(n488), .ZN(n607) );
  NAND2_X1 U581 ( .A1(n490), .A2(G221), .ZN(n491) );
  XNOR2_X1 U582 ( .A(n491), .B(KEYINPUT21), .ZN(n675) );
  INV_X1 U583 ( .A(n675), .ZN(n528) );
  NAND2_X1 U584 ( .A1(G234), .A2(G237), .ZN(n492) );
  XNOR2_X1 U585 ( .A(n492), .B(KEYINPUT14), .ZN(n495) );
  NAND2_X1 U586 ( .A1(G902), .A2(n495), .ZN(n493) );
  XOR2_X1 U587 ( .A(KEYINPUT94), .B(n493), .Z(n494) );
  NAND2_X1 U588 ( .A1(G953), .A2(n494), .ZN(n582) );
  NOR2_X1 U589 ( .A1(G900), .A2(n582), .ZN(n498) );
  NAND2_X1 U590 ( .A1(G952), .A2(n495), .ZN(n703) );
  OR2_X1 U591 ( .A1(n703), .A2(G953), .ZN(n583) );
  INV_X1 U592 ( .A(n583), .ZN(n497) );
  OR2_X1 U593 ( .A1(n498), .A2(n497), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n528), .A2(n530), .ZN(n499) );
  NOR2_X1 U595 ( .A1(n607), .A2(n499), .ZN(n559) );
  XNOR2_X1 U596 ( .A(n500), .B(G134), .ZN(n501) );
  XNOR2_X2 U597 ( .A(n502), .B(n501), .ZN(n515) );
  XOR2_X1 U598 ( .A(G113), .B(KEYINPUT5), .Z(n504) );
  XNOR2_X1 U599 ( .A(G137), .B(G146), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n504), .B(n503), .ZN(n507) );
  NAND2_X1 U601 ( .A1(n505), .A2(G210), .ZN(n506) );
  XNOR2_X1 U602 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U603 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U604 ( .A(n515), .B(n510), .ZN(n630) );
  INV_X1 U605 ( .A(KEYINPUT109), .ZN(n512) );
  XNOR2_X1 U606 ( .A(n513), .B(KEYINPUT28), .ZN(n524) );
  XOR2_X1 U607 ( .A(G104), .B(G107), .Z(n517) );
  XNOR2_X1 U608 ( .A(G101), .B(G146), .ZN(n516) );
  XNOR2_X1 U609 ( .A(n517), .B(n516), .ZN(n521) );
  NAND2_X1 U610 ( .A1(n496), .A2(G227), .ZN(n518) );
  XNOR2_X1 U611 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U612 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U613 ( .A(n523), .ZN(n532) );
  INV_X1 U614 ( .A(KEYINPUT114), .ZN(n525) );
  XNOR2_X1 U615 ( .A(n526), .B(n525), .ZN(n541) );
  NOR2_X1 U616 ( .A1(n704), .A2(n541), .ZN(n527) );
  XNOR2_X1 U617 ( .A(n527), .B(KEYINPUT42), .ZN(n753) );
  NOR2_X1 U618 ( .A1(n548), .A2(n550), .ZN(n665) );
  NAND2_X1 U619 ( .A1(n607), .A2(n528), .ZN(n529) );
  XNOR2_X1 U620 ( .A(n529), .B(KEYINPUT66), .ZN(n588) );
  INV_X1 U621 ( .A(n588), .ZN(n580) );
  NAND2_X1 U622 ( .A1(n580), .A2(n530), .ZN(n531) );
  NAND2_X1 U623 ( .A1(n533), .A2(n691), .ZN(n534) );
  XOR2_X1 U624 ( .A(KEYINPUT30), .B(n534), .Z(n535) );
  XNOR2_X1 U625 ( .A(KEYINPUT88), .B(KEYINPUT39), .ZN(n536) );
  XNOR2_X1 U626 ( .A(n537), .B(n536), .ZN(n576) );
  XNOR2_X1 U627 ( .A(KEYINPUT46), .B(KEYINPUT87), .ZN(n538) );
  INV_X1 U628 ( .A(n586), .ZN(n540) );
  NOR2_X1 U629 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X2 U630 ( .A(n542), .B(KEYINPUT77), .ZN(n656) );
  AND2_X1 U631 ( .A1(n550), .A2(n548), .ZN(n668) );
  NOR2_X1 U632 ( .A1(n665), .A2(n668), .ZN(n696) );
  NOR2_X1 U633 ( .A1(n656), .A2(n696), .ZN(n543) );
  NOR2_X1 U634 ( .A1(n543), .A2(KEYINPUT81), .ZN(n544) );
  XNOR2_X1 U635 ( .A(n544), .B(KEYINPUT47), .ZN(n555) );
  INV_X1 U636 ( .A(n696), .ZN(n545) );
  NAND2_X1 U637 ( .A1(n656), .A2(n545), .ZN(n546) );
  NAND2_X1 U638 ( .A1(KEYINPUT81), .A2(n546), .ZN(n553) );
  INV_X1 U639 ( .A(n547), .ZN(n552) );
  INV_X1 U640 ( .A(n548), .ZN(n549) );
  AND2_X1 U641 ( .A1(n550), .A2(n549), .ZN(n602) );
  NAND2_X1 U642 ( .A1(n602), .A2(n401), .ZN(n551) );
  NAND2_X1 U643 ( .A1(n553), .A2(n364), .ZN(n554) );
  NOR2_X1 U644 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U645 ( .A(n556), .B(KEYINPUT72), .ZN(n566) );
  INV_X1 U646 ( .A(n665), .ZN(n662) );
  XNOR2_X1 U647 ( .A(KEYINPUT107), .B(KEYINPUT6), .ZN(n558) );
  XNOR2_X1 U648 ( .A(n679), .B(n558), .ZN(n608) );
  NAND2_X1 U649 ( .A1(n608), .A2(n559), .ZN(n560) );
  XNOR2_X1 U650 ( .A(n560), .B(KEYINPUT111), .ZN(n561) );
  NAND2_X1 U651 ( .A1(n561), .A2(n691), .ZN(n562) );
  OR2_X1 U652 ( .A1(n662), .A2(n562), .ZN(n569) );
  NOR2_X1 U653 ( .A1(n569), .A2(n573), .ZN(n563) );
  XNOR2_X1 U654 ( .A(n563), .B(KEYINPUT36), .ZN(n565) );
  XNOR2_X1 U655 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n564) );
  XNOR2_X1 U656 ( .A(n681), .B(KEYINPUT91), .ZN(n610) );
  NAND2_X1 U657 ( .A1(n565), .A2(n610), .ZN(n672) );
  NOR2_X1 U658 ( .A1(n569), .A2(n605), .ZN(n572) );
  INV_X1 U659 ( .A(KEYINPUT112), .ZN(n570) );
  XNOR2_X1 U660 ( .A(n570), .B(KEYINPUT43), .ZN(n571) );
  XNOR2_X1 U661 ( .A(n572), .B(n571), .ZN(n574) );
  NAND2_X1 U662 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U663 ( .A(n575), .B(KEYINPUT113), .ZN(n751) );
  INV_X1 U664 ( .A(n751), .ZN(n621) );
  NAND2_X1 U665 ( .A1(n576), .A2(n668), .ZN(n673) );
  NAND2_X1 U666 ( .A1(n673), .A2(KEYINPUT2), .ZN(n577) );
  XNOR2_X1 U667 ( .A(n577), .B(KEYINPUT79), .ZN(n578) );
  NAND2_X1 U668 ( .A1(n621), .A2(n578), .ZN(n579) );
  NOR2_X1 U669 ( .A1(n623), .A2(n579), .ZN(n617) );
  INV_X1 U670 ( .A(n679), .ZN(n581) );
  OR2_X1 U671 ( .A1(n582), .A2(G898), .ZN(n584) );
  NAND2_X1 U672 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U673 ( .A(KEYINPUT0), .ZN(n587) );
  INV_X1 U674 ( .A(n592), .ZN(n598) );
  NOR2_X1 U675 ( .A1(n588), .A2(n679), .ZN(n589) );
  NOR2_X1 U676 ( .A1(n598), .A2(n590), .ZN(n652) );
  NOR2_X1 U677 ( .A1(n669), .A2(n652), .ZN(n591) );
  NOR2_X1 U678 ( .A1(n694), .A2(n675), .ZN(n593) );
  NAND2_X1 U679 ( .A1(n593), .A2(n592), .ZN(n594) );
  INV_X1 U680 ( .A(n607), .ZN(n676) );
  NOR2_X1 U681 ( .A1(n608), .A2(n676), .ZN(n595) );
  INV_X1 U682 ( .A(n596), .ZN(n650) );
  INV_X1 U683 ( .A(KEYINPUT34), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n602), .B(KEYINPUT76), .ZN(n603) );
  INV_X1 U685 ( .A(n614), .ZN(n638) );
  NOR2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n611), .B(KEYINPUT32), .ZN(n754) );
  NAND2_X1 U688 ( .A1(n614), .A2(KEYINPUT89), .ZN(n612) );
  NOR2_X1 U689 ( .A1(KEYINPUT44), .A2(KEYINPUT89), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n616) );
  INV_X1 U691 ( .A(n625), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U693 ( .A(n620), .B(KEYINPUT83), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n621), .A2(n673), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n624), .A2(n744), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n625), .B(KEYINPUT85), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n709), .A2(G472), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT62), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n634) );
  INV_X1 U702 ( .A(G952), .ZN(n633) );
  AND2_X1 U703 ( .A1(n633), .A2(G953), .ZN(n728) );
  NOR2_X2 U704 ( .A1(n634), .A2(n728), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(G57) );
  XNOR2_X1 U706 ( .A(n637), .B(G110), .ZN(G12) );
  XNOR2_X1 U707 ( .A(n638), .B(n639), .ZN(G24) );
  NAND2_X1 U708 ( .A1(n724), .A2(G217), .ZN(n641) );
  XNOR2_X1 U709 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X1 U710 ( .A1(n642), .A2(n728), .ZN(G66) );
  XOR2_X1 U711 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n643) );
  XNOR2_X1 U712 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U713 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X2 U714 ( .A1(n647), .A2(n728), .ZN(n649) );
  XNOR2_X1 U715 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n648) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(G60) );
  XOR2_X1 U717 ( .A(G101), .B(n650), .Z(G3) );
  NAND2_X1 U718 ( .A1(n652), .A2(n665), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n651), .B(G104), .ZN(G6) );
  XOR2_X1 U720 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n654) );
  NAND2_X1 U721 ( .A1(n652), .A2(n668), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U723 ( .A(G107), .B(n655), .ZN(G9) );
  INV_X1 U724 ( .A(n668), .ZN(n657) );
  NOR2_X1 U725 ( .A1(n656), .A2(n657), .ZN(n659) );
  XNOR2_X1 U726 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(n660) );
  XOR2_X1 U728 ( .A(G128), .B(n660), .Z(G30) );
  XOR2_X1 U729 ( .A(G143), .B(n661), .Z(G45) );
  NOR2_X1 U730 ( .A1(n662), .A2(n656), .ZN(n663) );
  XOR2_X1 U731 ( .A(KEYINPUT116), .B(n663), .Z(n664) );
  XNOR2_X1 U732 ( .A(G146), .B(n664), .ZN(G48) );
  XOR2_X1 U733 ( .A(G113), .B(KEYINPUT117), .Z(n667) );
  NAND2_X1 U734 ( .A1(n669), .A2(n665), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n667), .B(n666), .ZN(G15) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(G116), .ZN(G18) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(G27) );
  XNOR2_X1 U740 ( .A(G134), .B(n673), .ZN(G36) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n677), .B(KEYINPUT49), .ZN(n678) );
  NOR2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U744 ( .A(KEYINPUT118), .B(n680), .Z(n685) );
  NAND2_X1 U745 ( .A1(n681), .A2(n588), .ZN(n682) );
  XNOR2_X1 U746 ( .A(n682), .B(KEYINPUT119), .ZN(n683) );
  XNOR2_X1 U747 ( .A(KEYINPUT50), .B(n683), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n687) );
  XOR2_X1 U749 ( .A(KEYINPUT120), .B(n361), .Z(n688) );
  XNOR2_X1 U750 ( .A(n688), .B(KEYINPUT51), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n704), .A2(n689), .ZN(n690) );
  XOR2_X1 U752 ( .A(KEYINPUT121), .B(n690), .Z(n700) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U754 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U755 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U756 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U757 ( .A1(n700), .A2(n365), .ZN(n701) );
  XNOR2_X1 U758 ( .A(n701), .B(KEYINPUT52), .ZN(n702) );
  NOR2_X1 U759 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n704), .A2(n403), .ZN(n705) );
  NOR2_X1 U761 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n708), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U763 ( .A1(n709), .A2(G210), .ZN(n714) );
  XOR2_X1 U764 ( .A(KEYINPUT80), .B(KEYINPUT90), .Z(n711) );
  XNOR2_X1 U765 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n710) );
  XNOR2_X1 U766 ( .A(n711), .B(n710), .ZN(n713) );
  XNOR2_X1 U767 ( .A(n714), .B(n373), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n724), .A2(G469), .ZN(n722) );
  XOR2_X1 U769 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n719) );
  XNOR2_X1 U770 ( .A(n719), .B(KEYINPUT122), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n718), .B(n720), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U773 ( .A1(n728), .A2(n723), .ZN(G54) );
  NAND2_X1 U774 ( .A1(n724), .A2(G478), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U776 ( .A1(n728), .A2(n727), .ZN(G63) );
  NAND2_X1 U777 ( .A1(n729), .A2(n496), .ZN(n733) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n731), .A2(G898), .ZN(n732) );
  NAND2_X1 U781 ( .A1(n733), .A2(n732), .ZN(n739) );
  XOR2_X1 U782 ( .A(G110), .B(n734), .Z(n736) );
  NOR2_X1 U783 ( .A1(G898), .A2(n496), .ZN(n735) );
  NOR2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U785 ( .A(KEYINPUT125), .B(n737), .Z(n738) );
  XNOR2_X1 U786 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U787 ( .A(KEYINPUT126), .B(n740), .ZN(G69) );
  XNOR2_X1 U788 ( .A(n741), .B(KEYINPUT127), .ZN(n742) );
  XNOR2_X1 U789 ( .A(n743), .B(n742), .ZN(n746) );
  XNOR2_X1 U790 ( .A(n744), .B(n746), .ZN(n745) );
  NAND2_X1 U791 ( .A1(n745), .A2(n496), .ZN(n750) );
  XOR2_X1 U792 ( .A(G227), .B(n746), .Z(n747) );
  NAND2_X1 U793 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U794 ( .A1(G953), .A2(n748), .ZN(n749) );
  NAND2_X1 U795 ( .A1(n750), .A2(n749), .ZN(G72) );
  XOR2_X1 U796 ( .A(G140), .B(n751), .Z(G42) );
  XOR2_X1 U797 ( .A(G131), .B(n752), .Z(G33) );
  XOR2_X1 U798 ( .A(G137), .B(n753), .Z(G39) );
  XNOR2_X1 U799 ( .A(G119), .B(n754), .ZN(G21) );
endmodule

