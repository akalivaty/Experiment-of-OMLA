//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(KEYINPUT14), .B(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n205), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT96), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n204), .A2(KEYINPUT15), .A3(new_n208), .A4(new_n206), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT95), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT17), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n218), .ZN(new_n221));
  XOR2_X1   g020(.A(new_n221), .B(G8gat), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n222), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n223), .A2(KEYINPUT18), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n216), .B(new_n225), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n224), .B(KEYINPUT13), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n216), .B(new_n232), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n224), .B(new_n226), .C1(new_n233), .C2(new_n225), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT97), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n223), .A2(KEYINPUT97), .A3(new_n224), .A4(new_n226), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT98), .B(KEYINPUT18), .Z(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G113gat), .B(G141gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT94), .ZN(new_n241));
  XOR2_X1   g040(.A(G169gat), .B(G197gat), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(new_n245), .B(KEYINPUT12), .Z(new_n246));
  AND3_X1   g045(.A1(new_n231), .A2(new_n239), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n231), .B2(new_n239), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT99), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n239), .ZN(new_n250));
  INV_X1    g049(.A(new_n246), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT99), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n239), .A3(new_n246), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259));
  XNOR2_X1  g058(.A(G141gat), .B(G148gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G155gat), .ZN(new_n262));
  INV_X1    g061(.A(G162gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(KEYINPUT2), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n265), .B(new_n264), .C1(new_n260), .C2(KEYINPUT2), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n259), .B1(new_n270), .B2(KEYINPUT3), .ZN(new_n271));
  XNOR2_X1  g070(.A(G197gat), .B(G204gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT22), .ZN(new_n273));
  INV_X1    g072(.A(G211gat), .ZN(new_n274));
  INV_X1    g073(.A(G218gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G211gat), .B(G218gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n272), .A3(new_n276), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n271), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G228gat), .ZN(new_n285));
  INV_X1    g084(.A(G233gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT29), .B1(new_n280), .B2(new_n281), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n270), .B1(new_n288), .B2(KEYINPUT3), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT3), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n288), .B2(new_n291), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n270), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n284), .A2(KEYINPUT86), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT86), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n271), .A2(new_n297), .A3(new_n283), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n287), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n299), .A2(KEYINPUT87), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT87), .B1(new_n299), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n290), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G22gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305));
  INV_X1    g104(.A(G50gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G22gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n309), .B(new_n290), .C1(new_n301), .C2(new_n302), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n304), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n308), .B1(new_n304), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n258), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n313), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(new_n257), .A3(new_n311), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  NOR2_X1   g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G169gat), .ZN(new_n320));
  INV_X1    g119(.A(G176gat), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT23), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(KEYINPUT23), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n319), .A2(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT24), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G183gat), .B(G190gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(new_n329), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT64), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n325), .B(new_n326), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n332), .A2(new_n333), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n317), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n322), .A2(new_n319), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(KEYINPUT25), .A3(new_n323), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n338), .A2(new_n332), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n320), .A2(new_n321), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n341), .A2(KEYINPUT26), .A3(new_n318), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n318), .A2(KEYINPUT26), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n342), .A2(new_n328), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G183gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(KEYINPUT27), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(G190gat), .B1(new_n345), .B2(KEYINPUT27), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(KEYINPUT28), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n345), .B2(KEYINPUT27), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n352), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT67), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT67), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n355), .A2(new_n359), .A3(new_n356), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n350), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n344), .B1(new_n361), .B2(KEYINPUT68), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n355), .A2(new_n359), .A3(new_n356), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n359), .B1(new_n355), .B2(new_n356), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT68), .B(new_n349), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n340), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n368));
  INV_X1    g167(.A(G134gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G127gat), .ZN(new_n370));
  INV_X1    g169(.A(G127gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G134gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT1), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G113gat), .ZN(new_n375));
  INV_X1    g174(.A(G120gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G113gat), .A2(G120gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n368), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n378), .ZN(new_n381));
  NOR2_X1   g180(.A1(G113gat), .A2(G120gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G127gat), .B(G134gat), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT70), .A4(new_n373), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT69), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n381), .B2(new_n382), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(KEYINPUT69), .A3(new_n378), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n373), .ZN(new_n389));
  INV_X1    g188(.A(new_n384), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n380), .A2(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n367), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G227gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n286), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n349), .B1(new_n363), .B2(new_n364), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT68), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n365), .A3(new_n344), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n385), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n390), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n398), .A2(new_n401), .A3(new_n340), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n392), .A2(new_n394), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404));
  XOR2_X1   g203(.A(G15gat), .B(G43gat), .Z(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT71), .ZN(new_n406));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n403), .B(KEYINPUT32), .C1(new_n404), .C2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n411));
  INV_X1    g210(.A(new_n408), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n398), .A2(new_n401), .A3(new_n340), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n401), .B1(new_n398), .B2(new_n340), .ZN(new_n414));
  INV_X1    g213(.A(new_n394), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT32), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n416), .A2(KEYINPUT33), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n411), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n408), .B1(new_n403), .B2(KEYINPUT32), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n404), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT72), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n410), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n415), .B1(new_n413), .B2(new_n414), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT34), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT34), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n427), .B(new_n415), .C1(new_n413), .C2(new_n414), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n314), .A2(new_n316), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n426), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n426), .B2(new_n428), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT73), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n424), .B2(new_n438), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT73), .B(new_n410), .C1(new_n420), .C2(new_n423), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n439), .A2(KEYINPUT75), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT75), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n421), .A2(KEYINPUT72), .A3(new_n422), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT72), .B1(new_n421), .B2(new_n422), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n409), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n436), .B1(new_n445), .B2(KEYINPUT73), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n438), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n442), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n432), .B1(new_n441), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  INV_X1    g250(.A(G226gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(new_n286), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n344), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n395), .B2(new_n396), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n456), .A2(new_n365), .B1(new_n336), .B2(new_n339), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n454), .B1(new_n457), .B2(KEYINPUT29), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n457), .A2(KEYINPUT78), .A3(new_n454), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT78), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n367), .B2(new_n453), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n282), .B(new_n458), .C1(new_n459), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n367), .A2(new_n453), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n283), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(G8gat), .B(G36gat), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT79), .ZN(new_n468));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  AOI21_X1  g269(.A(new_n451), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n282), .B1(new_n458), .B2(new_n463), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n453), .B1(new_n367), .B2(new_n259), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n463), .A2(KEYINPUT78), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n367), .A2(new_n460), .A3(new_n453), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n476), .B2(new_n282), .ZN(new_n477));
  INV_X1    g276(.A(new_n470), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n451), .A3(new_n478), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n270), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n391), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n391), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G225gat), .A2(G233gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT80), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n399), .A2(new_n400), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n399), .B2(new_n400), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n268), .A2(new_n269), .A3(new_n293), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n293), .B1(new_n268), .B2(new_n269), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n493), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT5), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n491), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n401), .A2(KEYINPUT80), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n391), .A2(new_n494), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n401), .A2(new_n270), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n484), .A2(new_n487), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n506), .A2(new_n508), .A3(new_n492), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT82), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n488), .B1(new_n391), .B2(new_n483), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(KEYINPUT4), .B2(new_n507), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n501), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n504), .A2(new_n505), .A3(new_n270), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n484), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n502), .B1(new_n518), .B2(new_n493), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n503), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G1gat), .B(G29gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT0), .ZN(new_n522));
  XNOR2_X1  g321(.A(G57gat), .B(G85gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n522), .B(new_n523), .Z(new_n524));
  NOR2_X1   g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT6), .ZN(new_n526));
  INV_X1    g325(.A(new_n524), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n507), .B1(new_n497), .B2(new_n270), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT5), .B1(new_n528), .B2(new_n492), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n511), .B2(new_n515), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n527), .B1(new_n530), .B2(new_n503), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n519), .ZN(new_n532));
  INV_X1    g331(.A(new_n503), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n524), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n526), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n450), .B1(new_n482), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n482), .A2(new_n450), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT35), .B1(new_n449), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n535), .B1(new_n520), .B2(new_n524), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n530), .A2(new_n527), .A3(new_n503), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n531), .A2(new_n534), .A3(KEYINPUT90), .A4(new_n535), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n526), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n482), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT92), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT35), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n314), .A2(new_n316), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n445), .A2(new_n429), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n431), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n542), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n540), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n552), .B1(new_n558), .B2(new_n538), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n464), .B2(new_n282), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n283), .B(new_n458), .C1(new_n459), .C2(new_n461), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT38), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n462), .A2(new_n465), .A3(new_n560), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n470), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n479), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT91), .B1(new_n548), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n547), .A2(new_n526), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n466), .A2(new_n470), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n564), .A2(new_n470), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(new_n563), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n568), .A2(new_n571), .A3(new_n572), .A4(new_n546), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n560), .B2(new_n477), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT38), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n567), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT40), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n492), .B1(new_n491), .B2(new_n506), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n517), .A2(new_n492), .A3(new_n484), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(KEYINPUT39), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n579), .A3(KEYINPUT39), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n506), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n493), .B1(new_n585), .B2(new_n490), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n524), .B1(new_n586), .B2(KEYINPUT39), .ZN(new_n587));
  OAI211_X1 g386(.A(KEYINPUT89), .B(new_n577), .C1(new_n584), .C2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT89), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n582), .B2(new_n583), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(KEYINPUT40), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n525), .B1(KEYINPUT40), .B2(new_n590), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n592), .A2(new_n480), .A3(new_n481), .A4(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n594), .A2(new_n316), .A3(new_n314), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n576), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n420), .A2(new_n423), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n430), .B1(new_n599), .B2(new_n409), .ZN(new_n600));
  AOI211_X1 g399(.A(new_n429), .B(new_n410), .C1(new_n420), .C2(new_n423), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT77), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT77), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n554), .A2(new_n604), .A3(new_n598), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n431), .A2(KEYINPUT36), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT75), .B1(new_n439), .B2(new_n440), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n446), .A2(new_n442), .A3(new_n447), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n559), .B(new_n596), .C1(new_n606), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n256), .B1(new_n557), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT101), .ZN(new_n614));
  NOR2_X1   g413(.A1(G71gat), .A2(G78gat), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n615), .A2(KEYINPUT100), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n614), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G57gat), .B(G64gat), .Z(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(KEYINPUT9), .B2(new_n613), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OR3_X1    g419(.A1(new_n619), .A2(new_n613), .A3(new_n615), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(KEYINPUT21), .ZN(new_n623));
  AND2_X1   g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G127gat), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n225), .B1(KEYINPUT21), .B2(new_n622), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G155gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT7), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(G85gat), .B2(G92gat), .ZN(new_n637));
  OAI211_X1 g436(.A(G85gat), .B(G92gat), .C1(new_n636), .C2(KEYINPUT102), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n636), .A2(KEYINPUT102), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n640), .B2(KEYINPUT103), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(KEYINPUT103), .B2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  INV_X1    g442(.A(G85gat), .ZN(new_n644));
  INV_X1    g443(.A(G92gat), .ZN(new_n645));
  AOI22_X1  g444(.A1(KEYINPUT8), .A2(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G99gat), .B(G106gat), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n650), .A3(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n217), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n649), .A2(new_n651), .ZN(new_n654));
  AND2_X1   g453(.A1(G232gat), .A2(G233gat), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n654), .A2(new_n216), .B1(KEYINPUT41), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G190gat), .B(G218gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n655), .A2(KEYINPUT41), .ZN(new_n660));
  XNOR2_X1  g459(.A(G134gat), .B(G162gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n658), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n653), .A2(new_n663), .A3(new_n656), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n659), .B2(new_n664), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n635), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n622), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n652), .A2(new_n620), .A3(new_n621), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n654), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(G230gat), .A2(G233gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n671), .ZN(new_n678));
  INV_X1    g477(.A(new_n676), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G120gat), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(G176gat), .B(G204gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n677), .A2(new_n680), .A3(new_n684), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n669), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n612), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n537), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g491(.A1(new_n690), .A2(new_n482), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(G8gat), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT16), .B(G8gat), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(new_n694), .B2(new_n695), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n696), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(G1325gat));
  NAND2_X1  g502(.A1(new_n608), .A2(new_n609), .ZN(new_n704));
  INV_X1    g503(.A(new_n607), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n704), .A2(new_n705), .B1(new_n603), .B2(new_n605), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n690), .B2(new_n707), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n554), .A2(G15gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n690), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT106), .ZN(G1326gat));
  NAND3_X1  g510(.A1(new_n612), .A2(new_n552), .A3(new_n689), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT107), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT43), .B(G22gat), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n713), .B(new_n714), .Z(G1327gat));
  NOR3_X1   g514(.A1(new_n635), .A2(new_n668), .A3(new_n688), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n612), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(G29gat), .A3(new_n537), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT45), .Z(new_n719));
  INV_X1    g518(.A(KEYINPUT92), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n549), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n555), .A2(new_n551), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n314), .A2(new_n316), .A3(new_n431), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n608), .B2(new_n609), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n558), .A2(new_n538), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n551), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n596), .A2(new_n559), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n723), .A2(new_n727), .B1(new_n728), .B2(new_n706), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n667), .B(KEYINPUT108), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n668), .B1(new_n557), .B2(new_n611), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n730), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n635), .A2(new_n688), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n252), .A2(new_n254), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n537), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n719), .B1(new_n205), .B2(new_n740), .ZN(G1328gat));
  NOR3_X1   g540(.A1(new_n717), .A2(G36gat), .A3(new_n482), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT46), .ZN(new_n743));
  INV_X1    g542(.A(new_n482), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n745), .B2(new_n203), .ZN(G1329gat));
  NAND3_X1  g545(.A1(new_n734), .A2(new_n706), .A3(new_n737), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G43gat), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT47), .B1(new_n748), .B2(KEYINPUT109), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n554), .A2(G43gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n717), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n749), .B(new_n751), .ZN(G1330gat));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n552), .A3(new_n737), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G50gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n612), .A2(new_n306), .A3(new_n552), .A4(new_n716), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(KEYINPUT48), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT111), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n754), .A2(KEYINPUT111), .A3(new_n756), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n755), .B(KEYINPUT110), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(G50gat), .B2(new_n753), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n757), .A2(new_n758), .B1(new_n760), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI211_X1 g560(.A(new_n736), .B(new_n669), .C1(new_n557), .C2(new_n611), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n688), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n739), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  INV_X1    g565(.A(new_n688), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n482), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT49), .B(G64gat), .Z(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n763), .B2(new_n707), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n554), .A2(G71gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n763), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1334gat));
  NAND2_X1  g576(.A1(new_n764), .A2(new_n552), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT113), .B(G78gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n635), .A2(new_n736), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n767), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n734), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n537), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(KEYINPUT114), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n733), .B2(new_n781), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AND4_X1   g589(.A1(new_n729), .A2(new_n667), .A3(new_n781), .A4(new_n790), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n739), .A2(new_n644), .A3(new_n688), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n785), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  NOR3_X1   g594(.A1(new_n482), .A2(new_n767), .A3(G92gat), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n783), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n730), .B1(new_n729), .B2(new_n667), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n800), .B2(new_n732), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n645), .B1(new_n801), .B2(new_n744), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n784), .A2(new_n805), .A3(new_n482), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT115), .B1(new_n801), .B2(new_n744), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(new_n645), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n804), .B2(new_n808), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n784), .B2(new_n707), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n554), .A2(G99gat), .A3(new_n767), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n793), .B2(new_n811), .ZN(G1338gat));
  INV_X1    g611(.A(G106gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n552), .A2(new_n813), .A3(new_n688), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n788), .B2(new_n791), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n734), .A2(KEYINPUT116), .A3(new_n552), .A4(new_n783), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n731), .A2(new_n730), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n557), .B2(new_n611), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n552), .B(new_n783), .C1(new_n799), .C2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n813), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n818), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(G106gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n817), .B1(new_n826), .B2(new_n816), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n822), .A2(new_n823), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n819), .A3(G106gat), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n816), .A2(new_n817), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n826), .A2(new_n816), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n828), .A2(new_n836), .ZN(G1339gat));
  NAND3_X1  g636(.A1(new_n673), .A2(new_n674), .A3(new_n679), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n677), .A2(KEYINPUT54), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n679), .B1(new_n673), .B2(new_n674), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n684), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n687), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n839), .A2(new_n842), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n844), .B(new_n847), .C1(new_n247), .C2(new_n248), .ZN(new_n848));
  INV_X1    g647(.A(new_n245), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n224), .B1(new_n223), .B2(new_n226), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n228), .A2(new_n229), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n254), .A2(new_n688), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT118), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n254), .A2(new_n688), .A3(new_n855), .A4(new_n852), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n848), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT119), .ZN(new_n858));
  INV_X1    g657(.A(new_n731), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n848), .A2(new_n854), .A3(new_n860), .A4(new_n856), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n847), .A2(new_n687), .A3(new_n843), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n254), .A2(new_n852), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n731), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n635), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n669), .A2(new_n736), .A3(new_n688), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(new_n739), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n482), .A3(new_n725), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n375), .B(new_n736), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n868), .A2(new_n555), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n744), .A2(new_n537), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n256), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n874), .A2(new_n878), .ZN(G1340gat));
  OAI211_X1 g678(.A(new_n376), .B(new_n688), .C1(new_n872), .C2(new_n873), .ZN(new_n880));
  OAI21_X1  g679(.A(G120gat), .B1(new_n877), .B2(new_n767), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1341gat));
  INV_X1    g681(.A(new_n635), .ZN(new_n883));
  OAI21_X1  g682(.A(G127gat), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n635), .A2(new_n371), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n870), .B2(new_n885), .ZN(G1342gat));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n725), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n668), .A2(new_n744), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n369), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n887), .A2(KEYINPUT56), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT56), .B1(new_n887), .B2(new_n889), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n667), .A3(new_n876), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(G134gat), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n892), .B2(G134gat), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n890), .B(new_n891), .C1(new_n894), .C2(new_n895), .ZN(G1343gat));
  NAND2_X1  g695(.A1(new_n707), .A2(new_n876), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  XOR2_X1   g697(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n868), .B2(new_n552), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n552), .A2(KEYINPUT57), .ZN(new_n902));
  INV_X1    g701(.A(new_n865), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n249), .A2(new_n255), .A3(new_n863), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n667), .B1(new_n904), .B2(new_n853), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n883), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n867), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n898), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G141gat), .B1(new_n909), .B2(new_n256), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n707), .A2(new_n552), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AND4_X1   g711(.A1(new_n739), .A2(new_n868), .A3(new_n482), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n256), .A2(G141gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT58), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n736), .B(new_n898), .C1(new_n901), .C2(new_n908), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n918), .A2(G141gat), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(G148gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n913), .A2(new_n921), .A3(new_n688), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n844), .A2(new_n667), .A3(new_n847), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n863), .A2(new_n926), .A3(new_n667), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n925), .A2(new_n927), .A3(new_n864), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n883), .B1(new_n928), .B2(new_n905), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n689), .A2(new_n256), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n552), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n552), .B(new_n900), .C1(new_n866), .C2(new_n867), .ZN(new_n935));
  AOI211_X1 g734(.A(new_n767), .B(new_n897), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n921), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n935), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n688), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT124), .B1(new_n940), .B2(new_n897), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n923), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n909), .A2(new_n767), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n923), .A2(G148gat), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n922), .B1(new_n942), .B2(new_n945), .ZN(G1345gat));
  OAI21_X1  g745(.A(G155gat), .B1(new_n909), .B2(new_n883), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n913), .A2(new_n262), .A3(new_n635), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1346gat));
  OAI21_X1  g748(.A(G162gat), .B1(new_n909), .B2(new_n859), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n869), .A2(new_n263), .A3(new_n888), .A4(new_n912), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1347gat));
  NOR2_X1   g751(.A1(new_n482), .A2(new_n739), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n875), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n954), .A2(new_n320), .A3(new_n256), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n868), .A2(new_n537), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n449), .A2(new_n482), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n736), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n955), .B1(new_n320), .B2(new_n958), .ZN(G1348gat));
  NOR3_X1   g758(.A1(new_n954), .A2(new_n321), .A3(new_n767), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n956), .A2(new_n957), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n321), .B1(new_n961), .B2(new_n767), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g763(.A(KEYINPUT125), .B(new_n321), .C1(new_n961), .C2(new_n767), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(G1349gat));
  OAI21_X1  g765(.A(G183gat), .B1(new_n954), .B2(new_n883), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n353), .A2(G183gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n883), .A2(new_n346), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n956), .A2(new_n957), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT60), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n967), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1350gat));
  OR3_X1    g774(.A1(new_n961), .A2(G190gat), .A3(new_n859), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n868), .A2(new_n555), .A3(new_n667), .A4(new_n953), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G190gat), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(KEYINPUT126), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n981), .A3(G190gat), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n980), .B1(new_n979), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n976), .B1(new_n983), .B2(new_n984), .ZN(G1351gat));
  NAND2_X1  g784(.A1(new_n956), .A2(new_n912), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n986), .A2(new_n482), .ZN(new_n987));
  AOI21_X1  g786(.A(G197gat), .B1(new_n987), .B2(new_n736), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n707), .A2(new_n953), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n989), .B1(new_n934), .B2(new_n935), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n249), .A2(new_n255), .A3(G197gat), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(G1352gat));
  XNOR2_X1  g791(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n993));
  INV_X1    g792(.A(G204gat), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n768), .A2(new_n994), .ZN(new_n995));
  OR3_X1    g794(.A1(new_n986), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(G204gat), .B1(new_n940), .B2(new_n989), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n993), .B1(new_n986), .B2(new_n995), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(G1353gat));
  NAND3_X1  g798(.A1(new_n987), .A2(new_n274), .A3(new_n635), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n990), .A2(new_n635), .ZN(new_n1001));
  AND3_X1   g800(.A1(new_n1001), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(KEYINPUT63), .B1(new_n1001), .B2(G211gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(G1354gat));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n275), .A3(new_n731), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n990), .A2(new_n667), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1005), .B1(new_n275), .B2(new_n1006), .ZN(G1355gat));
endmodule


