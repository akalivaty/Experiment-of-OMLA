//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT65), .B(G77), .Z(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G87), .A2(G250), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  INV_X1    g0026(.A(G13), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n226), .B1(new_n208), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n209), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n214), .B(new_n225), .C1(new_n231), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n240), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n209), .A2(G33), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT70), .Z(new_n256));
  INV_X1    g0056(.A(G58), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(KEYINPUT8), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT69), .B(G58), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(KEYINPUT8), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n254), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n210), .A2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n230), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n227), .A2(new_n209), .A3(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n202), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n230), .A2(new_n262), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G1), .B2(new_n209), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n264), .B(new_n266), .C1(new_n202), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT73), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT72), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n275), .ZN(new_n282));
  INV_X1    g0082(.A(G226), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n278), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n228), .B(new_n229), .C1(new_n279), .C2(new_n280), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n285), .B1(new_n216), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n287), .A2(new_n288), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT68), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(G223), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(G223), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G222), .A2(G1698), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n291), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n284), .B1(new_n290), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(G190), .B2(new_n299), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n272), .A2(new_n274), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT10), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n269), .B1(G169), .B2(new_n299), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n260), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(new_n265), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n268), .B2(new_n311), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n314));
  OR2_X1    g0114(.A1(KEYINPUT74), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT74), .A2(G33), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n286), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n317), .A2(new_n318), .B1(KEYINPUT3), .B2(new_n279), .ZN(new_n319));
  AND2_X1   g0119(.A1(KEYINPUT74), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(KEYINPUT74), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT75), .A3(new_n286), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n314), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT7), .B1(new_n289), .B2(new_n209), .ZN(new_n325));
  OAI21_X1  g0125(.A(G68), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G68), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n232), .B1(new_n259), .B2(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(G20), .B1(G159), .B2(new_n253), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT3), .B1(new_n320), .B2(new_n321), .ZN(new_n333));
  AOI21_X1  g0133(.A(G20), .B1(new_n333), .B2(new_n287), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  OAI21_X1  g0135(.A(G68), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n287), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n315), .A2(new_n316), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(KEYINPUT3), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n339), .A2(KEYINPUT7), .A3(G20), .ZN(new_n340));
  OAI211_X1 g0140(.A(KEYINPUT16), .B(new_n329), .C1(new_n336), .C2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n341), .A2(new_n263), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n313), .B1(new_n332), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NOR2_X1   g0144(.A1(G223), .A2(G1698), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n283), .B2(G1698), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(new_n333), .A3(new_n287), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G87), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n285), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G232), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n278), .B1(new_n282), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n300), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n349), .A2(new_n354), .A3(new_n351), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n343), .A2(new_n344), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n313), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT16), .B1(new_n326), .B2(new_n329), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n341), .A2(new_n263), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n356), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT17), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n352), .A2(G179), .ZN(new_n364));
  OAI21_X1  g0164(.A(G169), .B1(new_n349), .B2(new_n351), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT76), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n358), .B(KEYINPUT76), .C1(new_n359), .C2(new_n360), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n363), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AOI211_X1 g0175(.A(KEYINPUT18), .B(new_n367), .C1(new_n370), .C2(new_n371), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n265), .A2(new_n327), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT12), .ZN(new_n380));
  INV_X1    g0180(.A(G77), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n256), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n253), .A2(G50), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n209), .B2(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n263), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT11), .ZN(new_n386));
  OAI221_X1 g0186(.A(new_n380), .B1(new_n327), .B2(new_n268), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n385), .A2(new_n386), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n281), .A2(G238), .A3(new_n275), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n350), .A2(G1698), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n291), .B(new_n392), .C1(G226), .C2(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n278), .B(new_n391), .C1(new_n395), .C2(new_n285), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(KEYINPUT13), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G179), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  INV_X1    g0201(.A(G169), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n397), .B2(new_n398), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n400), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n403), .A2(new_n401), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n390), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n390), .B1(new_n399), .B2(G190), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n300), .B2(new_n399), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n268), .A2(new_n381), .ZN(new_n410));
  XOR2_X1   g0210(.A(new_n410), .B(KEYINPUT71), .Z(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT8), .B(G58), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n253), .B1(new_n215), .B2(G20), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n255), .B2(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(new_n263), .B1(new_n216), .B2(new_n265), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n285), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G232), .A2(G1698), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n292), .A2(G238), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n291), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n419), .B(new_n422), .C1(G107), .C2(new_n291), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n282), .A2(new_n217), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n277), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n402), .ZN(new_n427));
  INV_X1    g0227(.A(new_n426), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n306), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n418), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n426), .A2(new_n354), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(G200), .B2(new_n426), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(new_n411), .A3(new_n417), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NOR4_X1   g0234(.A1(new_n310), .A2(new_n378), .A3(new_n409), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT80), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G283), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n292), .B1(KEYINPUT4), .B2(G244), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT4), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n333), .A2(new_n439), .A3(new_n287), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n440), .B2(G244), .ZN(new_n441));
  INV_X1    g0241(.A(G250), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G1698), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n439), .B1(new_n291), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n437), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT78), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(KEYINPUT78), .B(new_n437), .C1(new_n441), .C2(new_n444), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n419), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT79), .B1(new_n450), .B2(G41), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT79), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n280), .A3(KEYINPUT5), .ZN(new_n453));
  INV_X1    g0253(.A(G45), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G1), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(G41), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n451), .A2(new_n453), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n276), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n281), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n460), .B2(G257), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n449), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n436), .B1(new_n462), .B2(G179), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n265), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n265), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(G1), .B2(new_n279), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(new_n263), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n465), .B1(new_n469), .B2(new_n464), .ZN(new_n470));
  OAI21_X1  g0270(.A(G107), .B1(new_n324), .B2(new_n325), .ZN(new_n471));
  INV_X1    g0271(.A(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(KEYINPUT6), .A3(G97), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT77), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  XOR2_X1   g0276(.A(G97), .B(G107), .Z(new_n477));
  OAI211_X1 g0277(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(KEYINPUT6), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n470), .B1(new_n480), .B2(new_n263), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n462), .B2(new_n402), .ZN(new_n482));
  INV_X1    g0282(.A(new_n461), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n285), .B1(new_n445), .B2(new_n446), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n448), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(KEYINPUT80), .A3(new_n306), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n463), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(G190), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(new_n481), .C1(new_n300), .C2(new_n485), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT84), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n457), .A2(G270), .A3(new_n281), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT83), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n458), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n457), .A2(KEYINPUT83), .A3(G270), .A4(new_n281), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n289), .A2(G303), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n333), .A2(new_n287), .ZN(new_n499));
  INV_X1    g0299(.A(G264), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G1698), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(G257), .B2(G1698), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT85), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n285), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(KEYINPUT85), .B(new_n498), .C1(new_n499), .C2(new_n502), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n491), .A2(new_n497), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT84), .A4(new_n496), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G200), .ZN(new_n510));
  INV_X1    g0310(.A(G116), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G20), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n464), .A2(G33), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n437), .A2(new_n209), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n263), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT20), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n466), .A2(G116), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n468), .B2(G116), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n510), .B(new_n520), .C1(new_n354), .C2(new_n509), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n455), .A2(new_n442), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n281), .B1(G274), .B2(new_n455), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n338), .A2(new_n511), .ZN(new_n524));
  NOR2_X1   g0324(.A1(G238), .A2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n217), .B2(G1698), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n339), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n523), .B1(new_n527), .B2(new_n285), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G200), .ZN(new_n529));
  OAI211_X1 g0329(.A(G190), .B(new_n523), .C1(new_n527), .C2(new_n285), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n468), .A2(G87), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n209), .B1(new_n394), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g0333(.A(KEYINPUT82), .B(G87), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n206), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n255), .B2(new_n464), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n209), .A2(G68), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n536), .C1(new_n499), .C2(new_n537), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n538), .A2(new_n263), .B1(new_n265), .B2(new_n415), .ZN(new_n539));
  AND4_X1   g0339(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n539), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n527), .A2(new_n285), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n541), .A2(KEYINPUT81), .A3(new_n306), .A4(new_n523), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n539), .B1(new_n415), .B2(new_n469), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n528), .A2(new_n402), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n541), .A2(new_n306), .A3(new_n523), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT81), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n540), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  MUX2_X1   g0349(.A(G250), .B(G257), .S(G1698), .Z(new_n550));
  AOI22_X1  g0350(.A1(new_n339), .A2(new_n550), .B1(G294), .B2(new_n322), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(new_n285), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n459), .A2(new_n500), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n552), .A2(new_n458), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(KEYINPUT87), .A3(new_n354), .ZN(new_n555));
  OAI221_X1 g0355(.A(new_n495), .B1(new_n500), .B2(new_n459), .C1(new_n551), .C2(new_n285), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n300), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT87), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n556), .B2(G190), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n291), .A2(new_n209), .A3(G87), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT86), .B1(new_n472), .B2(G20), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n524), .ZN(new_n571));
  INV_X1    g0371(.A(G87), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n563), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n333), .A2(new_n287), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(G20), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n561), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n562), .A2(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n524), .B1(new_n339), .B2(new_n573), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(KEYINPUT24), .C1(new_n578), .C2(G20), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n579), .A3(new_n263), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n466), .B2(G107), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n265), .A2(KEYINPUT25), .A3(new_n472), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n468), .A2(G107), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n560), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n521), .A2(new_n549), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n517), .A2(new_n519), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n509), .A2(G169), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n497), .A2(new_n491), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n503), .A2(new_n504), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n506), .A3(new_n419), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n593), .A2(G179), .A3(new_n508), .A4(new_n595), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n520), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n509), .A2(KEYINPUT21), .A3(G169), .A4(new_n589), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n556), .A2(new_n402), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n585), .B(new_n599), .C1(G179), .C2(new_n556), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n592), .A2(new_n597), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n588), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n435), .A2(new_n490), .A3(new_n602), .ZN(G372));
  NAND2_X1  g0403(.A1(new_n368), .A2(new_n366), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n604), .B(new_n373), .ZN(new_n605));
  INV_X1    g0405(.A(new_n430), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n408), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n406), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT90), .ZN(new_n609));
  INV_X1    g0409(.A(new_n363), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n308), .B1(new_n611), .B2(new_n304), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n543), .A2(new_n546), .A3(new_n544), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT88), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n529), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n539), .A2(new_n531), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n528), .A2(KEYINPUT88), .A3(G200), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n530), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n613), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n586), .B2(new_n560), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n601), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n622), .B2(new_n490), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n463), .A2(new_n482), .A3(new_n486), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n549), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT89), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n549), .A2(new_n463), .A3(new_n482), .A4(new_n486), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n620), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(new_n463), .A3(new_n482), .A4(new_n486), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n628), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n625), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n435), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n612), .A2(new_n635), .ZN(G369));
  INV_X1    g0436(.A(KEYINPUT91), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n227), .A2(G20), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n208), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(G213), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n520), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n637), .B1(new_n638), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n638), .A2(new_n521), .A3(new_n647), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(KEYINPUT91), .A3(new_n646), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G330), .ZN(new_n653));
  INV_X1    g0453(.A(new_n645), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n600), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n645), .B1(new_n580), .B2(new_n584), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n560), .B2(new_n586), .ZN(new_n657));
  INV_X1    g0457(.A(new_n600), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n653), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n650), .A2(new_n600), .A3(new_n645), .A4(new_n657), .ZN(new_n662));
  INV_X1    g0462(.A(new_n655), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(G399));
  NOR3_X1   g0466(.A1(new_n534), .A2(G116), .A3(new_n206), .ZN(new_n667));
  XOR2_X1   g0467(.A(new_n667), .B(KEYINPUT92), .Z(new_n668));
  INV_X1    g0468(.A(new_n212), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(G1), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n233), .B2(new_n671), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n654), .B1(new_n623), .B2(new_n633), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT29), .ZN(new_n676));
  OR3_X1    g0476(.A1(new_n631), .A2(KEYINPUT95), .A3(new_n628), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n627), .A2(new_n628), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT95), .B1(new_n631), .B2(new_n628), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n654), .B1(new_n680), .B2(new_n623), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT29), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT31), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n556), .A2(new_n306), .A3(new_n528), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n462), .A2(new_n509), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT93), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n596), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n507), .A2(KEYINPUT93), .A3(G179), .A4(new_n508), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n528), .A2(new_n552), .A3(new_n553), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n449), .A2(new_n461), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n686), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n690), .A2(new_n693), .A3(KEYINPUT30), .ZN(new_n697));
  AOI211_X1 g0497(.A(new_n683), .B(new_n645), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n697), .A3(new_n685), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT31), .B1(new_n700), .B2(new_n654), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT94), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n692), .B1(new_n688), .B2(new_n689), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n685), .B1(new_n703), .B2(KEYINPUT30), .ZN(new_n704));
  INV_X1    g0504(.A(new_n697), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n654), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n683), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT94), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n602), .A2(new_n490), .A3(new_n645), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n702), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n676), .A2(new_n682), .B1(G330), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n674), .B1(new_n713), .B2(G1), .ZN(G364));
  AOI21_X1  g0514(.A(new_n208), .B1(new_n639), .B2(G45), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n670), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT96), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n652), .A2(new_n719), .A3(G330), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n719), .B1(new_n652), .B2(G330), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n718), .B1(G330), .B2(new_n652), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n230), .B1(G20), .B2(new_n402), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT97), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(KEYINPUT97), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n212), .A2(new_n291), .ZN(new_n733));
  INV_X1    g0533(.A(G355), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n733), .A2(new_n734), .B1(G116), .B2(new_n212), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n669), .A2(new_n339), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G45), .B2(new_n233), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n248), .A2(new_n454), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n717), .B1(new_n732), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n354), .A2(G20), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n300), .A2(G179), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G283), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n209), .A2(new_n354), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n306), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G322), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n745), .A2(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n742), .A2(new_n306), .A3(new_n300), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT33), .B(G317), .Z(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n743), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n751), .B(new_n755), .C1(G329), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n743), .A2(new_n748), .ZN(new_n760));
  INV_X1    g0560(.A(G311), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n306), .A2(new_n300), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n747), .ZN(new_n763));
  INV_X1    g0563(.A(G326), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n760), .A2(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n747), .A2(new_n744), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n291), .B(new_n765), .C1(G303), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G294), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n209), .B1(new_n756), .B2(G190), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n759), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n289), .B1(new_n767), .B2(new_n534), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT99), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n749), .B(KEYINPUT98), .ZN(new_n774));
  INV_X1    g0574(.A(new_n259), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n760), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n777), .A2(new_n215), .B1(new_n752), .B2(G68), .ZN(new_n778));
  INV_X1    g0578(.A(new_n763), .ZN(new_n779));
  INV_X1    g0579(.A(new_n745), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G50), .A2(new_n779), .B1(new_n780), .B2(G107), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n773), .A2(new_n776), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  OR3_X1    g0583(.A1(new_n757), .A2(KEYINPUT32), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(KEYINPUT32), .B1(new_n757), .B2(new_n783), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n464), .C2(new_n770), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n771), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n741), .B1(new_n787), .B2(new_n727), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n730), .B(KEYINPUT100), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n652), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n723), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  INV_X1    g0592(.A(new_n727), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n729), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n717), .B1(new_n794), .B2(G77), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n430), .A2(new_n654), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n418), .A2(new_n654), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n798), .A2(new_n433), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n797), .B1(new_n799), .B2(new_n606), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n729), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n753), .A2(new_n746), .B1(new_n472), .B2(new_n766), .ZN(new_n803));
  INV_X1    g0603(.A(new_n749), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n291), .B(new_n803), .C1(G294), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n745), .A2(new_n572), .ZN(new_n806));
  INV_X1    g0606(.A(G303), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n760), .A2(new_n511), .B1(new_n763), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(G311), .C2(new_n758), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n805), .B(new_n809), .C1(new_n464), .C2(new_n770), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n780), .A2(G68), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n811), .B1(new_n202), .B2(new_n766), .C1(new_n812), .C2(new_n757), .ZN(new_n813));
  INV_X1    g0613(.A(new_n770), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n499), .B(new_n813), .C1(new_n775), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n774), .A2(G143), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G159), .A2(new_n777), .B1(new_n779), .B2(G137), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n816), .B(new_n817), .C1(new_n818), .C2(new_n753), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n815), .B1(KEYINPUT34), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT34), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n810), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n795), .B(new_n802), .C1(new_n727), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n675), .A2(new_n801), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n654), .B(new_n800), .C1(new_n623), .C2(new_n633), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G330), .ZN(new_n831));
  INV_X1    g0631(.A(new_n711), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n707), .A2(new_n709), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(KEYINPUT94), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n834), .B2(new_n710), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n717), .B1(new_n830), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n830), .A2(new_n836), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n826), .B1(new_n838), .B2(new_n839), .ZN(G384));
  OAI211_X1 g0640(.A(G116), .B(new_n231), .C1(new_n478), .C2(KEYINPUT35), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(KEYINPUT35), .B2(new_n478), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT36), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n234), .B(new_n215), .C1(new_n327), .C2(new_n259), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n202), .A2(G68), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n208), .B(G13), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n707), .A2(new_n711), .A3(new_n709), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n435), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT102), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n370), .A2(new_n371), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n643), .B(KEYINPUT101), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n604), .A2(new_n361), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n361), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n372), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n857), .A2(KEYINPUT37), .B1(new_n860), .B2(new_n855), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n855), .B1(new_n605), .B2(new_n363), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n851), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n855), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n329), .B1(new_n336), .B2(new_n340), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(new_n331), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n358), .B1(new_n866), .B2(new_n360), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n644), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n366), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n361), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n868), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n374), .B2(new_n376), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n874), .A3(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n863), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n390), .A2(new_n654), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n406), .A2(new_n408), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n390), .B(new_n654), .C1(new_n404), .C2(new_n405), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n876), .A2(new_n801), .A3(new_n880), .A4(new_n848), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n848), .A2(new_n801), .A3(new_n880), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n872), .A2(new_n874), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n851), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT40), .B1(new_n885), .B2(new_n875), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n881), .A2(KEYINPUT40), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n850), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n850), .A2(new_n888), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(G330), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n676), .A2(new_n682), .A3(new_n435), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n612), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n891), .B(new_n893), .Z(new_n894));
  OR2_X1    g0694(.A1(new_n406), .A2(new_n654), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n885), .B2(new_n875), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n863), .A2(new_n897), .A3(new_n875), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n885), .A2(new_n875), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n880), .C1(new_n828), .C2(new_n796), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n605), .A2(new_n854), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n894), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n208), .B2(new_n639), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n894), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n847), .B1(new_n908), .B2(new_n909), .ZN(G367));
  OAI21_X1  g0710(.A(new_n731), .B1(new_n212), .B2(new_n415), .ZN(new_n911));
  INV_X1    g0711(.A(new_n736), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n240), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n717), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n774), .A2(G303), .B1(G311), .B2(new_n779), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT107), .Z(new_n916));
  NOR2_X1   g0716(.A1(new_n766), .A2(new_n511), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(KEYINPUT46), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(G107), .B2(new_n814), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n758), .A2(G317), .B1(new_n752), .B2(G294), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n745), .A2(new_n464), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(G283), .B2(new_n777), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n339), .B1(KEYINPUT46), .B2(new_n917), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n919), .A2(new_n920), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n749), .A2(new_n818), .B1(new_n770), .B2(new_n327), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(KEYINPUT108), .ZN(new_n926));
  INV_X1    g0726(.A(G143), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n216), .A2(new_n745), .B1(new_n927), .B2(new_n763), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n775), .B2(new_n767), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n925), .A2(KEYINPUT108), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n289), .B1(new_n758), .B2(G137), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n777), .A2(G50), .B1(new_n752), .B2(G159), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n929), .A2(new_n930), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n916), .A2(new_n924), .B1(new_n926), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT47), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n793), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n914), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n617), .A2(new_n645), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n614), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n620), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n938), .B1(new_n941), .B2(new_n789), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n481), .A2(new_n645), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n487), .A2(new_n489), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT103), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n624), .A2(new_n654), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT103), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n487), .A2(new_n947), .A3(new_n489), .A4(new_n943), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT42), .B1(new_n950), .B2(new_n662), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n600), .B1(new_n945), .B2(new_n948), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n645), .B1(new_n952), .B2(new_n624), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n662), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT42), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n951), .A2(new_n953), .A3(new_n954), .A4(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT104), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n951), .A2(new_n957), .A3(new_n953), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n941), .B(KEYINPUT43), .Z(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT105), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n660), .A2(new_n949), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n960), .A2(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n970));
  INV_X1    g0770(.A(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT105), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n971), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n670), .B(KEYINPUT41), .Z(new_n975));
  NAND2_X1  g0775(.A1(new_n949), .A2(new_n665), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT45), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n664), .A2(new_n946), .A3(new_n945), .A4(new_n948), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n660), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n638), .A2(new_n654), .B1(new_n659), .B2(new_n655), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n662), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n653), .B(new_n983), .C1(new_n719), .C2(KEYINPUT106), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT106), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n653), .A2(KEYINPUT96), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n985), .B1(new_n986), .B2(new_n720), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n984), .B1(new_n987), .B2(new_n983), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n976), .B(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n978), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(new_n992), .A3(new_n661), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n980), .A2(new_n988), .A3(new_n993), .A4(new_n713), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n975), .B1(new_n994), .B2(new_n713), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n974), .B1(new_n995), .B2(new_n716), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n942), .B1(new_n973), .B2(new_n996), .ZN(G387));
  AOI221_X4 g0797(.A(new_n982), .B1(KEYINPUT96), .B2(new_n985), .C1(G330), .C2(new_n652), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT106), .B1(new_n721), .B2(new_n722), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n982), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n676), .A2(new_n682), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n835), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n988), .A2(new_n713), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n1003), .A3(new_n670), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT114), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n760), .A2(new_n807), .B1(new_n763), .B2(new_n750), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n753), .A2(new_n761), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(G317), .C2(new_n774), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT48), .Z(new_n1009));
  OAI22_X1  g0809(.A1(new_n766), .A2(new_n769), .B1(new_n770), .B2(new_n746), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT112), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT113), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT49), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1012), .B(KEYINPUT113), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n745), .A2(new_n511), .B1(new_n757), .B2(new_n764), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n339), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1015), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G68), .A2(new_n777), .B1(new_n779), .B2(G159), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n818), .B2(new_n757), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n216), .A2(new_n766), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1023), .A2(new_n499), .A3(new_n921), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n770), .A2(new_n415), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G50), .B2(new_n804), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT111), .Z(new_n1028));
  OAI211_X1 g0828(.A(new_n1025), .B(new_n1028), .C1(new_n260), .C2(new_n753), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n793), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n668), .A2(new_n733), .B1(G107), .B2(new_n212), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n668), .B(new_n454), .C1(new_n327), .C2(new_n381), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT109), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n412), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n912), .B1(new_n244), .B2(G45), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1031), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n717), .B1(new_n1040), .B2(new_n732), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT110), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1005), .B1(new_n1030), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1021), .A2(new_n1029), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1005), .B(new_n1042), .C1(new_n1044), .C2(new_n727), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n659), .A2(new_n655), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1046), .A2(new_n789), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1043), .A2(new_n1048), .B1(new_n988), .B2(new_n716), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n1004), .A2(new_n1049), .A3(KEYINPUT115), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT115), .B1(new_n1004), .B2(new_n1049), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(G393));
  NAND3_X1  g0853(.A1(new_n980), .A2(new_n716), .A3(new_n993), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n912), .A2(new_n251), .B1(new_n464), .B2(new_n212), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n717), .B1(new_n732), .B2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G317), .A2(new_n779), .B1(new_n804), .B2(G311), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  AOI22_X1  g0858(.A1(new_n814), .A2(G116), .B1(new_n752), .B2(G303), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT116), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n289), .B1(new_n745), .B2(new_n472), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n766), .A2(new_n746), .B1(new_n757), .B2(new_n750), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G294), .C2(new_n777), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1058), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n763), .A2(new_n818), .B1(new_n749), .B2(new_n783), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT51), .Z(new_n1066));
  AOI211_X1 g0866(.A(new_n499), .B(new_n806), .C1(new_n413), .C2(new_n777), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n753), .A2(new_n202), .B1(new_n757), .B2(new_n927), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G68), .B2(new_n767), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n814), .A2(G77), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1064), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1056), .B1(new_n1072), .B2(new_n727), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n730), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1073), .B1(new_n949), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n994), .A2(new_n670), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n980), .A2(new_n993), .B1(new_n988), .B2(new_n713), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1054), .B(new_n1075), .C1(new_n1076), .C2(new_n1077), .ZN(G390));
  INV_X1    g0878(.A(KEYINPUT117), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n880), .B(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n848), .A2(G330), .A3(new_n801), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n712), .A2(G330), .A3(new_n801), .A4(new_n880), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n799), .A2(new_n606), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n796), .B1(new_n681), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1082), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n712), .A2(G330), .A3(new_n801), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n880), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n882), .A2(new_n831), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n796), .B1(new_n675), .B2(new_n801), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT118), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1091), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT118), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1097), .A2(new_n1098), .A3(new_n1094), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1087), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n872), .A2(new_n874), .A3(KEYINPUT38), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT38), .B1(new_n872), .B2(new_n874), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT39), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n863), .A2(new_n897), .A3(new_n875), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n880), .B1(new_n828), .B2(new_n796), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n895), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n876), .A2(new_n895), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n680), .A2(new_n623), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n645), .A3(new_n1085), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n797), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n880), .B(KEYINPUT117), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1091), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1105), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n895), .B1(new_n1094), .B2(new_n1089), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n895), .B(new_n876), .C1(new_n1086), .C2(new_n1080), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1083), .A3(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n849), .A2(G330), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n612), .A2(new_n1121), .A3(new_n892), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1100), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1087), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n880), .B1(new_n835), .B2(new_n801), .ZN(new_n1127));
  OAI211_X1 g0927(.A(KEYINPUT118), .B(new_n1095), .C1(new_n1127), .C2(new_n1091), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1098), .B1(new_n1097), .B2(new_n1094), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1125), .B1(new_n1130), .B2(new_n1122), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1124), .A2(new_n1131), .A3(new_n670), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1115), .A2(new_n728), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n717), .B1(new_n794), .B2(new_n311), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n766), .A2(new_n818), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n758), .A2(G125), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n780), .A2(G50), .B1(new_n804), .B2(G132), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT54), .B(G143), .Z(new_n1140));
  AOI22_X1  g0940(.A1(new_n777), .A2(new_n1140), .B1(new_n752), .B2(G137), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n289), .B1(new_n779), .B2(G128), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n783), .C2(new_n770), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n777), .A2(G97), .B1(new_n752), .B2(G107), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n572), .B2(new_n766), .C1(new_n746), .C2(new_n763), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n758), .A2(G294), .B1(new_n804), .B2(G116), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1146), .A2(new_n289), .A3(new_n811), .A4(new_n1070), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1139), .A2(new_n1143), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1134), .B1(new_n727), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1120), .A2(new_n716), .B1(new_n1133), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1132), .A2(new_n1150), .ZN(G378));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1122), .B1(new_n1100), .B2(new_n1120), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n903), .B1(new_n1105), .B2(new_n896), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n902), .C1(new_n887), .C2(new_n831), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n876), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT40), .B1(new_n1156), .B2(new_n882), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n883), .A2(new_n886), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n831), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n905), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n310), .A2(new_n269), .A3(new_n644), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n310), .B1(new_n269), .B2(new_n644), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  OR3_X1    g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1155), .A2(new_n1160), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1152), .B1(new_n1153), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n905), .A2(new_n1159), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n905), .A2(new_n1159), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1167), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1155), .A2(new_n1160), .A3(new_n1168), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1123), .B1(new_n1130), .B2(new_n1125), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n1178), .A3(KEYINPUT57), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1172), .A2(new_n670), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT121), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n715), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1168), .A2(new_n728), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n717), .B1(new_n794), .B2(G50), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT120), .Z(new_n1186));
  NOR2_X1   g0986(.A1(G33), .A2(G41), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G50), .B(new_n1187), .C1(new_n499), .C2(new_n280), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n758), .A2(G283), .B1(new_n752), .B2(G97), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n472), .B2(new_n749), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1190), .A2(G41), .A3(new_n339), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n259), .A2(new_n745), .B1(new_n760), .B2(new_n415), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1024), .B(new_n1192), .C1(G116), .C2(new_n779), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(new_n327), .C2(new_n770), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1188), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1140), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n766), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT119), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n814), .A2(G150), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n777), .A2(G137), .B1(new_n752), .B2(G132), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G125), .A2(new_n779), .B1(new_n804), .B2(G128), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT59), .ZN(new_n1204));
  INV_X1    g1004(.A(G124), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1187), .B1(new_n757), .B2(new_n1205), .C1(new_n783), .C2(new_n745), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1196), .B1(new_n1195), .B2(new_n1194), .C1(new_n1204), .C2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1186), .B1(new_n1207), .B2(new_n727), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1184), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1182), .B1(new_n1183), .B2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(KEYINPUT121), .B(new_n1209), .C1(new_n1171), .C2(new_n715), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1181), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(G375));
  NAND2_X1  g1016(.A1(new_n1100), .A2(new_n1123), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1122), .B(new_n1087), .C1(new_n1096), .C2(new_n1099), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n975), .B(KEYINPUT122), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G150), .A2(new_n777), .B1(new_n758), .B2(G128), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n812), .B2(new_n763), .C1(new_n783), .C2(new_n766), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G137), .B2(new_n774), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n753), .A2(new_n1197), .B1(new_n745), .B2(new_n259), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n499), .B(new_n1225), .C1(G50), .C2(new_n814), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n745), .A2(new_n381), .B1(new_n763), .B2(new_n769), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n760), .A2(new_n472), .B1(new_n749), .B2(new_n746), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n753), .A2(new_n511), .B1(new_n757), .B2(new_n807), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n289), .B1(new_n766), .B2(new_n464), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1230), .A2(new_n1026), .A3(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1224), .A2(new_n1226), .B1(new_n1229), .B2(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n717), .B1(G68), .B2(new_n794), .C1(new_n1233), .C2(new_n793), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1080), .B2(new_n728), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1100), .B2(new_n716), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1221), .A2(new_n1236), .ZN(G381));
  INV_X1    g1037(.A(KEYINPUT123), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1132), .B2(new_n1150), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1132), .A2(new_n1238), .A3(new_n1150), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1215), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1004), .A2(new_n1049), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT115), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1004), .A2(new_n1049), .A3(KEYINPUT115), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n791), .A3(new_n1246), .ZN(new_n1247));
  OR4_X1    g1047(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1247), .ZN(new_n1248));
  OR3_X1    g1048(.A1(new_n1242), .A2(G381), .A3(new_n1248), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1242), .ZN(G409));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  OAI21_X1  g1051(.A(G396), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1247), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n942), .B(G390), .C1(new_n973), .C2(new_n996), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n994), .A2(new_n713), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n715), .B1(new_n1256), .B2(new_n975), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1257), .A2(new_n974), .A3(new_n972), .A4(new_n969), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G390), .B1(new_n1258), .B2(new_n942), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1251), .B1(new_n1255), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(G390), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1262), .A2(KEYINPUT125), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1258), .A2(KEYINPUT124), .A3(new_n942), .A4(G390), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1254), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1266), .A3(new_n1262), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1253), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1260), .A2(new_n1263), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G343), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(G213), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1218), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n1122), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1217), .A3(new_n1274), .A4(new_n670), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1275), .A2(G384), .A3(new_n1236), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G384), .B1(new_n1275), .B2(new_n1236), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1180), .A2(new_n1213), .A3(G378), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1210), .B1(new_n1177), .B2(new_n716), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1177), .A2(new_n1178), .A3(new_n1220), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1240), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1271), .B(new_n1278), .C1(new_n1279), .C2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1180), .A2(new_n1213), .A3(G378), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1241), .A2(new_n1239), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(new_n1282), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1290), .A2(KEYINPUT62), .A3(new_n1271), .A4(new_n1278), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1287), .A2(KEYINPUT126), .A3(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1271), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1270), .A2(G213), .A3(G2897), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1275), .A2(new_n1236), .ZN(new_n1297));
  INV_X1    g1097(.A(G384), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1275), .A2(G384), .A3(new_n1236), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1300), .A3(new_n1294), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT61), .B1(new_n1293), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1287), .B2(KEYINPUT126), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1269), .B1(new_n1292), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  OR2_X1    g1106(.A1(new_n1285), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1285), .A2(new_n1306), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1307), .A2(new_n1310), .A3(new_n1303), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1305), .A2(new_n1312), .ZN(G405));
  AOI22_X1  g1113(.A1(new_n1283), .A2(new_n1240), .B1(new_n1180), .B2(new_n1213), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1314), .A2(new_n1279), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1269), .B1(new_n1279), .B2(new_n1314), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1320));
  OAI22_X1  g1120(.A1(new_n1319), .A2(new_n1320), .B1(new_n1277), .B2(new_n1276), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT127), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1278), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1321), .A2(new_n1325), .ZN(G402));
endmodule


