

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708;

  NOR2_X1 U362 ( .A1(n626), .A2(n676), .ZN(n627) );
  NOR2_X1 U363 ( .A1(n670), .A2(n676), .ZN(n671) );
  XNOR2_X1 U364 ( .A(n412), .B(n411), .ZN(n533) );
  XNOR2_X1 U365 ( .A(n677), .B(n410), .ZN(n620) );
  XNOR2_X1 U366 ( .A(n404), .B(n451), .ZN(n677) );
  XNOR2_X1 U367 ( .A(n340), .B(n348), .ZN(n410) );
  XNOR2_X1 U368 ( .A(n408), .B(n406), .ZN(n340) );
  XNOR2_X1 U369 ( .A(n396), .B(KEYINPUT65), .ZN(n422) );
  XNOR2_X2 U370 ( .A(n341), .B(n419), .ZN(n514) );
  NOR2_X2 U371 ( .A1(n388), .A2(n418), .ZN(n341) );
  XNOR2_X1 U372 ( .A(n403), .B(n402), .ZN(n451) );
  NOR2_X1 U373 ( .A1(n633), .A2(n676), .ZN(n350) );
  XNOR2_X2 U374 ( .A(n690), .B(G146), .ZN(n369) );
  XNOR2_X2 U375 ( .A(n458), .B(n457), .ZN(n579) );
  NOR2_X2 U376 ( .A1(n513), .A2(n548), .ZN(n458) );
  XNOR2_X2 U377 ( .A(n486), .B(n485), .ZN(n705) );
  INV_X1 U378 ( .A(KEYINPUT4), .ZN(n396) );
  AND2_X1 U379 ( .A1(n703), .A2(n518), .ZN(n394) );
  XNOR2_X1 U380 ( .A(n505), .B(KEYINPUT102), .ZN(n703) );
  OR2_X1 U381 ( .A1(n497), .A2(n360), .ZN(n359) );
  NAND2_X1 U382 ( .A1(n492), .A2(n589), .ZN(n513) );
  XNOR2_X1 U383 ( .A(n365), .B(n445), .ZN(n504) );
  XNOR2_X1 U384 ( .A(n369), .B(n361), .ZN(n660) );
  XNOR2_X1 U385 ( .A(n440), .B(n366), .ZN(n635) );
  XNOR2_X1 U386 ( .A(n370), .B(n481), .ZN(n690) );
  XNOR2_X1 U387 ( .A(n422), .B(G137), .ZN(n370) );
  XNOR2_X1 U388 ( .A(n405), .B(n371), .ZN(n481) );
  XNOR2_X1 U389 ( .A(n351), .B(G122), .ZN(n477) );
  XNOR2_X1 U390 ( .A(G143), .B(G128), .ZN(n405) );
  XNOR2_X1 U391 ( .A(G110), .B(KEYINPUT24), .ZN(n427) );
  XNOR2_X1 U392 ( .A(G128), .B(G119), .ZN(n428) );
  INV_X2 U393 ( .A(G953), .ZN(n696) );
  XOR2_X1 U394 ( .A(G131), .B(G140), .Z(n462) );
  XNOR2_X1 U395 ( .A(G146), .B(G125), .ZN(n431) );
  XOR2_X2 U396 ( .A(G110), .B(G104), .Z(n423) );
  NOR2_X1 U397 ( .A1(n705), .A2(n646), .ZN(n342) );
  BUF_X1 U398 ( .A(n664), .Z(n672) );
  NOR2_X2 U399 ( .A1(n484), .A2(n552), .ZN(n486) );
  XNOR2_X2 U400 ( .A(n544), .B(KEYINPUT1), .ZN(n492) );
  XNOR2_X2 U401 ( .A(n426), .B(n425), .ZN(n544) );
  OR2_X1 U402 ( .A1(n389), .A2(KEYINPUT84), .ZN(n360) );
  NOR2_X1 U403 ( .A1(G237), .A2(G953), .ZN(n453) );
  XNOR2_X1 U404 ( .A(n452), .B(n387), .ZN(n386) );
  INV_X1 U405 ( .A(G116), .ZN(n387) );
  XOR2_X1 U406 ( .A(KEYINPUT5), .B(G131), .Z(n452) );
  XNOR2_X1 U407 ( .A(G113), .B(G122), .ZN(n468) );
  XNOR2_X1 U408 ( .A(G143), .B(G104), .ZN(n463) );
  XOR2_X1 U409 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n464) );
  XNOR2_X1 U410 ( .A(n461), .B(n367), .ZN(n689) );
  INV_X1 U411 ( .A(n462), .ZN(n367) );
  XNOR2_X1 U412 ( .A(n401), .B(KEYINPUT69), .ZN(n402) );
  XNOR2_X1 U413 ( .A(G101), .B(KEYINPUT3), .ZN(n400) );
  OR2_X1 U414 ( .A1(n635), .A2(G902), .ZN(n365) );
  XNOR2_X1 U415 ( .A(n431), .B(KEYINPUT10), .ZN(n461) );
  XNOR2_X1 U416 ( .A(n364), .B(n362), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n424), .B(n363), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n352), .B(n477), .ZN(n404) );
  XNOR2_X1 U419 ( .A(n423), .B(n353), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n354), .B(KEYINPUT72), .ZN(n353) );
  NAND2_X1 U421 ( .A1(G234), .A2(G237), .ZN(n416) );
  AND2_X1 U422 ( .A1(n381), .A2(n380), .ZN(n569) );
  XNOR2_X1 U423 ( .A(n382), .B(KEYINPUT105), .ZN(n381) );
  NAND2_X1 U424 ( .A1(n383), .A2(n502), .ZN(n382) );
  XOR2_X1 U425 ( .A(G472), .B(n345), .Z(n594) );
  AND2_X1 U426 ( .A1(n358), .A2(n504), .ZN(n357) );
  NAND2_X1 U427 ( .A1(n389), .A2(KEYINPUT84), .ZN(n358) );
  XNOR2_X1 U428 ( .A(n491), .B(n490), .ZN(n497) );
  XNOR2_X1 U429 ( .A(n625), .B(n624), .ZN(n676) );
  XNOR2_X1 U430 ( .A(G119), .B(KEYINPUT68), .ZN(n401) );
  XNOR2_X1 U431 ( .A(G101), .B(G107), .ZN(n363) );
  INV_X1 U432 ( .A(KEYINPUT16), .ZN(n354) );
  INV_X1 U433 ( .A(n581), .ZN(n398) );
  NAND2_X1 U434 ( .A1(n493), .A2(n548), .ZN(n389) );
  XNOR2_X1 U435 ( .A(n451), .B(n385), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n454), .B(n386), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n391), .B(KEYINPUT70), .ZN(n390) );
  INV_X1 U438 ( .A(G134), .ZN(n371) );
  XNOR2_X1 U439 ( .A(G116), .B(G107), .ZN(n351) );
  XNOR2_X1 U440 ( .A(KEYINPUT7), .B(KEYINPUT100), .ZN(n474) );
  XOR2_X1 U441 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n475) );
  XNOR2_X1 U442 ( .A(n368), .B(n689), .ZN(n665) );
  XNOR2_X1 U443 ( .A(n471), .B(n467), .ZN(n368) );
  XNOR2_X1 U444 ( .A(n344), .B(n466), .ZN(n467) );
  OR2_X1 U445 ( .A1(n550), .A2(n551), .ZN(n379) );
  INV_X1 U446 ( .A(KEYINPUT36), .ZN(n378) );
  INV_X1 U447 ( .A(KEYINPUT0), .ZN(n419) );
  XNOR2_X1 U448 ( .A(n551), .B(n414), .ZN(n388) );
  INV_X1 U449 ( .A(KEYINPUT19), .ZN(n414) );
  XNOR2_X1 U450 ( .A(n510), .B(KEYINPUT94), .ZN(n521) );
  XNOR2_X1 U451 ( .A(n439), .B(n438), .ZN(n366) );
  XNOR2_X1 U452 ( .A(n375), .B(n374), .ZN(n700) );
  INV_X1 U453 ( .A(KEYINPUT110), .ZN(n374) );
  NAND2_X1 U454 ( .A1(n377), .A2(n376), .ZN(n375) );
  XNOR2_X1 U455 ( .A(n379), .B(n378), .ZN(n377) );
  OR2_X1 U456 ( .A1(n497), .A2(n376), .ZN(n503) );
  NAND2_X1 U457 ( .A1(n356), .A2(n355), .ZN(n505) );
  AND2_X1 U458 ( .A1(n359), .A2(n357), .ZN(n356) );
  XNOR2_X1 U459 ( .A(n349), .B(n347), .ZN(n663) );
  NAND2_X1 U460 ( .A1(n672), .A2(G469), .ZN(n349) );
  AND2_X1 U461 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U462 ( .A(n345), .B(n455), .ZN(n502) );
  INV_X1 U463 ( .A(n502), .ZN(n548) );
  NOR2_X1 U464 ( .A1(n528), .A2(n531), .ZN(n343) );
  XOR2_X1 U465 ( .A(n464), .B(n463), .Z(n344) );
  NOR2_X1 U466 ( .A1(n628), .A2(G902), .ZN(n345) );
  AND2_X1 U467 ( .A1(n706), .A2(n373), .ZN(n346) );
  INV_X1 U468 ( .A(n492), .ZN(n493) );
  INV_X1 U469 ( .A(n493), .ZN(n376) );
  INV_X1 U470 ( .A(n531), .ZN(n532) );
  INV_X1 U471 ( .A(n638), .ZN(n380) );
  XOR2_X1 U472 ( .A(n662), .B(n661), .Z(n347) );
  NAND2_X1 U473 ( .A1(n533), .A2(n584), .ZN(n551) );
  XNOR2_X1 U474 ( .A(n421), .B(n422), .ZN(n348) );
  XNOR2_X1 U475 ( .A(n350), .B(n634), .ZN(G57) );
  NAND2_X1 U476 ( .A1(n497), .A2(KEYINPUT84), .ZN(n355) );
  XNOR2_X1 U477 ( .A(n423), .B(n462), .ZN(n364) );
  XNOR2_X1 U478 ( .A(n369), .B(n384), .ZN(n628) );
  INV_X1 U479 ( .A(n405), .ZN(n421) );
  NAND2_X1 U480 ( .A1(n501), .A2(n706), .ZN(n372) );
  NAND2_X1 U481 ( .A1(n342), .A2(n346), .ZN(n391) );
  NAND2_X1 U482 ( .A1(n372), .A2(KEYINPUT44), .ZN(n395) );
  INV_X1 U483 ( .A(KEYINPUT44), .ZN(n373) );
  XNOR2_X1 U484 ( .A(n399), .B(n535), .ZN(n567) );
  INV_X1 U485 ( .A(n549), .ZN(n383) );
  NOR2_X1 U486 ( .A1(n555), .A2(n388), .ZN(n650) );
  NAND2_X1 U487 ( .A1(n392), .A2(n390), .ZN(n520) );
  XNOR2_X1 U488 ( .A(n393), .B(KEYINPUT85), .ZN(n392) );
  NAND2_X1 U489 ( .A1(n395), .A2(n394), .ZN(n393) );
  NOR2_X1 U490 ( .A1(n528), .A2(n397), .ZN(n399) );
  NAND2_X1 U491 ( .A1(n532), .A2(n398), .ZN(n397) );
  NOR2_X2 U492 ( .A1(n618), .A2(n617), .ZN(n664) );
  XNOR2_X1 U493 ( .A(G472), .B(KEYINPUT6), .ZN(n455) );
  XNOR2_X1 U494 ( .A(n456), .B(KEYINPUT33), .ZN(n457) );
  INV_X1 U495 ( .A(KEYINPUT34), .ZN(n459) );
  BUF_X1 U496 ( .A(n533), .Z(n572) );
  XNOR2_X1 U497 ( .A(KEYINPUT77), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U498 ( .A(n400), .B(G113), .ZN(n403) );
  XOR2_X1 U499 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n406) );
  NAND2_X1 U500 ( .A1(G224), .A2(n696), .ZN(n407) );
  XNOR2_X1 U501 ( .A(n431), .B(n407), .ZN(n408) );
  XNOR2_X1 U502 ( .A(KEYINPUT15), .B(G902), .ZN(n617) );
  NAND2_X1 U503 ( .A1(n620), .A2(n617), .ZN(n412) );
  OR2_X1 U504 ( .A1(G237), .A2(G902), .ZN(n413) );
  AND2_X1 U505 ( .A1(G210), .A2(n413), .ZN(n411) );
  NAND2_X1 U506 ( .A1(G214), .A2(n413), .ZN(n584) );
  XOR2_X1 U507 ( .A(G898), .B(KEYINPUT89), .Z(n682) );
  NOR2_X1 U508 ( .A1(n682), .A2(n696), .ZN(n679) );
  NAND2_X1 U509 ( .A1(n679), .A2(G902), .ZN(n415) );
  NAND2_X1 U510 ( .A1(G952), .A2(n696), .ZN(n523) );
  NAND2_X1 U511 ( .A1(n415), .A2(n523), .ZN(n417) );
  XNOR2_X1 U512 ( .A(n416), .B(KEYINPUT14), .ZN(n578) );
  NAND2_X1 U513 ( .A1(n417), .A2(n578), .ZN(n418) );
  XNOR2_X1 U514 ( .A(n514), .B(KEYINPUT90), .ZN(n509) );
  NAND2_X1 U515 ( .A1(G227), .A2(n696), .ZN(n424) );
  NOR2_X1 U516 ( .A1(n660), .A2(G902), .ZN(n426) );
  XNOR2_X1 U517 ( .A(KEYINPUT67), .B(G469), .ZN(n425) );
  XNOR2_X1 U518 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U519 ( .A(KEYINPUT23), .B(KEYINPUT76), .ZN(n429) );
  XNOR2_X1 U520 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U521 ( .A(n432), .B(n461), .ZN(n440) );
  NAND2_X1 U522 ( .A1(G234), .A2(n696), .ZN(n434) );
  INV_X1 U523 ( .A(KEYINPUT8), .ZN(n433) );
  XNOR2_X1 U524 ( .A(n434), .B(n433), .ZN(n478) );
  NAND2_X1 U525 ( .A1(n478), .A2(G221), .ZN(n439) );
  INV_X1 U526 ( .A(G140), .ZN(n435) );
  XNOR2_X1 U527 ( .A(n435), .B(G137), .ZN(n437) );
  XNOR2_X1 U528 ( .A(KEYINPUT80), .B(KEYINPUT91), .ZN(n436) );
  XNOR2_X1 U529 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U530 ( .A1(G234), .A2(n617), .ZN(n441) );
  XNOR2_X1 U531 ( .A(KEYINPUT20), .B(n441), .ZN(n446) );
  NAND2_X1 U532 ( .A1(n446), .A2(G217), .ZN(n444) );
  INV_X1 U533 ( .A(KEYINPUT92), .ZN(n442) );
  XNOR2_X1 U534 ( .A(n442), .B(KEYINPUT25), .ZN(n443) );
  XNOR2_X1 U535 ( .A(n444), .B(n443), .ZN(n445) );
  NAND2_X1 U536 ( .A1(n446), .A2(G221), .ZN(n449) );
  INV_X1 U537 ( .A(KEYINPUT93), .ZN(n447) );
  XNOR2_X1 U538 ( .A(n447), .B(KEYINPUT21), .ZN(n448) );
  XNOR2_X1 U539 ( .A(n449), .B(n448), .ZN(n591) );
  INV_X1 U540 ( .A(n591), .ZN(n450) );
  AND2_X1 U541 ( .A1(n504), .A2(n450), .ZN(n589) );
  XNOR2_X1 U542 ( .A(n453), .B(KEYINPUT74), .ZN(n465) );
  NAND2_X1 U543 ( .A1(G210), .A2(n465), .ZN(n454) );
  XNOR2_X1 U544 ( .A(KEYINPUT86), .B(KEYINPUT104), .ZN(n456) );
  NOR2_X1 U545 ( .A1(n509), .A2(n579), .ZN(n460) );
  XNOR2_X1 U546 ( .A(n460), .B(n459), .ZN(n484) );
  NAND2_X1 U547 ( .A1(G214), .A2(n465), .ZN(n466) );
  XOR2_X1 U548 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n469) );
  XNOR2_X1 U549 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U550 ( .A(KEYINPUT11), .B(n470), .Z(n471) );
  NOR2_X1 U551 ( .A1(G902), .A2(n665), .ZN(n473) );
  XOR2_X1 U552 ( .A(KEYINPUT13), .B(G475), .Z(n472) );
  XNOR2_X1 U553 ( .A(n473), .B(n472), .ZN(n508) );
  XNOR2_X1 U554 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U555 ( .A(n477), .B(n476), .Z(n480) );
  NAND2_X1 U556 ( .A1(G217), .A2(n478), .ZN(n479) );
  XNOR2_X1 U557 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U558 ( .A(n482), .B(n481), .ZN(n673) );
  NOR2_X1 U559 ( .A1(G902), .A2(n673), .ZN(n483) );
  XNOR2_X1 U560 ( .A(G478), .B(n483), .ZN(n506) );
  OR2_X1 U561 ( .A1(n508), .A2(n506), .ZN(n552) );
  NAND2_X1 U562 ( .A1(n508), .A2(n506), .ZN(n582) );
  NOR2_X1 U563 ( .A1(n591), .A2(n582), .ZN(n487) );
  XNOR2_X1 U564 ( .A(n487), .B(KEYINPUT101), .ZN(n488) );
  NOR2_X1 U565 ( .A1(n514), .A2(n488), .ZN(n491) );
  XNOR2_X1 U566 ( .A(KEYINPUT64), .B(KEYINPUT71), .ZN(n489) );
  XNOR2_X1 U567 ( .A(n489), .B(KEYINPUT22), .ZN(n490) );
  INV_X1 U568 ( .A(n504), .ZN(n592) );
  INV_X1 U569 ( .A(n594), .ZN(n542) );
  NAND2_X1 U570 ( .A1(n592), .A2(n542), .ZN(n494) );
  NOR2_X1 U571 ( .A1(n503), .A2(n494), .ZN(n646) );
  NOR2_X1 U572 ( .A1(n705), .A2(n646), .ZN(n501) );
  XNOR2_X1 U573 ( .A(n548), .B(KEYINPUT78), .ZN(n499) );
  NAND2_X1 U574 ( .A1(n492), .A2(n592), .ZN(n495) );
  XOR2_X1 U575 ( .A(KEYINPUT103), .B(n495), .Z(n496) );
  NOR2_X1 U576 ( .A1(n497), .A2(n496), .ZN(n498) );
  NAND2_X1 U577 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U578 ( .A(n500), .B(KEYINPUT32), .ZN(n706) );
  INV_X1 U579 ( .A(n506), .ZN(n507) );
  AND2_X1 U580 ( .A1(n508), .A2(n507), .ZN(n656) );
  INV_X1 U581 ( .A(n656), .ZN(n568) );
  OR2_X1 U582 ( .A1(n508), .A2(n507), .ZN(n638) );
  AND2_X1 U583 ( .A1(n568), .A2(n638), .ZN(n580) );
  INV_X1 U584 ( .A(n509), .ZN(n512) );
  NAND2_X1 U585 ( .A1(n544), .A2(n589), .ZN(n510) );
  NOR2_X1 U586 ( .A1(n521), .A2(n594), .ZN(n511) );
  AND2_X1 U587 ( .A1(n512), .A2(n511), .ZN(n641) );
  OR2_X1 U588 ( .A1(n513), .A2(n542), .ZN(n599) );
  NOR2_X1 U589 ( .A1(n514), .A2(n599), .ZN(n516) );
  XNOR2_X1 U590 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n515) );
  XNOR2_X1 U591 ( .A(n516), .B(n515), .ZN(n657) );
  NOR2_X1 U592 ( .A1(n641), .A2(n657), .ZN(n517) );
  OR2_X1 U593 ( .A1(n580), .A2(n517), .ZN(n518) );
  INV_X1 U594 ( .A(KEYINPUT45), .ZN(n519) );
  XNOR2_X1 U595 ( .A(n520), .B(n519), .ZN(n684) );
  XNOR2_X1 U596 ( .A(n521), .B(KEYINPUT106), .ZN(n526) );
  NOR2_X1 U597 ( .A1(G900), .A2(n696), .ZN(n522) );
  NAND2_X1 U598 ( .A1(G902), .A2(n522), .ZN(n524) );
  NAND2_X1 U599 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U600 ( .A1(n525), .A2(n578), .ZN(n539) );
  NOR2_X1 U601 ( .A1(n526), .A2(n539), .ZN(n527) );
  XNOR2_X1 U602 ( .A(n527), .B(KEYINPUT75), .ZN(n528) );
  NAND2_X1 U603 ( .A1(n584), .A2(n594), .ZN(n530) );
  XOR2_X1 U604 ( .A(KEYINPUT107), .B(KEYINPUT30), .Z(n529) );
  XNOR2_X1 U605 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U606 ( .A(KEYINPUT73), .B(KEYINPUT38), .Z(n534) );
  XNOR2_X1 U607 ( .A(n572), .B(n534), .ZN(n581) );
  XOR2_X1 U608 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n535) );
  NOR2_X1 U609 ( .A1(n567), .A2(n638), .ZN(n536) );
  XNOR2_X1 U610 ( .A(n536), .B(KEYINPUT40), .ZN(n616) );
  NOR2_X1 U611 ( .A1(n581), .A2(n582), .ZN(n587) );
  NAND2_X1 U612 ( .A1(n587), .A2(n584), .ZN(n538) );
  XOR2_X1 U613 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n537) );
  XNOR2_X1 U614 ( .A(n538), .B(n537), .ZN(n609) );
  NOR2_X1 U615 ( .A1(n591), .A2(n539), .ZN(n540) );
  NAND2_X1 U616 ( .A1(n592), .A2(n540), .ZN(n541) );
  XNOR2_X1 U617 ( .A(n541), .B(KEYINPUT66), .ZN(n549) );
  NOR2_X1 U618 ( .A1(n549), .A2(n542), .ZN(n543) );
  XNOR2_X1 U619 ( .A(KEYINPUT28), .B(n543), .ZN(n545) );
  NAND2_X1 U620 ( .A1(n545), .A2(n544), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n609), .A2(n555), .ZN(n546) );
  XNOR2_X1 U622 ( .A(n546), .B(KEYINPUT42), .ZN(n708) );
  NOR2_X1 U623 ( .A1(n616), .A2(n708), .ZN(n547) );
  XNOR2_X1 U624 ( .A(n547), .B(KEYINPUT46), .ZN(n564) );
  XNOR2_X1 U625 ( .A(n569), .B(KEYINPUT109), .ZN(n550) );
  INV_X1 U626 ( .A(n572), .ZN(n553) );
  NOR2_X1 U627 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U628 ( .A1(n343), .A2(n554), .ZN(n649) );
  INV_X1 U629 ( .A(n580), .ZN(n556) );
  NAND2_X1 U630 ( .A1(n650), .A2(n556), .ZN(n559) );
  NAND2_X1 U631 ( .A1(KEYINPUT47), .A2(n559), .ZN(n557) );
  NAND2_X1 U632 ( .A1(n649), .A2(n557), .ZN(n558) );
  XNOR2_X1 U633 ( .A(n558), .B(KEYINPUT79), .ZN(n561) );
  OR2_X1 U634 ( .A1(n559), .A2(KEYINPUT47), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U636 ( .A1(n700), .A2(n562), .ZN(n563) );
  NAND2_X1 U637 ( .A1(n564), .A2(n563), .ZN(n566) );
  XOR2_X1 U638 ( .A(KEYINPUT82), .B(KEYINPUT48), .Z(n565) );
  XNOR2_X1 U639 ( .A(n566), .B(n565), .ZN(n575) );
  NOR2_X1 U640 ( .A1(n567), .A2(n568), .ZN(n615) );
  NAND2_X1 U641 ( .A1(n569), .A2(n584), .ZN(n570) );
  NOR2_X1 U642 ( .A1(n492), .A2(n570), .ZN(n571) );
  XNOR2_X1 U643 ( .A(n571), .B(KEYINPUT43), .ZN(n573) );
  NOR2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n659) );
  NOR2_X1 U645 ( .A1(n615), .A2(n659), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n694) );
  NOR2_X1 U647 ( .A1(n684), .A2(n694), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT2), .ZN(n618) );
  XNOR2_X1 U649 ( .A(n618), .B(KEYINPUT81), .ZN(n577) );
  NOR2_X1 U650 ( .A1(n577), .A2(G953), .ZN(n613) );
  NAND2_X1 U651 ( .A1(G952), .A2(n578), .ZN(n607) );
  OR2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n585) );
  AND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U656 ( .A1(n579), .A2(n588), .ZN(n603) );
  NOR2_X1 U657 ( .A1(n492), .A2(n589), .ZN(n590) );
  XOR2_X1 U658 ( .A(KEYINPUT50), .B(n590), .Z(n597) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n593), .B(KEYINPUT49), .ZN(n595) );
  NOR2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U664 ( .A(KEYINPUT51), .B(n600), .ZN(n601) );
  NOR2_X1 U665 ( .A1(n609), .A2(n601), .ZN(n602) );
  NOR2_X1 U666 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U667 ( .A(KEYINPUT119), .B(n604), .Z(n605) );
  XNOR2_X1 U668 ( .A(KEYINPUT52), .B(n605), .ZN(n606) );
  NOR2_X1 U669 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U670 ( .A(n608), .B(KEYINPUT120), .ZN(n611) );
  NOR2_X1 U671 ( .A1(n579), .A2(n609), .ZN(n610) );
  NOR2_X1 U672 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U673 ( .A(n614), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U674 ( .A(G134), .B(n615), .Z(G36) );
  XOR2_X1 U675 ( .A(n616), .B(G131), .Z(G33) );
  NAND2_X1 U676 ( .A1(n664), .A2(G210), .ZN(n622) );
  XNOR2_X1 U677 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n619) );
  XNOR2_X1 U678 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U679 ( .A(n622), .B(n621), .ZN(n626) );
  INV_X1 U680 ( .A(G952), .ZN(n623) );
  NAND2_X1 U681 ( .A1(n623), .A2(G953), .ZN(n625) );
  INV_X1 U682 ( .A(KEYINPUT88), .ZN(n624) );
  XNOR2_X1 U683 ( .A(n627), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U684 ( .A1(n664), .A2(G472), .ZN(n632) );
  XOR2_X1 U685 ( .A(KEYINPUT87), .B(KEYINPUT62), .Z(n630) );
  XOR2_X1 U686 ( .A(n628), .B(KEYINPUT111), .Z(n629) );
  XNOR2_X1 U687 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U688 ( .A(n632), .B(n631), .ZN(n633) );
  INV_X1 U689 ( .A(KEYINPUT63), .ZN(n634) );
  NAND2_X1 U690 ( .A1(n672), .A2(G217), .ZN(n636) );
  XNOR2_X1 U691 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X1 U692 ( .A1(n637), .A2(n676), .ZN(G66) );
  XOR2_X1 U693 ( .A(G104), .B(KEYINPUT113), .Z(n640) );
  NAND2_X1 U694 ( .A1(n641), .A2(n380), .ZN(n639) );
  XNOR2_X1 U695 ( .A(n640), .B(n639), .ZN(G6) );
  XNOR2_X1 U696 ( .A(G107), .B(KEYINPUT27), .ZN(n645) );
  XOR2_X1 U697 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n643) );
  NAND2_X1 U698 ( .A1(n641), .A2(n656), .ZN(n642) );
  XNOR2_X1 U699 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U700 ( .A(n645), .B(n644), .ZN(G9) );
  XOR2_X1 U701 ( .A(G110), .B(n646), .Z(G12) );
  XOR2_X1 U702 ( .A(G128), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U703 ( .A1(n650), .A2(n656), .ZN(n647) );
  XNOR2_X1 U704 ( .A(n648), .B(n647), .ZN(G30) );
  XNOR2_X1 U705 ( .A(G143), .B(n649), .ZN(G45) );
  XOR2_X1 U706 ( .A(G146), .B(KEYINPUT115), .Z(n652) );
  NAND2_X1 U707 ( .A1(n650), .A2(n380), .ZN(n651) );
  XNOR2_X1 U708 ( .A(n652), .B(n651), .ZN(G48) );
  XOR2_X1 U709 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n654) );
  NAND2_X1 U710 ( .A1(n657), .A2(n380), .ZN(n653) );
  XNOR2_X1 U711 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U712 ( .A(G113), .B(n655), .ZN(G15) );
  NAND2_X1 U713 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U714 ( .A(n658), .B(G116), .ZN(G18) );
  XOR2_X1 U715 ( .A(G140), .B(n659), .Z(G42) );
  XOR2_X1 U716 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n662) );
  XNOR2_X1 U717 ( .A(n660), .B(KEYINPUT121), .ZN(n661) );
  NOR2_X1 U718 ( .A1(n676), .A2(n663), .ZN(G54) );
  NAND2_X1 U719 ( .A1(n664), .A2(G475), .ZN(n669) );
  XNOR2_X1 U720 ( .A(KEYINPUT59), .B(KEYINPUT122), .ZN(n667) );
  XNOR2_X1 U721 ( .A(n665), .B(KEYINPUT123), .ZN(n666) );
  XNOR2_X1 U722 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U723 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U724 ( .A(n671), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U725 ( .A1(n672), .A2(G478), .ZN(n674) );
  XNOR2_X1 U726 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U727 ( .A1(n676), .A2(n675), .ZN(G63) );
  XNOR2_X1 U728 ( .A(n677), .B(KEYINPUT124), .ZN(n678) );
  XNOR2_X1 U729 ( .A(n678), .B(KEYINPUT125), .ZN(n680) );
  NOR2_X1 U730 ( .A1(n680), .A2(n679), .ZN(n688) );
  NAND2_X1 U731 ( .A1(G953), .A2(G224), .ZN(n681) );
  XNOR2_X1 U732 ( .A(n681), .B(KEYINPUT61), .ZN(n683) );
  NAND2_X1 U733 ( .A1(n683), .A2(n682), .ZN(n686) );
  OR2_X1 U734 ( .A1(G953), .A2(n684), .ZN(n685) );
  NAND2_X1 U735 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U736 ( .A(n688), .B(n687), .ZN(G69) );
  XNOR2_X1 U737 ( .A(n690), .B(n689), .ZN(n695) );
  XNOR2_X1 U738 ( .A(G227), .B(n695), .ZN(n691) );
  NAND2_X1 U739 ( .A1(n691), .A2(G900), .ZN(n692) );
  NAND2_X1 U740 ( .A1(n692), .A2(G953), .ZN(n693) );
  XNOR2_X1 U741 ( .A(n693), .B(KEYINPUT126), .ZN(n699) );
  XNOR2_X1 U742 ( .A(n694), .B(n695), .ZN(n697) );
  NAND2_X1 U743 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U744 ( .A1(n699), .A2(n698), .ZN(G72) );
  XNOR2_X1 U745 ( .A(KEYINPUT118), .B(KEYINPUT37), .ZN(n701) );
  XNOR2_X1 U746 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U747 ( .A(G125), .B(n702), .ZN(G27) );
  XNOR2_X1 U748 ( .A(n703), .B(G101), .ZN(n704) );
  XNOR2_X1 U749 ( .A(n704), .B(KEYINPUT112), .ZN(G3) );
  XOR2_X1 U750 ( .A(n705), .B(G122), .Z(G24) );
  XOR2_X1 U751 ( .A(G119), .B(n706), .Z(n707) );
  XNOR2_X1 U752 ( .A(KEYINPUT127), .B(n707), .ZN(G21) );
  XOR2_X1 U753 ( .A(G137), .B(n708), .Z(G39) );
endmodule

