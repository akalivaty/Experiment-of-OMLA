

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U548 ( .A1(n695), .A2(n694), .ZN(n735) );
  NOR2_X1 U549 ( .A1(n979), .A2(n697), .ZN(n699) );
  NOR2_X1 U550 ( .A1(n710), .A2(n971), .ZN(n700) );
  NOR2_X1 U551 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  NOR2_X1 U552 ( .A1(G651), .A2(n628), .ZN(n634) );
  AND2_X1 U553 ( .A1(n523), .A2(n522), .ZN(n681) );
  XOR2_X1 U554 ( .A(KEYINPUT23), .B(KEYINPUT65), .Z(n514) );
  INV_X1 U555 ( .A(G2105), .ZN(n520) );
  AND2_X1 U556 ( .A1(n520), .A2(G2104), .ZN(n878) );
  NAND2_X1 U557 ( .A1(G101), .A2(n878), .ZN(n513) );
  XOR2_X1 U558 ( .A(n514), .B(n513), .Z(n680) );
  XOR2_X2 U559 ( .A(KEYINPUT17), .B(n515), .Z(n877) );
  NAND2_X1 U560 ( .A1(n877), .A2(G137), .ZN(n516) );
  XNOR2_X1 U561 ( .A(n516), .B(KEYINPUT66), .ZN(n518) );
  AND2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U563 ( .A1(G113), .A2(n882), .ZN(n517) );
  NAND2_X1 U564 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U565 ( .A(KEYINPUT67), .B(n519), .ZN(n523) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n520), .ZN(n881) );
  NAND2_X1 U567 ( .A1(G125), .A2(n881), .ZN(n521) );
  XNOR2_X1 U568 ( .A(n521), .B(KEYINPUT64), .ZN(n522) );
  AND2_X1 U569 ( .A1(n680), .A2(n681), .ZN(G160) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n631) );
  NAND2_X1 U571 ( .A1(G85), .A2(n631), .ZN(n525) );
  XOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  INV_X1 U573 ( .A(G651), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n628), .A2(n526), .ZN(n637) );
  NAND2_X1 U575 ( .A1(G72), .A2(n637), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U577 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n527), .Z(n633) );
  NAND2_X1 U579 ( .A1(G60), .A2(n633), .ZN(n529) );
  NAND2_X1 U580 ( .A1(G47), .A2(n634), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U582 ( .A1(n531), .A2(n530), .ZN(G290) );
  NAND2_X1 U583 ( .A1(G64), .A2(n633), .ZN(n533) );
  NAND2_X1 U584 ( .A1(G52), .A2(n634), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n539) );
  NAND2_X1 U586 ( .A1(n637), .A2(G77), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT68), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G90), .A2(n631), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U590 ( .A(KEYINPUT9), .B(n537), .Z(n538) );
  NOR2_X1 U591 ( .A1(n539), .A2(n538), .ZN(G171) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G57), .ZN(G237) );
  INV_X1 U594 ( .A(G132), .ZN(G219) );
  INV_X1 U595 ( .A(G82), .ZN(G220) );
  NAND2_X1 U596 ( .A1(n637), .A2(G76), .ZN(n540) );
  XNOR2_X1 U597 ( .A(KEYINPUT74), .B(n540), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n631), .A2(G89), .ZN(n541) );
  XNOR2_X1 U599 ( .A(KEYINPUT4), .B(n541), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n544), .B(KEYINPUT5), .ZN(n549) );
  NAND2_X1 U602 ( .A1(G63), .A2(n633), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G51), .A2(n634), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U607 ( .A(n550), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(G7), .A2(G661), .ZN(n551) );
  XNOR2_X1 U610 ( .A(n551), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U611 ( .A(G223), .ZN(n822) );
  NAND2_X1 U612 ( .A1(n822), .A2(G567), .ZN(n552) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(n552), .Z(G234) );
  NAND2_X1 U614 ( .A1(G56), .A2(n633), .ZN(n553) );
  XOR2_X1 U615 ( .A(KEYINPUT14), .B(n553), .Z(n559) );
  NAND2_X1 U616 ( .A1(n631), .A2(G81), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(KEYINPUT12), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G68), .A2(n637), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT13), .B(n557), .Z(n558) );
  NOR2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n634), .A2(G43), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n561), .A2(n560), .ZN(n979) );
  INV_X1 U624 ( .A(G860), .ZN(n585) );
  OR2_X1 U625 ( .A1(n979), .A2(n585), .ZN(G153) );
  INV_X1 U626 ( .A(G171), .ZN(G301) );
  NAND2_X1 U627 ( .A1(G868), .A2(G301), .ZN(n573) );
  NAND2_X1 U628 ( .A1(G66), .A2(n633), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G92), .A2(n631), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT71), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G79), .A2(n637), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n634), .A2(G54), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT72), .B(n567), .Z(n568) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(n570), .B(KEYINPUT15), .Z(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT73), .B(n571), .ZN(n971) );
  INV_X1 U639 ( .A(G868), .ZN(n654) );
  NAND2_X1 U640 ( .A1(n971), .A2(n654), .ZN(n572) );
  NAND2_X1 U641 ( .A1(n573), .A2(n572), .ZN(G284) );
  NAND2_X1 U642 ( .A1(G53), .A2(n634), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT70), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G91), .A2(n631), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G78), .A2(n637), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U647 ( .A1(G65), .A2(n633), .ZN(n577) );
  XNOR2_X1 U648 ( .A(KEYINPUT69), .B(n577), .ZN(n578) );
  NOR2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(G299) );
  NOR2_X1 U651 ( .A1(G286), .A2(n654), .ZN(n583) );
  NOR2_X1 U652 ( .A1(G868), .A2(G299), .ZN(n582) );
  NOR2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U654 ( .A(KEYINPUT75), .B(n584), .Z(G297) );
  NAND2_X1 U655 ( .A1(n585), .A2(G559), .ZN(n586) );
  INV_X1 U656 ( .A(n971), .ZN(n609) );
  NAND2_X1 U657 ( .A1(n586), .A2(n609), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U659 ( .A1(n609), .A2(G868), .ZN(n588) );
  NOR2_X1 U660 ( .A1(G559), .A2(n588), .ZN(n589) );
  XNOR2_X1 U661 ( .A(n589), .B(KEYINPUT76), .ZN(n591) );
  NOR2_X1 U662 ( .A1(n979), .A2(G868), .ZN(n590) );
  NOR2_X1 U663 ( .A1(n591), .A2(n590), .ZN(G282) );
  XOR2_X1 U664 ( .A(G2100), .B(KEYINPUT78), .Z(n601) );
  NAND2_X1 U665 ( .A1(G123), .A2(n881), .ZN(n592) );
  XOR2_X1 U666 ( .A(KEYINPUT18), .B(n592), .Z(n593) );
  XNOR2_X1 U667 ( .A(n593), .B(KEYINPUT77), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G111), .A2(n882), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U670 ( .A1(G135), .A2(n877), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G99), .A2(n878), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n914) );
  XNOR2_X1 U674 ( .A(G2096), .B(n914), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(G156) );
  NAND2_X1 U676 ( .A1(G67), .A2(n633), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G55), .A2(n634), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U679 ( .A(KEYINPUT80), .B(n604), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G93), .A2(n631), .ZN(n606) );
  NAND2_X1 U681 ( .A1(G80), .A2(n637), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n655) );
  NAND2_X1 U684 ( .A1(G559), .A2(n609), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n610), .B(n979), .ZN(n652) );
  NOR2_X1 U686 ( .A1(G860), .A2(n652), .ZN(n612) );
  XNOR2_X1 U687 ( .A(KEYINPUT79), .B(KEYINPUT81), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n655), .B(n613), .ZN(G145) );
  NAND2_X1 U690 ( .A1(n631), .A2(G86), .ZN(n614) );
  XOR2_X1 U691 ( .A(KEYINPUT83), .B(n614), .Z(n616) );
  NAND2_X1 U692 ( .A1(n633), .A2(G61), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U694 ( .A(KEYINPUT84), .B(n617), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G73), .A2(n637), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT85), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT2), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n634), .A2(G48), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(G305) );
  NAND2_X1 U701 ( .A1(G49), .A2(n634), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U704 ( .A(KEYINPUT82), .B(n626), .ZN(n627) );
  NOR2_X1 U705 ( .A1(n633), .A2(n627), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U708 ( .A1(G88), .A2(n631), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT86), .ZN(n642) );
  NAND2_X1 U710 ( .A1(G62), .A2(n633), .ZN(n636) );
  NAND2_X1 U711 ( .A1(G50), .A2(n634), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G75), .A2(n637), .ZN(n638) );
  XNOR2_X1 U714 ( .A(KEYINPUT87), .B(n638), .ZN(n639) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(G303) );
  INV_X1 U717 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U718 ( .A(KEYINPUT91), .B(KEYINPUT88), .ZN(n644) );
  XNOR2_X1 U719 ( .A(G288), .B(KEYINPUT19), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U721 ( .A(KEYINPUT89), .B(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(G290), .B(KEYINPUT90), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U724 ( .A(G305), .B(n648), .ZN(n650) );
  INV_X1 U725 ( .A(G299), .ZN(n964) );
  XNOR2_X1 U726 ( .A(n964), .B(G166), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U728 ( .A(n655), .B(n651), .Z(n838) );
  XNOR2_X1 U729 ( .A(n652), .B(n838), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n653), .A2(G868), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U733 ( .A(KEYINPUT92), .B(n658), .Z(G295) );
  NAND2_X1 U734 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n662), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U740 ( .A1(G220), .A2(G219), .ZN(n663) );
  XOR2_X1 U741 ( .A(KEYINPUT22), .B(n663), .Z(n664) );
  NOR2_X1 U742 ( .A1(G218), .A2(n664), .ZN(n665) );
  NAND2_X1 U743 ( .A1(G96), .A2(n665), .ZN(n826) );
  NAND2_X1 U744 ( .A1(n826), .A2(G2106), .ZN(n669) );
  NAND2_X1 U745 ( .A1(G108), .A2(G120), .ZN(n666) );
  NOR2_X1 U746 ( .A1(G237), .A2(n666), .ZN(n667) );
  NAND2_X1 U747 ( .A1(G69), .A2(n667), .ZN(n827) );
  NAND2_X1 U748 ( .A1(n827), .A2(G567), .ZN(n668) );
  NAND2_X1 U749 ( .A1(n669), .A2(n668), .ZN(n903) );
  NAND2_X1 U750 ( .A1(G661), .A2(G483), .ZN(n670) );
  NOR2_X1 U751 ( .A1(n903), .A2(n670), .ZN(n671) );
  XOR2_X1 U752 ( .A(KEYINPUT93), .B(n671), .Z(n825) );
  NAND2_X1 U753 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U754 ( .A1(G126), .A2(n881), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n672), .B(KEYINPUT94), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G114), .A2(n882), .ZN(n673) );
  XOR2_X1 U757 ( .A(KEYINPUT95), .B(n673), .Z(n674) );
  NAND2_X1 U758 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U759 ( .A1(G138), .A2(n877), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G102), .A2(n878), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U762 ( .A1(n679), .A2(n678), .ZN(G164) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n695) );
  AND2_X1 U764 ( .A1(n680), .A2(G40), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n682), .A2(n681), .ZN(n693) );
  NOR2_X1 U766 ( .A1(n695), .A2(n693), .ZN(n817) );
  XNOR2_X1 U767 ( .A(G2067), .B(KEYINPUT37), .ZN(n683) );
  XNOR2_X1 U768 ( .A(n683), .B(KEYINPUT96), .ZN(n815) );
  NAND2_X1 U769 ( .A1(G140), .A2(n877), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G104), .A2(n878), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n686), .ZN(n691) );
  NAND2_X1 U773 ( .A1(G128), .A2(n881), .ZN(n688) );
  NAND2_X1 U774 ( .A1(G116), .A2(n882), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U776 ( .A(KEYINPUT35), .B(n689), .Z(n690) );
  NOR2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U778 ( .A(KEYINPUT36), .B(n692), .ZN(n895) );
  NOR2_X1 U779 ( .A1(n815), .A2(n895), .ZN(n921) );
  NAND2_X1 U780 ( .A1(n817), .A2(n921), .ZN(n813) );
  INV_X1 U781 ( .A(n813), .ZN(n781) );
  INV_X1 U782 ( .A(n693), .ZN(n694) );
  INV_X2 U783 ( .A(n735), .ZN(n721) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n721), .ZN(n696) );
  XOR2_X1 U785 ( .A(KEYINPUT26), .B(n696), .Z(n697) );
  NAND2_X1 U786 ( .A1(G1341), .A2(n735), .ZN(n698) );
  NAND2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n710) );
  XOR2_X1 U788 ( .A(n700), .B(KEYINPUT104), .Z(n708) );
  NOR2_X1 U789 ( .A1(n721), .A2(G1348), .ZN(n702) );
  NOR2_X1 U790 ( .A1(G2067), .A2(n735), .ZN(n701) );
  NOR2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U792 ( .A1(n721), .A2(G2072), .ZN(n703) );
  XNOR2_X1 U793 ( .A(n703), .B(KEYINPUT27), .ZN(n705) );
  XOR2_X1 U794 ( .A(G1956), .B(KEYINPUT102), .Z(n987) );
  NOR2_X1 U795 ( .A1(n721), .A2(n987), .ZN(n704) );
  NOR2_X1 U796 ( .A1(n705), .A2(n704), .ZN(n713) );
  NAND2_X1 U797 ( .A1(n964), .A2(n713), .ZN(n709) );
  AND2_X1 U798 ( .A1(n706), .A2(n709), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n719) );
  INV_X1 U800 ( .A(n709), .ZN(n712) );
  NAND2_X1 U801 ( .A1(n710), .A2(n971), .ZN(n711) );
  OR2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U803 ( .A1(n964), .A2(n713), .ZN(n715) );
  XNOR2_X1 U804 ( .A(KEYINPUT28), .B(KEYINPUT103), .ZN(n714) );
  XNOR2_X1 U805 ( .A(n715), .B(n714), .ZN(n716) );
  AND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U808 ( .A(n720), .B(KEYINPUT29), .ZN(n725) );
  XNOR2_X1 U809 ( .A(KEYINPUT25), .B(G2078), .ZN(n940) );
  NOR2_X1 U810 ( .A1(n735), .A2(n940), .ZN(n723) );
  INV_X1 U811 ( .A(G1961), .ZN(n986) );
  NOR2_X1 U812 ( .A1(n721), .A2(n986), .ZN(n722) );
  NOR2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n731) );
  AND2_X1 U814 ( .A1(G171), .A2(n731), .ZN(n724) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U816 ( .A(n726), .B(KEYINPUT105), .ZN(n750) );
  NAND2_X1 U817 ( .A1(G8), .A2(n735), .ZN(n774) );
  NOR2_X1 U818 ( .A1(G1966), .A2(n774), .ZN(n752) );
  NOR2_X1 U819 ( .A1(G2084), .A2(n735), .ZN(n748) );
  NOR2_X1 U820 ( .A1(n752), .A2(n748), .ZN(n727) );
  NAND2_X1 U821 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U822 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  XNOR2_X1 U823 ( .A(KEYINPUT106), .B(n729), .ZN(n730) );
  NOR2_X1 U824 ( .A1(G168), .A2(n730), .ZN(n733) );
  NOR2_X1 U825 ( .A1(G171), .A2(n731), .ZN(n732) );
  NOR2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U827 ( .A(KEYINPUT31), .B(n734), .Z(n749) );
  INV_X1 U828 ( .A(G8), .ZN(n741) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n774), .ZN(n737) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U832 ( .A(KEYINPUT107), .B(n738), .Z(n739) );
  NAND2_X1 U833 ( .A1(n739), .A2(G303), .ZN(n740) );
  OR2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n743) );
  AND2_X1 U835 ( .A1(n749), .A2(n743), .ZN(n742) );
  NAND2_X1 U836 ( .A1(n750), .A2(n742), .ZN(n746) );
  INV_X1 U837 ( .A(n743), .ZN(n744) );
  OR2_X1 U838 ( .A1(n744), .A2(G286), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U840 ( .A(n747), .B(KEYINPUT32), .ZN(n756) );
  NAND2_X1 U841 ( .A1(G8), .A2(n748), .ZN(n754) );
  AND2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n773) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n762) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n762), .A2(n757), .ZN(n965) );
  INV_X1 U849 ( .A(KEYINPUT33), .ZN(n758) );
  AND2_X1 U850 ( .A1(n965), .A2(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n773), .A2(n759), .ZN(n767) );
  INV_X1 U852 ( .A(n774), .ZN(n760) );
  NAND2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n967) );
  AND2_X1 U854 ( .A1(n760), .A2(n967), .ZN(n761) );
  NOR2_X1 U855 ( .A1(KEYINPUT33), .A2(n761), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n762), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U857 ( .A1(n763), .A2(n774), .ZN(n764) );
  NOR2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n766) );
  AND2_X1 U859 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U860 ( .A(G1981), .B(G305), .Z(n961) );
  NAND2_X1 U861 ( .A1(n768), .A2(n961), .ZN(n779) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U863 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  NOR2_X1 U864 ( .A1(n774), .A2(n770), .ZN(n777) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U866 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U867 ( .A1(n773), .A2(n772), .ZN(n775) );
  AND2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  AND2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n805) );
  NAND2_X1 U872 ( .A1(n878), .A2(G105), .ZN(n782) );
  XNOR2_X1 U873 ( .A(KEYINPUT38), .B(n782), .ZN(n788) );
  NAND2_X1 U874 ( .A1(n881), .A2(G129), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT99), .B(n783), .Z(n785) );
  NAND2_X1 U876 ( .A1(n882), .A2(G117), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U878 ( .A(KEYINPUT100), .B(n786), .Z(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U880 ( .A(n789), .B(KEYINPUT101), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G141), .A2(n877), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n898) );
  NAND2_X1 U883 ( .A1(n898), .A2(G1996), .ZN(n801) );
  NAND2_X1 U884 ( .A1(G131), .A2(n877), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G95), .A2(n878), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U887 ( .A(KEYINPUT98), .B(n794), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G119), .A2(n881), .ZN(n795) );
  XNOR2_X1 U889 ( .A(KEYINPUT97), .B(n795), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n882), .A2(G107), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n890) );
  NAND2_X1 U893 ( .A1(n890), .A2(G1991), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n917) );
  INV_X1 U895 ( .A(n917), .ZN(n802) );
  XOR2_X1 U896 ( .A(G1986), .B(G290), .Z(n968) );
  NAND2_X1 U897 ( .A1(n802), .A2(n968), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n803), .A2(n817), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n820) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n898), .ZN(n912) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n890), .ZN(n915) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n806) );
  XNOR2_X1 U903 ( .A(KEYINPUT108), .B(n806), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n915), .A2(n807), .ZN(n808) );
  XOR2_X1 U905 ( .A(KEYINPUT109), .B(n808), .Z(n809) );
  NOR2_X1 U906 ( .A1(n917), .A2(n809), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n810), .B(KEYINPUT110), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n912), .A2(n811), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n815), .A2(n895), .ZN(n926) );
  NAND2_X1 U912 ( .A1(n816), .A2(n926), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U915 ( .A(KEYINPUT40), .B(n821), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U918 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U921 ( .A(G120), .B(KEYINPUT113), .ZN(G236) );
  XOR2_X1 U922 ( .A(G96), .B(KEYINPUT114), .Z(G221) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  NOR2_X1 U925 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U927 ( .A(G1348), .B(G2454), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n828), .B(G2430), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n829), .B(G1341), .ZN(n835) );
  XOR2_X1 U930 ( .A(G2443), .B(G2427), .Z(n831) );
  XNOR2_X1 U931 ( .A(G2438), .B(G2446), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n833) );
  XOR2_X1 U933 ( .A(G2451), .B(G2435), .Z(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U936 ( .A1(n836), .A2(G14), .ZN(n837) );
  XOR2_X1 U937 ( .A(KEYINPUT111), .B(n837), .Z(n906) );
  XOR2_X1 U938 ( .A(KEYINPUT112), .B(n906), .Z(G401) );
  XNOR2_X1 U939 ( .A(n838), .B(n971), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n839), .B(n979), .ZN(n841) );
  XOR2_X1 U941 ( .A(G286), .B(G171), .Z(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  NOR2_X1 U943 ( .A1(G37), .A2(n842), .ZN(G397) );
  XOR2_X1 U944 ( .A(G2096), .B(G2100), .Z(n844) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2090), .Z(n846) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U950 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U953 ( .A(G1976), .B(G1971), .Z(n852) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1961), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U959 ( .A(G2474), .B(G1981), .Z(n857) );
  XNOR2_X1 U960 ( .A(G1966), .B(G1956), .ZN(n856) );
  XNOR2_X1 U961 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G100), .A2(n878), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G112), .A2(n882), .ZN(n861) );
  NAND2_X1 U965 ( .A1(G136), .A2(n877), .ZN(n860) );
  NAND2_X1 U966 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n881), .A2(G124), .ZN(n862) );
  XOR2_X1 U968 ( .A(KEYINPUT44), .B(n862), .Z(n863) );
  NOR2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n867), .B(KEYINPUT115), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G130), .A2(n881), .ZN(n869) );
  NAND2_X1 U973 ( .A1(G118), .A2(n882), .ZN(n868) );
  NAND2_X1 U974 ( .A1(n869), .A2(n868), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G142), .A2(n877), .ZN(n871) );
  NAND2_X1 U976 ( .A1(G106), .A2(n878), .ZN(n870) );
  NAND2_X1 U977 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U978 ( .A(KEYINPUT116), .B(n872), .Z(n873) );
  XNOR2_X1 U979 ( .A(KEYINPUT45), .B(n873), .ZN(n874) );
  NOR2_X1 U980 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U981 ( .A(n876), .B(G162), .Z(n889) );
  NAND2_X1 U982 ( .A1(G139), .A2(n877), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G103), .A2(n878), .ZN(n879) );
  NAND2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G127), .A2(n881), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G115), .A2(n882), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n928) );
  XNOR2_X1 U990 ( .A(G164), .B(n928), .ZN(n888) );
  XNOR2_X1 U991 ( .A(n889), .B(n888), .ZN(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n890), .B(KEYINPUT117), .ZN(n891) );
  XNOR2_X1 U994 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n895), .B(n914), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n898), .B(G160), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n901), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(KEYINPUT118), .B(n902), .ZN(G395) );
  INV_X1 U1002 ( .A(n903), .ZN(G319) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1005 ( .A1(G397), .A2(n905), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(n906), .A2(G319), .ZN(n907) );
  XOR2_X1 U1007 ( .A(KEYINPUT119), .B(n907), .Z(n908) );
  NOR2_X1 U1008 ( .A1(G395), .A2(n908), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1012 ( .A(G2090), .B(G162), .Z(n911) );
  NOR2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1014 ( .A(KEYINPUT51), .B(n913), .Z(n924) );
  NOR2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n919) );
  XOR2_X1 U1016 ( .A(G160), .B(G2084), .Z(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT120), .B(n922), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n925), .B(KEYINPUT121), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1024 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n931), .Z(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n934), .ZN(n935) );
  XOR2_X1 U1030 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n957) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n957), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n936), .A2(G29), .ZN(n937) );
  XOR2_X1 U1033 ( .A(KEYINPUT123), .B(n937), .Z(n1016) );
  XNOR2_X1 U1034 ( .A(G1991), .B(G25), .ZN(n948) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G1996), .B(G32), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G27), .B(KEYINPUT124), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(n941), .B(n940), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT125), .B(n946), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(G28), .A2(n949), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(n950), .B(KEYINPUT53), .ZN(n953) );
  XOR2_X1 U1047 ( .A(G2084), .B(G34), .Z(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT54), .B(n951), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G35), .B(G2090), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1052 ( .A(n957), .B(n956), .Z(n959) );
  INV_X1 U1053 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n960), .A2(G11), .ZN(n1014) );
  XNOR2_X1 U1056 ( .A(G16), .B(KEYINPUT56), .ZN(n985) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G168), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n963), .B(KEYINPUT57), .ZN(n983) );
  XNOR2_X1 U1060 ( .A(n964), .B(G1956), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n977) );
  AND2_X1 U1062 ( .A1(G303), .A2(G1971), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(G301), .B(G1961), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n971), .B(G1348), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1070 ( .A(KEYINPUT126), .B(n978), .Z(n981) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n979), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n1012) );
  INV_X1 U1075 ( .A(G16), .ZN(n1010) );
  XNOR2_X1 U1076 ( .A(G5), .B(n986), .ZN(n1005) );
  XNOR2_X1 U1077 ( .A(n987), .B(G20), .ZN(n995) );
  XNOR2_X1 U1078 ( .A(KEYINPUT59), .B(G1348), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n988), .B(G4), .ZN(n990) );
  XOR2_X1 U1080 ( .A(G1341), .B(G19), .Z(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1082 ( .A(KEYINPUT127), .B(G1981), .Z(n991) );
  XNOR2_X1 U1083 ( .A(G6), .B(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n996), .B(KEYINPUT60), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(G23), .B(G1976), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XOR2_X1 U1090 ( .A(G1986), .B(G24), .Z(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT58), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G21), .B(G1966), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT61), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1017), .Z(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

