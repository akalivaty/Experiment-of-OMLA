//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT66), .A2(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT66), .A2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(G131), .B1(new_n191), .B2(G137), .ZN(new_n196));
  OAI211_X1 g010(.A(KEYINPUT65), .B(new_n190), .C1(new_n191), .C2(G137), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G134), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT65), .B1(new_n200), .B2(new_n190), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n195), .B(new_n196), .C1(new_n198), .C2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(G134), .B1(new_n193), .B2(new_n194), .ZN(new_n203));
  INV_X1    g017(.A(new_n200), .ZN(new_n204));
  OAI21_X1  g018(.A(G131), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  OAI211_X1 g025(.A(G128), .B(new_n208), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(G146), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n213), .B(new_n214), .C1(KEYINPUT1), .C2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n216), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT0), .A4(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n209), .B2(new_n211), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n223), .B2(KEYINPUT64), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n222), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n191), .A2(G137), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n195), .B(new_n229), .C1(new_n198), .C2(new_n201), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n228), .B1(new_n231), .B2(new_n202), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n189), .B1(new_n221), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n228), .ZN(new_n237));
  INV_X1    g051(.A(G131), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT65), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT66), .A2(G137), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT66), .A2(G137), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n241), .A2(new_n197), .B1(new_n244), .B2(new_n192), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n238), .B1(new_n245), .B2(new_n229), .ZN(new_n246));
  INV_X1    g060(.A(new_n202), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n237), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n217), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT68), .B1(new_n212), .B2(new_n216), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n202), .B(new_n205), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n251), .A3(KEYINPUT71), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n233), .A2(new_n236), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n251), .A3(new_n236), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n236), .B1(new_n248), .B2(new_n251), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n255), .B1(new_n259), .B2(new_n254), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT69), .B(G237), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(G210), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT29), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n188), .B1(new_n260), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n236), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n212), .A2(new_n216), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n271), .A2(KEYINPUT67), .A3(new_n202), .A4(new_n205), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n230), .A2(G131), .B1(new_n245), .B2(new_n196), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n228), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n200), .B1(new_n244), .B2(G134), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n245), .A2(new_n196), .B1(new_n275), .B2(G131), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT67), .B1(new_n276), .B2(new_n271), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n270), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n256), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n255), .A3(new_n267), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n280), .A2(new_n255), .A3(KEYINPUT72), .A4(new_n267), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n274), .B2(new_n277), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n248), .A2(new_n251), .A3(KEYINPUT30), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n270), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n256), .ZN(new_n289));
  INV_X1    g103(.A(new_n267), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n283), .A2(new_n284), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n269), .B1(new_n292), .B2(KEYINPUT73), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n283), .A2(new_n294), .A3(new_n284), .A4(new_n291), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n187), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n288), .A2(new_n256), .A3(new_n267), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT31), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n256), .A4(new_n267), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n280), .A2(new_n255), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n290), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n297), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n300), .A2(new_n301), .B1(new_n303), .B2(new_n290), .ZN(new_n308));
  INV_X1    g122(.A(new_n306), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n308), .A2(KEYINPUT32), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT74), .B1(new_n296), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n291), .A2(new_n284), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n249), .A2(new_n250), .ZN(new_n314));
  OAI22_X1  g128(.A1(new_n314), .A2(new_n206), .B1(new_n273), .B2(new_n228), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n270), .B1(new_n315), .B2(new_n189), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT28), .B1(new_n316), .B2(new_n252), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n254), .B1(new_n278), .B2(new_n256), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT72), .B1(new_n319), .B2(new_n267), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT73), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n269), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n295), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G472), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n305), .A2(new_n297), .A3(new_n306), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT32), .B1(new_n308), .B2(new_n309), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n215), .A2(G119), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G128), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n331), .B2(G128), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n330), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n340), .A3(new_n332), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT76), .B1(new_n341), .B2(G110), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n341), .A2(KEYINPUT76), .A3(G110), .ZN(new_n343));
  XNOR2_X1  g157(.A(G125), .B(G140), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G125), .ZN(new_n347));
  OR3_X1    g161(.A1(new_n345), .A2(new_n347), .A3(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(KEYINPUT16), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT16), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n347), .B2(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(G146), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n210), .B1(new_n349), .B2(new_n351), .ZN(new_n354));
  OAI221_X1 g168(.A(new_n335), .B1(new_n342), .B2(new_n343), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n354), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n344), .B(KEYINPUT79), .Z(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n210), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT78), .B(G110), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n341), .A2(new_n359), .B1(new_n333), .B2(new_n334), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G137), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n362), .B(new_n363), .Z(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n355), .B2(new_n361), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT80), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n355), .A2(new_n361), .ZN(new_n369));
  INV_X1    g183(.A(new_n364), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n365), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(G234), .B2(new_n188), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(G902), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT81), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n379));
  INV_X1    g193(.A(new_n377), .ZN(new_n380));
  AOI211_X1 g194(.A(new_n379), .B(new_n380), .C1(new_n368), .C2(new_n373), .ZN(new_n381));
  INV_X1    g195(.A(new_n376), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(new_n188), .A3(new_n365), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT25), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n371), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n365), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n378), .A2(new_n381), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n312), .A2(new_n329), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G469), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G104), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT82), .B(KEYINPUT3), .C1(new_n393), .C2(KEYINPUT83), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n392), .A2(G104), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n397));
  INV_X1    g211(.A(G104), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G107), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n399), .B2(new_n397), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n394), .B(new_n396), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n405), .A3(G101), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT82), .B1(new_n393), .B2(KEYINPUT83), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n393), .B2(KEYINPUT82), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G101), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n394), .A4(new_n396), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT4), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n395), .B1(new_n407), .B2(new_n408), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n410), .B1(new_n413), .B2(new_n394), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n237), .B(new_n406), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT10), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n220), .B2(new_n217), .ZN(new_n417));
  OAI21_X1  g231(.A(G101), .B1(new_n399), .B2(new_n395), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n411), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n411), .A2(new_n271), .A3(new_n418), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n415), .A2(new_n420), .A3(new_n423), .A4(new_n273), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n228), .B1(new_n414), .B2(new_n405), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n404), .A2(G101), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT4), .A3(new_n411), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n426), .A2(new_n428), .B1(new_n417), .B2(new_n419), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n273), .A4(new_n423), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G140), .ZN(new_n433));
  INV_X1    g247(.A(G227), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G953), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n429), .A2(new_n423), .ZN(new_n438));
  INV_X1    g252(.A(new_n273), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n442));
  INV_X1    g256(.A(new_n421), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n271), .B1(new_n411), .B2(new_n418), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n439), .B(new_n442), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n444), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n273), .B1(new_n446), .B2(new_n421), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT12), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n425), .B2(new_n431), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n441), .B1(new_n437), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n391), .B1(new_n452), .B2(new_n188), .ZN(new_n453));
  INV_X1    g267(.A(new_n450), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n432), .A2(new_n437), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n432), .A2(new_n440), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n455), .A2(new_n456), .B1(new_n457), .B2(new_n436), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n451), .A2(KEYINPUT87), .A3(new_n437), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n453), .B1(new_n460), .B2(new_n391), .ZN(new_n461));
  AND2_X1   g275(.A1(KEYINPUT69), .A2(G237), .ZN(new_n462));
  NOR2_X1   g276(.A1(KEYINPUT69), .A2(G237), .ZN(new_n463));
  OAI211_X1 g277(.A(G214), .B(new_n262), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n207), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n261), .A2(G143), .A3(G214), .A4(new_n262), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G131), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT17), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(KEYINPUT94), .A3(G131), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n238), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n470), .A2(new_n471), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n353), .A2(new_n354), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT94), .B1(new_n467), .B2(G131), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n469), .B(new_n238), .C1(new_n465), .C2(new_n466), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT17), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G113), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n398), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n346), .A2(new_n348), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G146), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n358), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n473), .B1(new_n486), .B2(new_n238), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n467), .A2(KEYINPUT18), .A3(G131), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n482), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT95), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n480), .A2(KEYINPUT95), .A3(new_n482), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n470), .A2(new_n472), .A3(new_n474), .ZN(new_n495));
  MUX2_X1   g309(.A(new_n357), .B(new_n483), .S(KEYINPUT19), .Z(new_n496));
  OAI211_X1 g310(.A(new_n495), .B(new_n356), .C1(new_n496), .C2(G146), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n489), .ZN(new_n498));
  INV_X1    g312(.A(new_n482), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n492), .A2(new_n493), .B1(new_n499), .B2(new_n498), .ZN(new_n505));
  INV_X1    g319(.A(new_n503), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT20), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G122), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT96), .B1(new_n509), .B2(G116), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT96), .ZN(new_n511));
  INV_X1    g325(.A(G116), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(G122), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n512), .B2(G122), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(G107), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n207), .A2(G128), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n215), .A2(G143), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(new_n191), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G134), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n514), .A2(KEYINPUT14), .B1(G116), .B2(new_n509), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(KEYINPUT14), .B2(new_n514), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G107), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT97), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n517), .B2(new_n527), .ZN(new_n529));
  AOI211_X1 g343(.A(KEYINPUT97), .B(KEYINPUT13), .C1(new_n207), .C2(G128), .ZN(new_n530));
  OAI221_X1 g344(.A(new_n518), .B1(new_n527), .B2(new_n517), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G134), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n515), .A2(G107), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n532), .B(new_n519), .C1(new_n533), .C2(new_n516), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT9), .B(G234), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n536), .A2(new_n375), .A3(G953), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n526), .A2(new_n534), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n188), .ZN(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n542), .B(new_n544), .Z(new_n545));
  AOI21_X1  g359(.A(new_n482), .B1(new_n480), .B2(new_n489), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n492), .B2(new_n493), .ZN(new_n547));
  OAI21_X1  g361(.A(G475), .B1(new_n547), .B2(G902), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n508), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G221), .B1(new_n536), .B2(G902), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n461), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(G234), .A2(G237), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(G952), .A3(new_n262), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT21), .B(G898), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(G902), .A3(G953), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G214), .B1(G237), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G210), .B1(G237), .B2(G902), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT93), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n234), .A2(KEYINPUT5), .ZN(new_n566));
  INV_X1    g380(.A(G113), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n512), .A2(G119), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT5), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n566), .A2(KEYINPUT88), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT88), .B1(new_n566), .B2(new_n570), .ZN(new_n572));
  INV_X1    g386(.A(new_n234), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n235), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n411), .A2(new_n418), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n566), .A2(new_n570), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n411), .B(new_n418), .C1(new_n574), .C2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(G110), .B(G122), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT8), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n212), .A2(new_n347), .A3(new_n216), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n228), .B2(new_n347), .ZN(new_n584));
  INV_X1    g398(.A(G224), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT7), .B1(new_n585), .B2(G953), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n584), .B(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n582), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n582), .B2(new_n587), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n270), .B(new_n406), .C1(new_n412), .C2(new_n414), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n419), .A2(new_n575), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n580), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT89), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n236), .B1(new_n414), .B2(new_n405), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n597), .A2(new_n428), .B1(new_n419), .B2(new_n575), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(KEYINPUT89), .A3(new_n580), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n591), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n592), .A2(new_n593), .ZN(new_n602));
  INV_X1    g416(.A(new_n580), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT6), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT89), .B1(new_n598), .B2(new_n580), .ZN(new_n607));
  AND4_X1   g421(.A1(KEYINPUT89), .A2(new_n592), .A3(new_n580), .A4(new_n593), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT6), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n609), .B2(new_n604), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n585), .A2(G953), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT90), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n584), .B(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n601), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n565), .B1(new_n615), .B2(KEYINPUT92), .ZN(new_n616));
  INV_X1    g430(.A(new_n606), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n605), .B1(new_n596), .B2(new_n599), .ZN(new_n618));
  INV_X1    g432(.A(new_n604), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n613), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT92), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n601), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n564), .B(new_n601), .C1(new_n610), .C2(new_n614), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n563), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n552), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n390), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT98), .B(G101), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G3));
  OAI21_X1  g444(.A(G472), .B1(new_n308), .B2(G902), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n308), .B2(new_n309), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n388), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n455), .A2(new_n456), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n457), .A2(new_n436), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n459), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n391), .A3(new_n188), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n432), .A2(new_n437), .A3(new_n440), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n437), .B1(new_n432), .B2(new_n454), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(G469), .B1(new_n640), .B2(G902), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n551), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT99), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n502), .B1(new_n501), .B2(new_n503), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n505), .A2(KEYINPUT20), .A3(new_n506), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n548), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT102), .B(G478), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n542), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n541), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT100), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n541), .A2(new_n653), .A3(new_n650), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n540), .A2(KEYINPUT101), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n540), .A2(KEYINPUT101), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(KEYINPUT33), .A3(new_n656), .A4(new_n539), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n652), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n188), .A2(G478), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n649), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n647), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n625), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n564), .B1(new_n621), .B2(new_n601), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n558), .B(new_n560), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n644), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT103), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  INV_X1    g483(.A(new_n545), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n508), .A2(new_n670), .A3(new_n548), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n644), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT35), .B(G107), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  NOR2_X1   g489(.A1(new_n370), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n369), .B(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n677), .A2(new_n377), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n387), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n632), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n549), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n626), .A2(new_n680), .A3(new_n681), .A4(new_n642), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT37), .B(G110), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G12));
  NAND2_X1  g498(.A1(new_n637), .A2(new_n641), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n550), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n387), .A2(new_n678), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n687), .B(new_n560), .C1(new_n662), .C2(new_n663), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n557), .A2(G900), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n554), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n671), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n689), .A2(new_n312), .A3(new_n329), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  NAND2_X1  g509(.A1(new_n624), .A2(new_n625), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n691), .B(KEYINPUT39), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n642), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n647), .A2(new_n670), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n290), .B1(new_n257), .B2(new_n258), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n298), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n188), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n326), .A2(new_n327), .B1(G472), .B2(new_n709), .ZN(new_n710));
  NOR4_X1   g524(.A1(new_n703), .A2(new_n710), .A3(new_n561), .A4(new_n687), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n698), .A2(new_n701), .A3(new_n702), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND2_X1  g527(.A1(new_n312), .A2(new_n329), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n647), .A2(new_n660), .A3(new_n691), .ZN(new_n715));
  INV_X1    g529(.A(new_n564), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n615), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n561), .B1(new_n717), .B2(new_n625), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(new_n642), .A3(new_n718), .A4(new_n687), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n210), .ZN(G48));
  NAND2_X1  g535(.A1(new_n636), .A2(new_n188), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(G469), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n550), .A3(new_n637), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n723), .A2(KEYINPUT106), .A3(new_n550), .A4(new_n637), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n665), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n390), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT41), .B(G113), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n726), .A2(new_n672), .A3(new_n727), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n390), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n512), .ZN(G18));
  AND3_X1   g548(.A1(new_n726), .A2(new_n718), .A3(new_n727), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n549), .A2(new_n559), .A3(new_n679), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n312), .A2(new_n329), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n737), .A3(KEYINPUT107), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n726), .A2(new_n718), .A3(new_n727), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n312), .A2(new_n329), .A3(new_n736), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G119), .ZN(G21));
  OAI21_X1  g558(.A(new_n560), .B1(new_n662), .B2(new_n663), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n703), .A2(new_n745), .A3(new_n559), .ZN(new_n746));
  INV_X1    g560(.A(new_n260), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n302), .B1(new_n747), .B2(new_n267), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n306), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT108), .B(G472), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n308), .B2(G902), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n388), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n746), .A2(new_n726), .A3(new_n727), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  NAND3_X1  g569(.A1(new_n647), .A2(new_n660), .A3(new_n691), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n687), .A2(new_n749), .A3(new_n751), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n726), .A2(new_n758), .A3(new_n718), .A4(new_n727), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  AOI21_X1  g574(.A(new_n551), .B1(new_n685), .B2(KEYINPUT109), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n561), .B(new_n662), .C1(new_n616), .C2(new_n623), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n637), .A2(new_n763), .A3(new_n641), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n390), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT42), .B1(new_n766), .B2(new_n715), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n324), .A2(new_n328), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n715), .A3(KEYINPUT42), .A4(new_n389), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT110), .B1(new_n769), .B2(new_n765), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n323), .A2(G472), .B1(new_n327), .B2(new_n326), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n647), .A2(KEYINPUT42), .A3(new_n660), .A4(new_n691), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n771), .A2(new_n772), .A3(new_n388), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n685), .A2(KEYINPUT109), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n550), .A3(new_n764), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n773), .A2(new_n775), .A3(new_n776), .A4(new_n762), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n767), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT111), .B(G131), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(G33));
  NAND2_X1  g595(.A1(new_n766), .A2(new_n693), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  NAND2_X1  g597(.A1(new_n632), .A2(new_n687), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT112), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n508), .A2(new_n548), .A3(new_n660), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT43), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n786), .A2(KEYINPUT43), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT44), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n640), .A2(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n640), .A2(KEYINPUT45), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(G469), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(G469), .A2(G902), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(KEYINPUT46), .A3(new_n794), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n637), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n550), .A3(new_n699), .ZN(new_n800));
  INV_X1    g614(.A(new_n762), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  AND3_X1   g618(.A1(new_n799), .A2(KEYINPUT47), .A3(new_n550), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT47), .B1(new_n799), .B2(new_n550), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n801), .A2(new_n389), .A3(new_n756), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n714), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND2_X1  g625(.A1(new_n723), .A2(new_n637), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n550), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n753), .ZN(new_n815));
  INV_X1    g629(.A(new_n554), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n788), .A2(new_n816), .A3(new_n787), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT116), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(KEYINPUT116), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n762), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT51), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n726), .A2(new_n727), .A3(new_n762), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n389), .A2(new_n816), .A3(new_n710), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n647), .A3(new_n660), .ZN(new_n826));
  INV_X1    g640(.A(new_n757), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n823), .B1(new_n818), .B2(new_n819), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n698), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n561), .A2(new_n830), .A3(new_n726), .A4(new_n727), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n831), .A2(KEYINPUT50), .A3(new_n820), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT50), .B1(new_n831), .B2(new_n820), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n834), .A2(KEYINPUT118), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(KEYINPUT118), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n822), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n807), .A2(KEYINPUT117), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n813), .B1(new_n807), .B2(KEYINPUT117), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n821), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n771), .A2(new_n388), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n828), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT119), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n828), .A2(new_n846), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT120), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n845), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n851), .A3(KEYINPUT48), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n262), .A2(G952), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n825), .A2(new_n661), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n853), .B(new_n854), .C1(new_n735), .C2(new_n820), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT48), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n848), .A2(KEYINPUT120), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n842), .A2(new_n852), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n837), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n661), .A2(new_n671), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n626), .A2(new_n860), .A3(new_n633), .A4(new_n642), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n682), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n628), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n679), .A2(new_n692), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n625), .A2(new_n624), .A3(new_n560), .A4(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n312), .A3(new_n552), .A4(new_n329), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n758), .A2(new_n762), .A3(new_n764), .A4(new_n761), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n782), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n779), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n694), .A2(new_n759), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n312), .A2(new_n329), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n686), .A2(new_n688), .A3(new_n756), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n718), .A2(new_n670), .A3(new_n647), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n679), .A2(new_n691), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n710), .A3(new_n876), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n873), .A2(new_n874), .B1(new_n877), .B2(new_n775), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT115), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n694), .A2(new_n759), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n703), .A2(new_n745), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n709), .A2(G472), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n876), .B1(new_n328), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n881), .A2(new_n761), .A3(new_n764), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n714), .B2(new_n719), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n871), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT52), .B1(new_n880), .B2(new_n885), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n754), .B1(new_n390), .B2(new_n728), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n733), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n891), .A2(new_n743), .A3(KEYINPUT53), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n870), .A2(new_n888), .A3(new_n889), .A4(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n891), .A2(new_n743), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n891), .B2(new_n743), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n872), .A2(new_n878), .A3(KEYINPUT115), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(KEYINPUT52), .A3(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n897), .A2(new_n870), .A3(new_n888), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT53), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n893), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n891), .A2(new_n743), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT114), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n891), .A2(new_n743), .A3(new_n894), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n870), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n888), .A2(new_n889), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n901), .A2(KEYINPUT53), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT54), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n859), .A2(new_n914), .B1(G952), .B2(G953), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n812), .A2(KEYINPUT49), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT113), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n812), .A2(KEYINPUT49), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n786), .A2(new_n561), .A3(new_n551), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n389), .A2(new_n918), .A3(new_n919), .A4(new_n710), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n830), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n915), .A2(new_n921), .ZN(G75));
  XNOR2_X1  g736(.A(new_n620), .B(new_n614), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT55), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n888), .A2(new_n900), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n902), .B1(new_n909), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n870), .A2(new_n888), .A3(new_n889), .A4(new_n892), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(G902), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(G210), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n924), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n262), .A2(G952), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n929), .A2(new_n565), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n924), .A2(new_n932), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n933), .A2(new_n938), .ZN(G51));
  XOR2_X1   g753(.A(new_n794), .B(KEYINPUT57), .Z(new_n940));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n926), .A2(new_n941), .A3(new_n904), .A4(new_n927), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n903), .B2(new_n904), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n903), .B2(new_n904), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n636), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n929), .A2(new_n793), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n934), .B1(new_n946), .B2(new_n947), .ZN(G54));
  NAND2_X1  g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n505), .B1(new_n929), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n935), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n929), .A2(new_n505), .A3(new_n949), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(G60));
  NOR2_X1   g767(.A1(new_n943), .A2(new_n944), .ZN(new_n954));
  NAND2_X1  g768(.A1(G478), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT59), .Z(new_n956));
  OR2_X1    g770(.A1(new_n658), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n905), .B2(new_n913), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n652), .A2(new_n654), .A3(new_n657), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n935), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(G63));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT123), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT122), .Z(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT60), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n926), .B2(new_n927), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n677), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n935), .B1(new_n970), .B2(new_n374), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n964), .B(new_n965), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n928), .A2(new_n968), .ZN(new_n975));
  INV_X1    g789(.A(new_n374), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n934), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(KEYINPUT123), .A3(new_n963), .A4(new_n971), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n974), .A2(new_n978), .ZN(G66));
  AOI21_X1  g793(.A(new_n262), .B1(new_n556), .B2(G224), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n897), .A2(new_n863), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n262), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n610), .B1(G898), .B2(new_n262), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT124), .Z(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  XOR2_X1   g799(.A(new_n496), .B(KEYINPUT125), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n286), .A2(new_n287), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n810), .A2(new_n803), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n880), .A2(new_n720), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n712), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n762), .A2(new_n860), .ZN(new_n994));
  OR3_X1    g808(.A1(new_n390), .A2(new_n700), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n989), .A2(new_n992), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n988), .B1(new_n996), .B2(new_n262), .ZN(new_n997));
  INV_X1    g811(.A(new_n779), .ZN(new_n998));
  NOR4_X1   g812(.A1(new_n800), .A2(new_n771), .A3(new_n388), .A4(new_n875), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n693), .B2(new_n766), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n989), .A2(new_n998), .A3(new_n990), .A4(new_n1000), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n1001), .A2(G953), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G900), .A2(G953), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n988), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n997), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(G900), .ZN(new_n1006));
  OAI21_X1  g820(.A(G953), .B1(new_n434), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1005), .B(new_n1007), .ZN(G72));
  XNOR2_X1  g822(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n187), .A2(new_n188), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(new_n1001), .B2(new_n981), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n289), .B(KEYINPUT127), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1013), .A2(new_n267), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n934), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n289), .A2(new_n290), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n298), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n911), .A2(new_n912), .A3(new_n1017), .A4(new_n1011), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1011), .B1(new_n996), .B2(new_n981), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n267), .A3(new_n1013), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1015), .A2(new_n1018), .A3(new_n1020), .ZN(G57));
endmodule


