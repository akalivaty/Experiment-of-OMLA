//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  AND2_X1   g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208));
  NAND2_X1  g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT72), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n207), .ZN(new_n213));
  NOR2_X1   g012(.A1(G197gat), .A2(G204gat), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n213), .A2(new_n214), .B1(new_n203), .B2(KEYINPUT22), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n203), .A2(new_n204), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT72), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G162gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G148gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G141gat), .ZN(new_n226));
  INV_X1    g025(.A(G141gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G148gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n229), .B1(new_n226), .B2(new_n228), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n224), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n226), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT78), .B(G141gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT2), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n221), .A3(new_n223), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n237), .A2(KEYINPUT80), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT78), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT78), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G141gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n245), .A3(G148gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n226), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n239), .A2(new_n221), .A3(new_n223), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n242), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n219), .B(new_n234), .C1(new_n241), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT29), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n218), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT80), .B1(new_n237), .B2(new_n240), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(new_n242), .A3(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n226), .A2(new_n228), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT77), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(new_n231), .A3(new_n230), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n253), .A2(new_n254), .B1(new_n224), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT29), .B1(new_n215), .B2(new_n216), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n210), .A2(new_n205), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT3), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n202), .B1(new_n252), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G22gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n234), .B1(new_n241), .B2(new_n249), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n212), .A2(new_n251), .A3(new_n217), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n219), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n202), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT29), .B1(new_n258), .B2(new_n219), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(new_n218), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n263), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT85), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n263), .A2(new_n270), .A3(new_n273), .A4(new_n264), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(new_n270), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G22gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G78gat), .B(G106gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT31), .B(G50gat), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n278), .B(new_n279), .Z(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT86), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT86), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n280), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n286), .A3(new_n271), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT87), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT87), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n276), .A2(new_n289), .A3(new_n286), .A4(new_n271), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT88), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n277), .A2(new_n283), .A3(new_n280), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n283), .B1(new_n277), .B2(new_n280), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT88), .B(new_n291), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT89), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n301), .B2(KEYINPUT23), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n307), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n307), .A2(G169gat), .A3(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT64), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n304), .A2(new_n309), .A3(new_n311), .A4(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n310), .A2(new_n300), .A3(new_n318), .ZN(new_n320));
  INV_X1    g119(.A(G183gat), .ZN(new_n321));
  INV_X1    g120(.A(G190gat), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n315), .A2(KEYINPUT67), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(KEYINPUT67), .B2(new_n315), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT66), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n326), .A2(KEYINPUT24), .A3(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n309), .B(new_n320), .C1(new_n324), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n298), .B2(new_n299), .ZN(new_n332));
  NOR3_X1   g131(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n313), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT68), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(new_n313), .C1(new_n332), .C2(new_n333), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT27), .B(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(new_n322), .ZN(new_n340));
  INV_X1    g139(.A(new_n338), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT28), .B1(new_n341), .B2(G190gat), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n335), .A2(new_n337), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n330), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n345), .B(KEYINPUT73), .Z(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT29), .B1(new_n330), .B2(new_n343), .ZN(new_n348));
  INV_X1    g147(.A(new_n345), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n347), .B(new_n218), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(G8gat), .B(G36gat), .Z(new_n351));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n324), .A2(new_n328), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n320), .A2(new_n309), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n354), .A2(new_n355), .B1(new_n317), .B2(new_n318), .ZN(new_n356));
  AND4_X1   g155(.A1(new_n335), .A2(new_n337), .A3(new_n340), .A4(new_n342), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n251), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n346), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(new_n344), .B2(new_n349), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n350), .B(new_n353), .C1(new_n360), .C2(new_n218), .ZN(new_n361));
  XOR2_X1   g160(.A(KEYINPUT76), .B(KEYINPUT30), .Z(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n350), .B1(new_n360), .B2(new_n218), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n353), .B(KEYINPUT74), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n369));
  OR3_X1    g168(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n361), .B2(new_n369), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(G120gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G113gat), .ZN(new_n376));
  INV_X1    g175(.A(G113gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G120gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n379), .B(new_n380), .C1(new_n381), .C2(KEYINPUT69), .ZN(new_n382));
  INV_X1    g181(.A(G127gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G134gat), .ZN(new_n384));
  INV_X1    g183(.A(G134gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G127gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n380), .A2(KEYINPUT69), .ZN(new_n388));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n387), .B(new_n388), .C1(new_n389), .C2(KEYINPUT1), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n382), .A2(new_n390), .A3(KEYINPUT81), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT81), .B1(new_n382), .B2(new_n390), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n265), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n382), .A2(new_n390), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n395), .B(new_n234), .C1(new_n241), .C2(new_n249), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n374), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n373), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(KEYINPUT4), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n258), .A2(new_n401), .A3(new_n395), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n250), .A3(new_n393), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n404), .A2(new_n374), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n382), .A2(new_n390), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n382), .A2(new_n390), .A3(KEYINPUT81), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n396), .B1(new_n413), .B2(new_n258), .ZN(new_n414));
  INV_X1    g213(.A(new_n374), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n408), .A3(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G1gat), .B(G29gat), .Z(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n400), .A2(new_n402), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n425), .A2(new_n406), .A3(new_n398), .A4(new_n374), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n418), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n424), .B1(new_n418), .B2(new_n426), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT6), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n430), .B(new_n424), .C1(new_n418), .C2(new_n426), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n372), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n295), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n297), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n344), .A2(new_n409), .ZN(new_n440));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n330), .A2(new_n395), .A3(new_n343), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT34), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n440), .A2(new_n445), .A3(new_n441), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(G15gat), .B(G43gat), .Z(new_n449));
  XNOR2_X1  g248(.A(G71gat), .B(G99gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(KEYINPUT33), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n453), .A2(new_n455), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT70), .B(new_n448), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n453), .A2(new_n455), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n447), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n444), .A2(KEYINPUT70), .A3(new_n446), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n456), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n439), .B1(new_n465), .B2(KEYINPUT71), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT71), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n459), .A2(new_n464), .A3(new_n467), .A4(KEYINPUT36), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n365), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n218), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n360), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(new_n218), .ZN(new_n475));
  OAI221_X1 g274(.A(new_n471), .B1(new_n473), .B2(new_n475), .C1(KEYINPUT37), .C2(new_n364), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n361), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n364), .A2(KEYINPUT37), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n364), .A2(KEYINPUT37), .ZN(new_n479));
  OR3_X1    g278(.A1(new_n478), .A2(new_n479), .A3(new_n353), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(KEYINPUT38), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n429), .A2(new_n431), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n374), .B1(new_n425), .B2(new_n406), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT39), .B1(new_n414), .B2(new_n415), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT39), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n424), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT40), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n490), .A2(new_n491), .A3(new_n428), .ZN(new_n492));
  INV_X1    g291(.A(new_n372), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n481), .A2(new_n482), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n435), .A2(new_n295), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n469), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n438), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n432), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n459), .A2(new_n464), .A3(KEYINPUT90), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT90), .B1(new_n459), .B2(new_n464), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n502));
  NAND4_X1  g301(.A1(new_n495), .A2(new_n498), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n465), .ZN(new_n504));
  AOI211_X1 g303(.A(new_n504), .B(new_n432), .C1(new_n435), .C2(new_n295), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT35), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n497), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509));
  INV_X1    g308(.A(G85gat), .ZN(new_n510));
  INV_X1    g309(.A(G92gat), .ZN(new_n511));
  AOI22_X1  g310(.A1(KEYINPUT8), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT102), .ZN(new_n513));
  XOR2_X1   g312(.A(G99gat), .B(G106gat), .Z(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(KEYINPUT103), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OR3_X1    g315(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT7), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT7), .B1(new_n510), .B2(new_n511), .ZN(new_n518));
  AOI22_X1  g317(.A1(KEYINPUT103), .A2(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n513), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n516), .B1(new_n513), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT92), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT14), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n526), .B(new_n529), .C1(G29gat), .C2(G36gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n523), .B2(new_n524), .ZN(new_n532));
  NAND3_X1  g331(.A1(KEYINPUT93), .A2(G29gat), .A3(G36gat), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(new_n530), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(G43gat), .A2(G50gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g335(.A1(G43gat), .A2(G50gat), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n535), .A2(KEYINPUT94), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n534), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT14), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n532), .A2(new_n530), .A3(new_n533), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(new_n540), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT96), .B1(new_n549), .B2(KEYINPUT17), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT96), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  NOR4_X1   g351(.A1(new_n544), .A2(new_n548), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  OAI221_X1 g352(.A(new_n522), .B1(KEYINPUT17), .B2(new_n549), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n522), .A2(new_n549), .ZN(new_n555));
  AND2_X1   g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(KEYINPUT41), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G190gat), .B(G218gat), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n556), .A2(KEYINPUT41), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n559), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n560), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n563), .B1(new_n560), .B2(new_n565), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G71gat), .B(G78gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT99), .B(KEYINPUT21), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G8gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G15gat), .B(G22gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(G1gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n581), .B2(KEYINPUT95), .ZN(new_n582));
  INV_X1    g381(.A(G1gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT16), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(G1gat), .B2(new_n580), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n582), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n574), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(KEYINPUT21), .B2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n578), .B(new_n589), .Z(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT101), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT100), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n590), .B(new_n597), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n569), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT13), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n582), .B(new_n586), .Z(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n549), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n534), .A2(KEYINPUT15), .A3(new_n539), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n543), .A2(new_n538), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n605), .B2(new_n534), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n587), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n601), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n587), .B1(new_n552), .B2(new_n606), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n609), .B1(new_n550), .B2(new_n553), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(new_n600), .A3(new_n607), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n600), .A4(new_n607), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n551), .B1(new_n606), .B2(new_n552), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n549), .A2(KEYINPUT96), .A3(KEYINPUT17), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n619), .A2(new_n609), .B1(new_n587), .B2(new_n606), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n620), .A2(KEYINPUT97), .A3(KEYINPUT18), .A4(new_n600), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n613), .A2(new_n616), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G113gat), .B(G141gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G197gat), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT11), .B(G169gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629));
  INV_X1    g428(.A(new_n627), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n613), .A2(new_n621), .A3(new_n616), .A4(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n622), .A2(KEYINPUT98), .A3(new_n627), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT105), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n588), .B1(new_n520), .B2(new_n521), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n513), .A2(new_n519), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n515), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n513), .A2(new_n519), .A3(new_n516), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n574), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(KEYINPUT10), .B(new_n588), .C1(new_n520), .C2(new_n521), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n639), .B1(new_n641), .B2(new_n645), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n638), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(new_n648), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n647), .A2(KEYINPUT104), .A3(new_n648), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n657), .A3(new_n639), .ZN(new_n658));
  INV_X1    g457(.A(new_n637), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n599), .A2(new_n634), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n508), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n482), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n583), .ZN(G1324gat));
  INV_X1    g466(.A(new_n664), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n579), .B1(new_n668), .B2(new_n493), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n664), .A2(new_n372), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(KEYINPUT42), .B2(new_n671), .ZN(G1325gat));
  INV_X1    g472(.A(new_n501), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n664), .A2(G15gat), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n469), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n664), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n297), .A2(new_n437), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  NOR3_X1   g481(.A1(new_n634), .A2(new_n598), .A3(new_n662), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n508), .A2(new_n568), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n523), .A3(new_n482), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n495), .A2(new_n498), .A3(new_n465), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT35), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n689), .A2(new_n503), .B1(new_n438), .B2(new_n496), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n690), .B2(new_n569), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n508), .A2(KEYINPUT44), .A3(new_n568), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n683), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n665), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n686), .A2(new_n695), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n684), .A2(new_n524), .A3(new_n493), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT46), .Z(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n694), .B2(new_n372), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1329gat));
  NAND4_X1  g499(.A1(new_n691), .A2(new_n692), .A3(new_n469), .A4(new_n683), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G43gat), .ZN(new_n702));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n684), .A2(new_n703), .A3(new_n501), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT47), .B1(new_n705), .B2(KEYINPUT107), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  AOI211_X1 g507(.A(new_n707), .B(new_n708), .C1(new_n702), .C2(new_n704), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n706), .A2(new_n709), .ZN(G1330gat));
  INV_X1    g509(.A(new_n495), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n691), .A2(new_n692), .A3(new_n711), .A4(new_n683), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n679), .A2(G50gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n684), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(KEYINPUT48), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n679), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n693), .A2(new_n717), .A3(new_n683), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n718), .A2(G50gat), .B1(new_n684), .B2(new_n714), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g519(.A(new_n634), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n690), .A2(new_n721), .A3(new_n599), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n662), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n482), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g525(.A(new_n372), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n722), .A2(new_n662), .A3(new_n727), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(G1333gat));
  OAI21_X1  g533(.A(G71gat), .B1(new_n723), .B2(new_n676), .ZN(new_n735));
  INV_X1    g534(.A(G71gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n662), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n674), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n717), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g543(.A1(new_n721), .A2(new_n598), .A3(new_n737), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n693), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n665), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n721), .A2(new_n598), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n508), .A2(new_n568), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n508), .A2(KEYINPUT51), .A3(new_n568), .A4(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n482), .A2(new_n510), .A3(new_n662), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n747), .B1(new_n754), .B2(new_n755), .ZN(G1336gat));
  NOR3_X1   g555(.A1(new_n737), .A2(G92gat), .A3(new_n372), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n691), .A2(new_n692), .A3(new_n493), .A4(new_n745), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n759), .A2(new_n760), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n753), .A2(new_n757), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n759), .A2(G92gat), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT52), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n746), .B2(new_n676), .ZN(new_n769));
  OR3_X1    g568(.A1(new_n674), .A2(G99gat), .A3(new_n737), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n754), .B2(new_n770), .ZN(G1338gat));
  NAND4_X1  g570(.A1(new_n691), .A2(new_n692), .A3(new_n717), .A4(new_n745), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G106gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n495), .A2(G106gat), .A3(new_n737), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n751), .B2(new_n752), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI211_X1 g577(.A(KEYINPUT111), .B(new_n775), .C1(new_n751), .C2(new_n752), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT53), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n776), .A2(KEYINPUT53), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n691), .A2(new_n692), .A3(new_n711), .A4(new_n745), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT112), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n782), .A2(KEYINPUT112), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n780), .A2(new_n786), .ZN(G1339gat));
  NAND4_X1  g586(.A1(new_n634), .A2(new_n598), .A3(new_n569), .A4(new_n737), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n603), .A2(new_n607), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n601), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n792), .A3(new_n601), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n620), .A2(new_n600), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n626), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT114), .B(new_n626), .C1(new_n794), .C2(new_n795), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n631), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n647), .A2(new_n648), .A3(new_n640), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n640), .B1(new_n654), .B2(new_n655), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n657), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n649), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n659), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n801), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n803), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n658), .A2(new_n810), .ZN(new_n811));
  AOI211_X1 g610(.A(new_n801), .B(new_n637), .C1(new_n649), .C2(new_n806), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n809), .A2(new_n661), .A3(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n800), .A2(new_n569), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n662), .A2(new_n798), .A3(new_n631), .A4(new_n799), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n634), .B2(new_n814), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n817), .B2(new_n569), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n788), .B1(new_n818), .B2(new_n598), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n482), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n495), .A2(new_n465), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n493), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n721), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n819), .A2(new_n679), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n482), .A2(new_n372), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n501), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n377), .A3(new_n634), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n826), .A2(new_n831), .ZN(G1340gat));
  OAI21_X1  g631(.A(new_n375), .B1(new_n824), .B2(new_n737), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(G120gat), .A3(new_n738), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT115), .ZN(G1341gat));
  NAND3_X1  g635(.A1(new_n825), .A2(new_n383), .A3(new_n598), .ZN(new_n837));
  INV_X1    g636(.A(new_n598), .ZN(new_n838));
  OAI21_X1  g637(.A(G127gat), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(G1342gat));
  NAND4_X1  g639(.A1(new_n821), .A2(new_n385), .A3(new_n568), .A4(new_n823), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n842));
  OAI21_X1  g641(.A(G134gat), .B1(new_n830), .B2(new_n569), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT116), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n842), .A2(new_n843), .A3(new_n847), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1343gat));
  XNOR2_X1  g648(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n808), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n811), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n659), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n661), .B1(new_n805), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT117), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n809), .A2(new_n813), .A3(new_n857), .A4(new_n661), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n856), .A2(new_n632), .A3(new_n633), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n568), .B1(new_n859), .B2(new_n816), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n838), .B1(new_n860), .B2(new_n815), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n788), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n717), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n469), .A2(new_n828), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n819), .A2(new_n711), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n679), .B1(new_n861), .B2(new_n788), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT118), .B1(new_n869), .B2(KEYINPUT57), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n865), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n236), .B1(new_n871), .B2(new_n721), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n820), .A2(KEYINPUT119), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n820), .A2(KEYINPUT119), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n469), .A2(new_n495), .A3(new_n493), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n721), .A2(new_n227), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n851), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n236), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n870), .A2(new_n868), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n863), .A3(new_n864), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n882), .B2(new_n634), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n876), .A2(new_n877), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n884), .A3(new_n850), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n879), .A2(new_n885), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n737), .A2(G148gat), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n866), .A2(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n869), .A2(new_n867), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n737), .B1(new_n864), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT122), .B1(new_n469), .B2(new_n828), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n892), .A2(new_n893), .A3(new_n894), .A4(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(G148gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n892), .A2(new_n893), .A3(new_n898), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT123), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n891), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n891), .A2(G148gat), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n904), .B1(new_n871), .B2(new_n662), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n890), .B1(new_n903), .B2(new_n905), .ZN(G1345gat));
  NOR2_X1   g705(.A1(new_n882), .A2(new_n838), .ZN(new_n907));
  XOR2_X1   g706(.A(KEYINPUT79), .B(G155gat), .Z(new_n908));
  NAND2_X1  g707(.A1(new_n598), .A2(new_n908), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n907), .A2(new_n908), .B1(new_n876), .B2(new_n909), .ZN(G1346gat));
  OR2_X1    g709(.A1(new_n876), .A2(new_n569), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n569), .A2(new_n220), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n911), .A2(new_n220), .B1(new_n871), .B2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n482), .A2(new_n372), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n819), .A2(new_n679), .A3(new_n501), .A4(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(new_n298), .A3(new_n634), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n819), .A2(new_n665), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(new_n372), .A3(new_n822), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n721), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n919), .B2(new_n298), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT124), .Z(G1348gat));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n299), .A3(new_n662), .ZN(new_n922));
  OAI21_X1  g721(.A(G176gat), .B1(new_n915), .B2(new_n737), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT125), .ZN(G1349gat));
  NOR2_X1   g724(.A1(new_n838), .A2(new_n341), .ZN(new_n926));
  AOI22_X1  g725(.A1(new_n918), .A2(new_n926), .B1(KEYINPUT126), .B2(KEYINPUT60), .ZN(new_n927));
  OAI21_X1  g726(.A(G183gat), .B1(new_n915), .B2(new_n838), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g728(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n915), .B2(new_n569), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT61), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n322), .A3(new_n568), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1351gat));
  AND2_X1   g734(.A1(new_n892), .A2(new_n893), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n469), .A2(new_n482), .A3(new_n372), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n936), .A2(G197gat), .A3(new_n721), .A4(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G197gat), .ZN(new_n939));
  INV_X1    g738(.A(new_n917), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n676), .A2(new_n711), .A3(new_n493), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT127), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n939), .B1(new_n943), .B2(new_n634), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n938), .A2(new_n944), .ZN(G1352gat));
  NOR3_X1   g744(.A1(new_n943), .A2(G204gat), .A3(new_n737), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT62), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n936), .A2(new_n937), .ZN(new_n948));
  OAI21_X1  g747(.A(G204gat), .B1(new_n948), .B2(new_n737), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1353gat));
  OR3_X1    g749(.A1(new_n943), .A2(G211gat), .A3(new_n838), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n936), .A2(new_n598), .A3(new_n937), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  OAI21_X1  g754(.A(G218gat), .B1(new_n948), .B2(new_n569), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n569), .A2(G218gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n943), .B2(new_n957), .ZN(G1355gat));
endmodule


