

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753;

  XNOR2_X1 U371 ( .A(KEYINPUT76), .B(G110), .ZN(n430) );
  XNOR2_X1 U372 ( .A(n552), .B(KEYINPUT109), .ZN(n399) );
  NOR2_X2 U373 ( .A1(G902), .A2(n707), .ZN(n437) );
  XNOR2_X2 U374 ( .A(n366), .B(n428), .ZN(n739) );
  XNOR2_X2 U375 ( .A(n441), .B(KEYINPUT4), .ZN(n366) );
  NOR2_X2 U376 ( .A1(n750), .A2(n751), .ZN(n553) );
  INV_X1 U377 ( .A(n654), .ZN(n651) );
  XNOR2_X1 U378 ( .A(n495), .B(n494), .ZN(n507) );
  NOR2_X1 U379 ( .A1(n631), .A2(n721), .ZN(n632) );
  BUF_X1 U380 ( .A(n706), .Z(n717) );
  AND2_X1 U381 ( .A1(n574), .A2(n573), .ZN(n744) );
  XNOR2_X1 U382 ( .A(n539), .B(KEYINPUT32), .ZN(n575) );
  NOR2_X1 U383 ( .A1(n687), .A2(n596), .ZN(n597) );
  XNOR2_X1 U384 ( .A(n595), .B(n594), .ZN(n687) );
  NAND2_X1 U385 ( .A1(n399), .A2(n670), .ZN(n419) );
  NAND2_X1 U386 ( .A1(n416), .A2(n668), .ZN(n552) );
  XNOR2_X1 U387 ( .A(n679), .B(KEYINPUT6), .ZN(n591) );
  NAND2_X2 U388 ( .A1(n385), .A2(n386), .ZN(n679) );
  INV_X2 U389 ( .A(n525), .ZN(n546) );
  AND2_X1 U390 ( .A1(n361), .A2(n358), .ZN(n385) );
  XNOR2_X1 U391 ( .A(n507), .B(n506), .ZN(n728) );
  XNOR2_X1 U392 ( .A(n398), .B(G119), .ZN(n495) );
  XOR2_X1 U393 ( .A(G137), .B(G140), .Z(n461) );
  XNOR2_X1 U394 ( .A(G104), .B(G107), .ZN(n429) );
  XNOR2_X1 U395 ( .A(KEYINPUT16), .B(G122), .ZN(n506) );
  INV_X1 U396 ( .A(KEYINPUT73), .ZN(n493) );
  NOR2_X1 U397 ( .A1(n681), .A2(n682), .ZN(n593) );
  XNOR2_X1 U398 ( .A(n410), .B(KEYINPUT103), .ZN(n654) );
  OR2_X1 U399 ( .A1(n551), .A2(n682), .ZN(n598) );
  XNOR2_X2 U400 ( .A(KEYINPUT68), .B(G101), .ZN(n485) );
  XNOR2_X2 U401 ( .A(n727), .B(n485), .ZN(n508) );
  XNOR2_X2 U402 ( .A(n431), .B(n430), .ZN(n727) );
  XNOR2_X2 U403 ( .A(n580), .B(n579), .ZN(n666) );
  AND2_X1 U404 ( .A1(n647), .A2(n356), .ZN(n412) );
  INV_X1 U405 ( .A(KEYINPUT69), .ZN(n413) );
  INV_X1 U406 ( .A(G237), .ZN(n500) );
  XNOR2_X1 U407 ( .A(n401), .B(G125), .ZN(n512) );
  INV_X1 U408 ( .A(G146), .ZN(n401) );
  NAND2_X1 U409 ( .A1(n675), .A2(n676), .ZN(n682) );
  OR2_X1 U410 ( .A1(n633), .A2(n387), .ZN(n386) );
  NAND2_X1 U411 ( .A1(n388), .A2(n501), .ZN(n387) );
  INV_X1 U412 ( .A(G472), .ZN(n388) );
  XNOR2_X1 U413 ( .A(n562), .B(KEYINPUT104), .ZN(n667) );
  XNOR2_X1 U414 ( .A(n571), .B(KEYINPUT48), .ZN(n574) );
  AND2_X1 U415 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U416 ( .A1(n373), .A2(n372), .ZN(n371) );
  INV_X1 U417 ( .A(KEYINPUT2), .ZN(n372) );
  NOR2_X1 U418 ( .A1(n523), .A2(n369), .ZN(n368) );
  INV_X1 U419 ( .A(n416), .ZN(n369) );
  OR2_X1 U420 ( .A1(n499), .A2(n591), .ZN(n554) );
  XNOR2_X1 U421 ( .A(G128), .B(G119), .ZN(n462) );
  XNOR2_X1 U422 ( .A(G110), .B(KEYINPUT93), .ZN(n466) );
  XOR2_X1 U423 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n467) );
  XOR2_X1 U424 ( .A(G122), .B(G104), .Z(n452) );
  XNOR2_X1 U425 ( .A(G113), .B(G140), .ZN(n451) );
  XNOR2_X1 U426 ( .A(n407), .B(KEYINPUT11), .ZN(n406) );
  NAND2_X1 U427 ( .A1(n486), .A2(G214), .ZN(n407) );
  XNOR2_X1 U428 ( .A(n454), .B(n409), .ZN(n408) );
  XNOR2_X1 U429 ( .A(KEYINPUT12), .B(KEYINPUT98), .ZN(n409) );
  XNOR2_X1 U430 ( .A(n512), .B(n400), .ZN(n735) );
  INV_X1 U431 ( .A(KEYINPUT10), .ZN(n400) );
  XNOR2_X1 U432 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n510) );
  NAND2_X1 U433 ( .A1(n628), .A2(n609), .ZN(n389) );
  AND2_X1 U434 ( .A1(n415), .A2(n414), .ZN(n647) );
  INV_X1 U435 ( .A(n551), .ZN(n414) );
  XNOR2_X1 U436 ( .A(n411), .B(n459), .ZN(n560) );
  OR2_X1 U437 ( .A1(n620), .A2(G902), .ZN(n411) );
  XNOR2_X1 U438 ( .A(n472), .B(n403), .ZN(n402) );
  OR2_X1 U439 ( .A1(n718), .A2(G902), .ZN(n404) );
  INV_X1 U440 ( .A(KEYINPUT25), .ZN(n403) );
  NOR2_X1 U441 ( .A1(n660), .A2(n567), .ZN(n568) );
  AND2_X1 U442 ( .A1(n412), .A2(n667), .ZN(n564) );
  NAND2_X1 U443 ( .A1(n384), .A2(n668), .ZN(n383) );
  XOR2_X1 U444 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n490) );
  NOR2_X1 U445 ( .A1(G953), .A2(G237), .ZN(n486) );
  NOR2_X1 U446 ( .A1(n359), .A2(n350), .ZN(n394) );
  NOR2_X1 U447 ( .A1(n385), .A2(n383), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n555), .B(n528), .ZN(n563) );
  XOR2_X1 U449 ( .A(G122), .B(G107), .Z(n439) );
  XNOR2_X1 U450 ( .A(G134), .B(G116), .ZN(n438) );
  XNOR2_X1 U451 ( .A(KEYINPUT7), .B(KEYINPUT101), .ZN(n444) );
  XOR2_X1 U452 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n445) );
  AND2_X1 U453 ( .A1(n722), .A2(n374), .ZN(n665) );
  XNOR2_X1 U454 ( .A(n376), .B(n375), .ZN(n374) );
  INV_X1 U455 ( .A(KEYINPUT86), .ZN(n375) );
  INV_X1 U456 ( .A(n554), .ZN(n502) );
  XNOR2_X1 U457 ( .A(n370), .B(n426), .ZN(n397) );
  INV_X1 U458 ( .A(KEYINPUT97), .ZN(n594) );
  XNOR2_X1 U459 ( .A(n471), .B(n470), .ZN(n718) );
  XNOR2_X1 U460 ( .A(n408), .B(n406), .ZN(n455) );
  XNOR2_X1 U461 ( .A(n421), .B(n420), .ZN(n628) );
  XNOR2_X1 U462 ( .A(n728), .B(n422), .ZN(n421) );
  AND2_X1 U463 ( .A1(n623), .A2(G953), .ZN(n721) );
  XNOR2_X1 U464 ( .A(n418), .B(n417), .ZN(n750) );
  INV_X1 U465 ( .A(KEYINPUT42), .ZN(n417) );
  XNOR2_X1 U466 ( .A(n548), .B(KEYINPUT40), .ZN(n751) );
  AND2_X1 U467 ( .A1(n397), .A2(n651), .ZN(n548) );
  NOR2_X1 U468 ( .A1(n561), .A2(n560), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n395), .B(KEYINPUT22), .ZN(n541) );
  AND2_X1 U470 ( .A1(n424), .A2(KEYINPUT85), .ZN(n350) );
  OR2_X1 U471 ( .A1(n524), .A2(n523), .ZN(n351) );
  AND2_X1 U472 ( .A1(n664), .A2(n663), .ZN(n352) );
  XOR2_X1 U473 ( .A(n516), .B(n515), .Z(n353) );
  AND2_X1 U474 ( .A1(n386), .A2(n520), .ZN(n354) );
  NOR2_X1 U475 ( .A1(n416), .A2(n668), .ZN(n355) );
  AND2_X1 U476 ( .A1(n646), .A2(n413), .ZN(n356) );
  AND2_X1 U477 ( .A1(n540), .A2(n681), .ZN(n357) );
  NAND2_X1 U478 ( .A1(G902), .A2(G472), .ZN(n358) );
  NOR2_X1 U479 ( .A1(n614), .A2(n613), .ZN(n359) );
  INV_X1 U480 ( .A(n611), .ZN(n424) );
  AND2_X1 U481 ( .A1(n391), .A2(n615), .ZN(n360) );
  NAND2_X1 U482 ( .A1(n525), .A2(n668), .ZN(n555) );
  XNOR2_X2 U483 ( .A(n389), .B(n353), .ZN(n525) );
  NAND2_X1 U484 ( .A1(n633), .A2(G472), .ZN(n361) );
  INV_X1 U485 ( .A(n598), .ZN(n518) );
  XNOR2_X1 U486 ( .A(n550), .B(KEYINPUT28), .ZN(n415) );
  NAND2_X1 U487 ( .A1(n362), .A2(n589), .ZN(n607) );
  NAND2_X1 U488 ( .A1(n587), .A2(n588), .ZN(n362) );
  NAND2_X1 U489 ( .A1(n405), .A2(n394), .ZN(n393) );
  NAND2_X1 U490 ( .A1(n363), .A2(n357), .ZN(n543) );
  INV_X1 U491 ( .A(n541), .ZN(n363) );
  AND2_X1 U492 ( .A1(n392), .A2(n360), .ZN(n390) );
  XNOR2_X1 U493 ( .A(n364), .B(n605), .ZN(n606) );
  NAND2_X1 U494 ( .A1(n603), .A2(n604), .ZN(n364) );
  NAND2_X1 U495 ( .A1(n365), .A2(n667), .ZN(n601) );
  NAND2_X1 U496 ( .A1(n656), .A2(n642), .ZN(n365) );
  NAND2_X1 U497 ( .A1(n393), .A2(n390), .ZN(n617) );
  NAND2_X1 U498 ( .A1(n593), .A2(n679), .ZN(n595) );
  XNOR2_X1 U499 ( .A(n366), .B(n508), .ZN(n420) );
  NAND2_X1 U500 ( .A1(n368), .A2(n367), .ZN(n370) );
  INV_X1 U501 ( .A(n524), .ZN(n367) );
  NAND2_X1 U502 ( .A1(n574), .A2(n371), .ZN(n376) );
  INV_X1 U503 ( .A(n573), .ZN(n373) );
  NAND2_X1 U504 ( .A1(n378), .A2(n377), .ZN(n522) );
  NAND2_X1 U505 ( .A1(n385), .A2(n354), .ZN(n377) );
  NOR2_X1 U506 ( .A1(n382), .A2(n379), .ZN(n378) );
  NAND2_X1 U507 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U508 ( .A1(n527), .A2(n520), .ZN(n380) );
  OR2_X1 U509 ( .A1(n386), .A2(n383), .ZN(n381) );
  INV_X1 U510 ( .A(n520), .ZN(n384) );
  NAND2_X1 U511 ( .A1(n394), .A2(n611), .ZN(n391) );
  NAND2_X1 U512 ( .A1(n664), .A2(KEYINPUT85), .ZN(n392) );
  NAND2_X1 U513 ( .A1(n600), .A2(n535), .ZN(n395) );
  XNOR2_X2 U514 ( .A(n532), .B(n425), .ZN(n600) );
  INV_X1 U515 ( .A(n396), .ZN(n587) );
  NAND2_X1 U516 ( .A1(n576), .A2(n575), .ZN(n396) );
  NAND2_X1 U517 ( .A1(n545), .A2(n544), .ZN(n576) );
  NAND2_X1 U518 ( .A1(n396), .A2(n577), .ZN(n589) );
  NAND2_X1 U519 ( .A1(n397), .A2(n648), .ZN(n662) );
  XNOR2_X2 U520 ( .A(G116), .B(KEYINPUT3), .ZN(n398) );
  NAND2_X1 U521 ( .A1(n399), .A2(n667), .ZN(n673) );
  XNOR2_X2 U522 ( .A(n404), .B(n402), .ZN(n675) );
  INV_X1 U523 ( .A(n664), .ZN(n405) );
  XNOR2_X2 U524 ( .A(n546), .B(KEYINPUT38), .ZN(n416) );
  NAND2_X1 U525 ( .A1(n691), .A2(n647), .ZN(n418) );
  XNOR2_X2 U526 ( .A(n419), .B(KEYINPUT41), .ZN(n691) );
  XNOR2_X1 U527 ( .A(n511), .B(n423), .ZN(n422) );
  XNOR2_X1 U528 ( .A(n512), .B(n510), .ZN(n423) );
  XNOR2_X1 U529 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U530 ( .A1(n744), .A2(n722), .ZN(n664) );
  XNOR2_X2 U531 ( .A(n551), .B(KEYINPUT1), .ZN(n681) );
  XNOR2_X2 U532 ( .A(n437), .B(n436), .ZN(n551) );
  XOR2_X1 U533 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n425) );
  XOR2_X1 U534 ( .A(n547), .B(KEYINPUT39), .Z(n426) );
  INV_X1 U535 ( .A(KEYINPUT30), .ZN(n519) );
  XNOR2_X1 U536 ( .A(n519), .B(KEYINPUT108), .ZN(n520) );
  INV_X1 U537 ( .A(KEYINPUT88), .ZN(n605) );
  XNOR2_X1 U538 ( .A(n554), .B(KEYINPUT110), .ZN(n556) );
  XNOR2_X1 U539 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U540 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n557) );
  XNOR2_X2 U541 ( .A(G128), .B(KEYINPUT79), .ZN(n427) );
  XNOR2_X2 U542 ( .A(n427), .B(G143), .ZN(n441) );
  XNOR2_X1 U543 ( .A(G131), .B(G134), .ZN(n428) );
  XNOR2_X2 U544 ( .A(n739), .B(G146), .ZN(n498) );
  XOR2_X1 U545 ( .A(KEYINPUT92), .B(n461), .Z(n736) );
  INV_X1 U546 ( .A(n736), .ZN(n432) );
  INV_X1 U547 ( .A(n429), .ZN(n431) );
  XNOR2_X1 U548 ( .A(n432), .B(n508), .ZN(n434) );
  INV_X2 U549 ( .A(G953), .ZN(n746) );
  NAND2_X1 U550 ( .A1(G227), .A2(n746), .ZN(n433) );
  XNOR2_X1 U551 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U552 ( .A(n435), .B(n498), .ZN(n707) );
  XNOR2_X1 U553 ( .A(KEYINPUT72), .B(G469), .ZN(n436) );
  INV_X1 U554 ( .A(n681), .ZN(n504) );
  XNOR2_X1 U555 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U556 ( .A(n441), .B(n440), .ZN(n449) );
  NAND2_X1 U557 ( .A1(G234), .A2(n746), .ZN(n443) );
  XOR2_X1 U558 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n442) );
  XNOR2_X1 U559 ( .A(n443), .B(n442), .ZN(n465) );
  NAND2_X1 U560 ( .A1(G217), .A2(n465), .ZN(n447) );
  XNOR2_X1 U561 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U562 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U563 ( .A(n449), .B(n448), .ZN(n713) );
  NOR2_X1 U564 ( .A1(G902), .A2(n713), .ZN(n450) );
  XNOR2_X1 U565 ( .A(G478), .B(n450), .ZN(n533) );
  INV_X1 U566 ( .A(n533), .ZN(n561) );
  XNOR2_X1 U567 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U568 ( .A(n735), .B(n453), .ZN(n456) );
  XNOR2_X1 U569 ( .A(G143), .B(G131), .ZN(n454) );
  XNOR2_X1 U570 ( .A(n456), .B(n455), .ZN(n620) );
  XOR2_X1 U571 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n458) );
  XNOR2_X1 U572 ( .A(KEYINPUT13), .B(G475), .ZN(n457) );
  XNOR2_X1 U573 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U574 ( .A(G902), .B(KEYINPUT15), .ZN(n609) );
  NAND2_X1 U575 ( .A1(n609), .A2(G234), .ZN(n460) );
  XNOR2_X1 U576 ( .A(n460), .B(KEYINPUT20), .ZN(n473) );
  NAND2_X1 U577 ( .A1(n473), .A2(G217), .ZN(n472) );
  INV_X1 U578 ( .A(n461), .ZN(n463) );
  XNOR2_X1 U579 ( .A(n735), .B(n464), .ZN(n471) );
  NAND2_X1 U580 ( .A1(G221), .A2(n465), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U582 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U583 ( .A1(n473), .A2(G221), .ZN(n475) );
  XOR2_X1 U584 ( .A(KEYINPUT94), .B(KEYINPUT21), .Z(n474) );
  XNOR2_X1 U585 ( .A(n475), .B(n474), .ZN(n676) );
  NAND2_X1 U586 ( .A1(G234), .A2(G237), .ZN(n476) );
  XNOR2_X1 U587 ( .A(n476), .B(KEYINPUT14), .ZN(n696) );
  NOR2_X1 U588 ( .A1(G902), .A2(n746), .ZN(n478) );
  NOR2_X1 U589 ( .A1(G953), .A2(G952), .ZN(n477) );
  NOR2_X1 U590 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U591 ( .A1(n696), .A2(n479), .ZN(n530) );
  INV_X1 U592 ( .A(n530), .ZN(n481) );
  NAND2_X1 U593 ( .A1(G953), .A2(G900), .ZN(n480) );
  NAND2_X1 U594 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U595 ( .A(KEYINPUT81), .B(n482), .ZN(n521) );
  NAND2_X1 U596 ( .A1(n676), .A2(n521), .ZN(n483) );
  XOR2_X1 U597 ( .A(KEYINPUT71), .B(n483), .Z(n484) );
  NOR2_X1 U598 ( .A1(n675), .A2(n484), .ZN(n549) );
  NAND2_X1 U599 ( .A1(n651), .A2(n549), .ZN(n499) );
  XNOR2_X1 U600 ( .A(n485), .B(KEYINPUT75), .ZN(n488) );
  NAND2_X1 U601 ( .A1(n486), .A2(G210), .ZN(n487) );
  XNOR2_X1 U602 ( .A(n488), .B(n487), .ZN(n492) );
  XNOR2_X1 U603 ( .A(G137), .B(KEYINPUT95), .ZN(n489) );
  XNOR2_X1 U604 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U605 ( .A(n492), .B(n491), .ZN(n496) );
  XNOR2_X1 U606 ( .A(n493), .B(G113), .ZN(n494) );
  XNOR2_X1 U607 ( .A(n507), .B(n496), .ZN(n497) );
  XNOR2_X1 U608 ( .A(n498), .B(n497), .ZN(n633) );
  INV_X1 U609 ( .A(G902), .ZN(n501) );
  NAND2_X1 U610 ( .A1(n501), .A2(n500), .ZN(n513) );
  NAND2_X1 U611 ( .A1(n513), .A2(G214), .ZN(n668) );
  NAND2_X1 U612 ( .A1(n502), .A2(n668), .ZN(n503) );
  NOR2_X1 U613 ( .A1(n504), .A2(n503), .ZN(n505) );
  XOR2_X1 U614 ( .A(n505), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U615 ( .A1(n746), .A2(G224), .ZN(n509) );
  XNOR2_X1 U616 ( .A(n509), .B(KEYINPUT90), .ZN(n511) );
  NAND2_X1 U617 ( .A1(n513), .A2(G210), .ZN(n516) );
  INV_X1 U618 ( .A(KEYINPUT80), .ZN(n514) );
  XNOR2_X1 U619 ( .A(n514), .B(KEYINPUT91), .ZN(n515) );
  NAND2_X1 U620 ( .A1(n517), .A2(n546), .ZN(n572) );
  XNOR2_X1 U621 ( .A(n572), .B(G140), .ZN(G42) );
  OR2_X1 U622 ( .A1(n533), .A2(n560), .ZN(n583) );
  XNOR2_X1 U623 ( .A(n518), .B(KEYINPUT107), .ZN(n524) );
  NAND2_X1 U624 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U625 ( .A1(n583), .A2(n351), .ZN(n526) );
  NAND2_X1 U626 ( .A1(n526), .A2(n525), .ZN(n565) );
  XNOR2_X1 U627 ( .A(n565), .B(G143), .ZN(G45) );
  INV_X1 U628 ( .A(n668), .ZN(n527) );
  INV_X1 U629 ( .A(KEYINPUT19), .ZN(n528) );
  AND2_X1 U630 ( .A1(G953), .A2(G898), .ZN(n529) );
  OR2_X1 U631 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X2 U632 ( .A1(n563), .A2(n531), .ZN(n532) );
  NAND2_X1 U633 ( .A1(n533), .A2(n560), .ZN(n534) );
  XNOR2_X1 U634 ( .A(n534), .B(KEYINPUT105), .ZN(n670) );
  AND2_X1 U635 ( .A1(n670), .A2(n676), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n591), .B(KEYINPUT78), .ZN(n537) );
  NOR2_X1 U637 ( .A1(n681), .A2(n675), .ZN(n536) );
  NAND2_X1 U638 ( .A1(n537), .A2(n536), .ZN(n538) );
  OR2_X1 U639 ( .A1(n541), .A2(n538), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n575), .B(G119), .ZN(G21) );
  INV_X1 U641 ( .A(n679), .ZN(n540) );
  INV_X1 U642 ( .A(KEYINPUT64), .ZN(n542) );
  XNOR2_X1 U643 ( .A(n543), .B(n542), .ZN(n545) );
  INV_X1 U644 ( .A(n675), .ZN(n544) );
  XNOR2_X1 U645 ( .A(n576), .B(G110), .ZN(G12) );
  XNOR2_X1 U646 ( .A(KEYINPUT74), .B(KEYINPUT87), .ZN(n547) );
  AND2_X1 U647 ( .A1(n679), .A2(n549), .ZN(n550) );
  XNOR2_X1 U648 ( .A(n553), .B(KEYINPUT46), .ZN(n570) );
  NOR2_X1 U649 ( .A1(n556), .A2(n555), .ZN(n558) );
  NOR2_X1 U650 ( .A1(n681), .A2(n559), .ZN(n660) );
  NAND2_X1 U651 ( .A1(n561), .A2(n560), .ZN(n657) );
  NAND2_X1 U652 ( .A1(n657), .A2(n654), .ZN(n562) );
  INV_X1 U653 ( .A(n563), .ZN(n646) );
  XNOR2_X1 U654 ( .A(n564), .B(KEYINPUT47), .ZN(n566) );
  NAND2_X1 U655 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U656 ( .A(KEYINPUT70), .B(n568), .ZN(n569) );
  INV_X1 U657 ( .A(n657), .ZN(n648) );
  AND2_X1 U658 ( .A1(n662), .A2(n572), .ZN(n573) );
  INV_X1 U659 ( .A(KEYINPUT44), .ZN(n577) );
  INV_X1 U660 ( .A(n591), .ZN(n578) );
  NAND2_X1 U661 ( .A1(n578), .A2(n593), .ZN(n580) );
  XNOR2_X1 U662 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n579) );
  NAND2_X1 U663 ( .A1(n666), .A2(n600), .ZN(n582) );
  XNOR2_X1 U664 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n581) );
  XNOR2_X1 U665 ( .A(n582), .B(n581), .ZN(n585) );
  INV_X1 U666 ( .A(n583), .ZN(n584) );
  NAND2_X1 U667 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X2 U668 ( .A(n586), .B(KEYINPUT35), .ZN(n752) );
  OR2_X1 U669 ( .A1(n752), .A2(KEYINPUT44), .ZN(n588) );
  NAND2_X1 U670 ( .A1(n752), .A2(KEYINPUT44), .ZN(n604) );
  AND2_X1 U671 ( .A1(n681), .A2(n675), .ZN(n590) );
  AND2_X1 U672 ( .A1(n591), .A2(n590), .ZN(n592) );
  AND2_X1 U673 ( .A1(n363), .A2(n592), .ZN(n639) );
  INV_X1 U674 ( .A(n639), .ZN(n602) );
  INV_X1 U675 ( .A(n600), .ZN(n596) );
  XNOR2_X1 U676 ( .A(n597), .B(KEYINPUT31), .ZN(n656) );
  NOR2_X1 U677 ( .A1(n598), .A2(n679), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n642) );
  AND2_X1 U679 ( .A1(n601), .A2(n602), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X2 U681 ( .A(n608), .B(KEYINPUT45), .ZN(n722) );
  INV_X1 U682 ( .A(n609), .ZN(n614) );
  NAND2_X1 U683 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n614), .A2(n610), .ZN(n611) );
  INV_X1 U685 ( .A(KEYINPUT85), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n612), .A2(KEYINPUT66), .ZN(n613) );
  OR2_X1 U687 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n615) );
  INV_X1 U688 ( .A(n665), .ZN(n616) );
  AND2_X2 U689 ( .A1(n617), .A2(n616), .ZN(n706) );
  AND2_X2 U690 ( .A1(n706), .A2(G475), .ZN(n622) );
  XNOR2_X1 U691 ( .A(KEYINPUT65), .B(KEYINPUT120), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(KEYINPUT59), .ZN(n619) );
  XOR2_X1 U693 ( .A(n620), .B(n619), .Z(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(n624) );
  INV_X1 U695 ( .A(G952), .ZN(n623) );
  NOR2_X2 U696 ( .A1(n624), .A2(n721), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n625), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U698 ( .A1(n706), .A2(G210), .ZN(n630) );
  XNOR2_X1 U699 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(KEYINPUT55), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U704 ( .A(KEYINPUT63), .ZN(n638) );
  NAND2_X1 U705 ( .A1(n706), .A2(G472), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n633), .B(KEYINPUT62), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X2 U708 ( .A1(n636), .A2(n721), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(G57) );
  XOR2_X1 U710 ( .A(G101), .B(n639), .Z(G3) );
  NOR2_X1 U711 ( .A1(n654), .A2(n642), .ZN(n641) );
  XNOR2_X1 U712 ( .A(G104), .B(KEYINPUT111), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(G6) );
  NOR2_X1 U714 ( .A1(n657), .A2(n642), .ZN(n644) );
  XNOR2_X1 U715 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U717 ( .A(G107), .B(n645), .ZN(G9) );
  XOR2_X1 U718 ( .A(G128), .B(KEYINPUT29), .Z(n650) );
  AND2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n652) );
  NAND2_X1 U720 ( .A1(n652), .A2(n648), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(G30) );
  NAND2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n653), .B(G146), .ZN(G48) );
  NOR2_X1 U724 ( .A1(n654), .A2(n656), .ZN(n655) );
  XOR2_X1 U725 ( .A(G113), .B(n655), .Z(G15) );
  NOR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U727 ( .A(KEYINPUT112), .B(n658), .Z(n659) );
  XNOR2_X1 U728 ( .A(G116), .B(n659), .ZN(G18) );
  XNOR2_X1 U729 ( .A(G125), .B(n660), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U731 ( .A(G134), .B(n662), .ZN(G36) );
  XNOR2_X1 U732 ( .A(KEYINPUT83), .B(KEYINPUT2), .ZN(n663) );
  NOR2_X1 U733 ( .A1(n665), .A2(n352), .ZN(n702) );
  NAND2_X1 U734 ( .A1(n691), .A2(n666), .ZN(n700) );
  XOR2_X1 U735 ( .A(KEYINPUT116), .B(n355), .Z(n669) );
  NAND2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U737 ( .A(KEYINPUT117), .B(n671), .Z(n672) );
  NAND2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U739 ( .A1(n674), .A2(n666), .ZN(n694) );
  NOR2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U741 ( .A(KEYINPUT49), .B(n677), .Z(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U743 ( .A(KEYINPUT113), .B(n680), .Z(n686) );
  NAND2_X1 U744 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n683), .B(KEYINPUT50), .ZN(n684) );
  XNOR2_X1 U746 ( .A(KEYINPUT114), .B(n684), .ZN(n685) );
  NAND2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n688) );
  NAND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U749 ( .A(n689), .B(KEYINPUT51), .ZN(n690) );
  XNOR2_X1 U750 ( .A(KEYINPUT115), .B(n690), .ZN(n692) );
  NAND2_X1 U751 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U752 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U753 ( .A(KEYINPUT52), .B(n695), .Z(n698) );
  NAND2_X1 U754 ( .A1(n696), .A2(G952), .ZN(n697) );
  OR2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U756 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U758 ( .A(KEYINPUT118), .B(n703), .Z(n704) );
  NOR2_X1 U759 ( .A1(G953), .A2(n704), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n705), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U761 ( .A1(n717), .A2(G469), .ZN(n711) );
  XNOR2_X1 U762 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n707), .B(KEYINPUT57), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n721), .A2(n712), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n717), .A2(G478), .ZN(n715) );
  XOR2_X1 U768 ( .A(n713), .B(KEYINPUT121), .Z(n714) );
  XNOR2_X1 U769 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U770 ( .A1(n721), .A2(n716), .ZN(G63) );
  NAND2_X1 U771 ( .A1(n717), .A2(G217), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n721), .A2(n720), .ZN(G66) );
  NAND2_X1 U774 ( .A1(n722), .A2(n746), .ZN(n726) );
  NAND2_X1 U775 ( .A1(G953), .A2(G224), .ZN(n723) );
  XNOR2_X1 U776 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U777 ( .A1(n724), .A2(G898), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n726), .A2(n725), .ZN(n734) );
  XOR2_X1 U779 ( .A(n727), .B(KEYINPUT122), .Z(n729) );
  XNOR2_X1 U780 ( .A(n728), .B(n729), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n730), .B(G101), .ZN(n732) );
  NOR2_X1 U782 ( .A1(n746), .A2(G898), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U784 ( .A(n734), .B(n733), .ZN(G69) );
  XOR2_X1 U785 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n738) );
  XNOR2_X1 U786 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n738), .B(n737), .ZN(n740) );
  XOR2_X1 U788 ( .A(n739), .B(n740), .Z(n745) );
  XOR2_X1 U789 ( .A(G227), .B(n745), .Z(n741) );
  NAND2_X1 U790 ( .A1(n741), .A2(G900), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n742), .A2(G953), .ZN(n743) );
  XOR2_X1 U792 ( .A(KEYINPUT125), .B(n743), .Z(n749) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U796 ( .A(G137), .B(n750), .Z(G39) );
  XOR2_X1 U797 ( .A(G131), .B(n751), .Z(G33) );
  XOR2_X1 U798 ( .A(n752), .B(G122), .Z(n753) );
  XNOR2_X1 U799 ( .A(KEYINPUT126), .B(n753), .ZN(G24) );
endmodule

