//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n201), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(G50), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n212), .B1(new_n215), .B2(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n213), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI22_X1  g0053(.A1(new_n250), .A2(new_n252), .B1(new_n207), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT15), .B(G87), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n207), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n249), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT69), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G77), .ZN(new_n261));
  INV_X1    g0061(.A(new_n249), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G1), .B2(new_n207), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n261), .B1(new_n264), .B2(G77), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n271), .B1(G244), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n283), .A2(G238), .B1(G107), .B2(new_n281), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n279), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G232), .A3(new_n282), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n213), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n276), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G200), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n267), .B(new_n294), .C1(new_n295), .C2(new_n293), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n293), .A2(G179), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n266), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT70), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n271), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n275), .A2(G226), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n283), .A2(G223), .B1(G77), .B2(new_n281), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n287), .A2(G222), .A3(new_n282), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n307), .B2(new_n268), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G179), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n251), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT67), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n250), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G58), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n311), .B1(new_n316), .B2(new_n256), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n249), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT68), .ZN(new_n320));
  INV_X1    g0120(.A(new_n260), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(new_n249), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n320), .A2(new_n322), .B1(new_n202), .B2(new_n321), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n308), .B2(G169), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n310), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n301), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n271), .B1(G238), .B2(new_n275), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n278), .A2(new_n280), .A3(G232), .A4(G1698), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n278), .A2(new_n280), .A3(G226), .A4(new_n282), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n268), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT13), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n328), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n341), .A3(G169), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n335), .A2(KEYINPUT73), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n336), .B1(new_n328), .B2(new_n333), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n337), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n340), .B(new_n342), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n242), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n253), .B2(new_n256), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n351), .A2(KEYINPUT11), .A3(new_n249), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT12), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n321), .B2(new_n242), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n260), .A2(KEYINPUT12), .A3(G68), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n263), .A2(new_n242), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT11), .B1(new_n351), .B2(new_n249), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n352), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n349), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT9), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n324), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n318), .A2(KEYINPUT9), .A3(new_n323), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT10), .B1(new_n308), .B2(G190), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT71), .B1(new_n308), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n309), .A2(new_n369), .A3(G200), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n365), .A2(new_n366), .A3(new_n368), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n308), .A2(G190), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n367), .B2(new_n308), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT10), .B1(new_n373), .B2(new_n364), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n296), .A2(new_n300), .A3(KEYINPUT70), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n327), .A2(new_n360), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT74), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT72), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n338), .B2(G200), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n328), .A2(new_n336), .A3(new_n333), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n379), .B(G200), .C1(new_n381), .C2(new_n344), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n343), .A2(G190), .A3(new_n337), .A4(new_n346), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n358), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n378), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n380), .A2(new_n383), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n385), .A2(new_n358), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT74), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n377), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT76), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n314), .A2(new_n242), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n393), .A2(new_n201), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  AOI211_X1 g0196(.A(new_n396), .B(G20), .C1(new_n278), .C2(new_n280), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n285), .B2(new_n286), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT75), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n207), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n401), .B2(new_n396), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT16), .B(new_n395), .C1(new_n402), .C2(new_n242), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n287), .B2(G20), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n242), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n395), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n409), .A3(new_n249), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n316), .A2(new_n260), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n316), .B2(new_n264), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n278), .A2(new_n280), .A3(G226), .A4(G1698), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n278), .A2(new_n280), .A3(G223), .A4(new_n282), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n268), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n269), .B1(new_n290), .B2(new_n291), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n275), .A2(G232), .B1(new_n418), .B2(new_n274), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n417), .A2(new_n419), .A3(G190), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n367), .B1(new_n417), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n410), .A2(new_n412), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n392), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n410), .A2(new_n412), .A3(new_n422), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT76), .A3(KEYINPUT17), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n410), .A2(new_n412), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n428), .A2(KEYINPUT77), .A3(new_n424), .A4(new_n422), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n410), .A2(new_n424), .A3(new_n412), .A4(new_n422), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n425), .A2(new_n427), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n410), .A2(new_n412), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n417), .A2(new_n419), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(new_n298), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(G179), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT18), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n391), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n281), .A2(G303), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n278), .A2(new_n280), .A3(G264), .A4(G1698), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n278), .A2(new_n280), .A3(G257), .A4(new_n282), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT82), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n443), .A2(KEYINPUT82), .A3(new_n444), .A4(new_n445), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n292), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT5), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT79), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(G41), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n272), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n273), .A2(G1), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n456), .A2(new_n292), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G270), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n418), .A2(new_n454), .A3(new_n453), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  INV_X1    g0262(.A(G97), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n207), .C1(G33), .C2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n249), .C1(new_n207), .C2(G116), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G116), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n321), .A2(new_n468), .ZN(new_n469));
  AOI211_X1 g0269(.A(new_n249), .B(new_n321), .C1(new_n206), .C2(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G116), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n461), .A2(G179), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT84), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n473), .B(new_n474), .ZN(new_n475));
  OR3_X1    g0275(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n460), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT83), .B1(new_n450), .B2(new_n460), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(G169), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT21), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT21), .ZN(new_n482));
  AOI211_X1 g0282(.A(new_n482), .B(new_n479), .C1(new_n476), .C2(new_n477), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n475), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n472), .B1(new_n478), .B2(G200), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n295), .B2(new_n478), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n287), .A2(new_n207), .A3(G68), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT80), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n287), .A2(new_n490), .A3(new_n207), .A4(G68), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  INV_X1    g0292(.A(G87), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n492), .A2(new_n493), .B1(new_n331), .B2(new_n207), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT19), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G97), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n494), .A2(new_n495), .B1(new_n256), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n489), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(new_n249), .B1(new_n321), .B2(new_n255), .ZN(new_n499));
  INV_X1    g0299(.A(new_n255), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n470), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n499), .A2(KEYINPUT81), .A3(new_n501), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n287), .A2(G238), .A3(new_n282), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n287), .A2(G244), .A3(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n268), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n292), .B(G250), .C1(G1), .C2(new_n273), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n418), .A2(new_n455), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(G169), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n513), .B1(new_n509), .B2(new_n268), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n348), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n504), .A2(new_n505), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n470), .A2(G87), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n499), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(G190), .ZN(new_n521));
  INV_X1    g0321(.A(new_n516), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n278), .A2(new_n280), .A3(G257), .A4(G1698), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n278), .A2(new_n280), .A3(G250), .A4(new_n282), .ZN(new_n527));
  INV_X1    g0327(.A(G294), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n277), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n268), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n457), .A2(G264), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n459), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n367), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n533), .B(KEYINPUT88), .C1(G190), .C2(new_n532), .ZN(new_n534));
  AND2_X1   g0334(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n287), .A2(new_n207), .A3(G87), .A4(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n278), .A2(new_n280), .A3(new_n207), .A4(G87), .ZN(new_n537));
  NOR2_X1   g0337(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  INV_X1    g0341(.A(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(G20), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(KEYINPUT86), .B1(KEYINPUT23), .B2(G107), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT86), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n508), .A2(new_n541), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n207), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n536), .A2(new_n540), .A3(new_n544), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT24), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n548), .A2(new_n544), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT24), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n536), .A4(new_n540), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n262), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n260), .A2(G107), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n470), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(new_n542), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  OR3_X1    g0360(.A1(new_n532), .A2(KEYINPUT88), .A3(G190), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n534), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n542), .B1(new_n405), .B2(new_n406), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT6), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n564), .A2(new_n463), .A3(G107), .ZN(new_n565));
  XNOR2_X1  g0365(.A(G97), .B(G107), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n567), .A2(new_n207), .B1(new_n253), .B2(new_n252), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n249), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n321), .A2(new_n463), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n470), .A2(G97), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n457), .A2(G257), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n459), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n278), .A2(new_n280), .A3(G250), .A4(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n278), .A2(new_n280), .A3(G244), .A4(new_n282), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n462), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT78), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT78), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n582), .A3(new_n578), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n575), .B(G190), .C1(new_n584), .C2(new_n292), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n292), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(new_n574), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n572), .B(new_n585), .C1(new_n587), .C2(new_n367), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n575), .B(new_n348), .C1(new_n584), .C2(new_n292), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n587), .C2(G169), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n532), .A2(new_n298), .ZN(new_n592));
  OAI221_X1 g0392(.A(new_n592), .B1(G179), .B2(new_n532), .C1(new_n554), .C2(new_n559), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n562), .A2(new_n588), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  NOR4_X1   g0394(.A1(new_n442), .A2(new_n487), .A3(new_n525), .A4(new_n594), .ZN(G372));
  INV_X1    g0395(.A(new_n442), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n513), .A2(KEYINPUT89), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT89), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n511), .B2(new_n512), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n510), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n298), .B1(new_n348), .B2(new_n516), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n502), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n478), .A2(new_n480), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n482), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n473), .B(KEYINPUT84), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n478), .A2(KEYINPUT21), .A3(new_n480), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n593), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n600), .A2(G200), .B1(G190), .B2(new_n516), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n520), .A2(new_n610), .B1(new_n601), .B2(new_n502), .ZN(new_n611));
  AND4_X1   g0411(.A1(new_n591), .A2(new_n611), .A3(new_n588), .A4(new_n562), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n604), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n591), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n611), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n518), .A3(new_n524), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(KEYINPUT26), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n596), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n410), .A2(new_n412), .B1(new_n436), .B2(new_n437), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT18), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n388), .A2(new_n389), .ZN(new_n623));
  INV_X1    g0423(.A(new_n300), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(new_n359), .B2(new_n349), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(new_n433), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT10), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n308), .A2(new_n367), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(G190), .B2(new_n308), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n627), .B1(new_n629), .B2(new_n365), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n370), .A2(new_n368), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n366), .A2(new_n363), .A3(new_n362), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT90), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT90), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n371), .A2(new_n635), .A3(new_n374), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n326), .B1(new_n626), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n620), .A2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(new_n484), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n472), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n487), .B2(new_n647), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n593), .A2(new_n646), .ZN(new_n652));
  INV_X1    g0452(.A(new_n646), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n562), .B1(new_n560), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n654), .B2(new_n593), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n484), .A2(new_n646), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n655), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n210), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G1), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n492), .A2(new_n493), .A3(new_n468), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n665), .A2(new_n666), .B1(new_n219), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n619), .A2(new_n653), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n617), .A2(KEYINPUT26), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n615), .B1(new_n611), .B2(new_n614), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n646), .B1(new_n613), .B2(new_n672), .ZN(new_n673));
  MUX2_X1   g0473(.A(new_n669), .B(new_n673), .S(KEYINPUT29), .Z(new_n674));
  NOR2_X1   g0474(.A1(new_n594), .A2(new_n525), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n484), .A2(new_n675), .A3(new_n486), .A4(new_n653), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n461), .A2(G179), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n516), .A2(new_n531), .A3(new_n530), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n678), .A2(KEYINPUT30), .A3(new_n587), .A4(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n587), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n677), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n600), .A2(new_n348), .A3(new_n532), .ZN(new_n685));
  AOI211_X1 g0485(.A(new_n587), .B(new_n685), .C1(new_n476), .C2(new_n477), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n646), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g0489(.A(KEYINPUT31), .B(new_n646), .C1(new_n684), .C2(new_n686), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n676), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n674), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n668), .B1(new_n696), .B2(G1), .ZN(G364));
  AND2_X1   g0497(.A1(new_n207), .A2(G13), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n206), .B1(new_n698), .B2(G45), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n663), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n651), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(G330), .B2(new_n649), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n662), .A2(new_n281), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n704), .A2(G355), .B1(new_n468), .B2(new_n662), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n399), .A2(new_n400), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n662), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(G45), .B2(new_n219), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n246), .A2(new_n273), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n710), .A2(KEYINPUT91), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n213), .B1(G20), .B2(new_n298), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n710), .A2(KEYINPUT91), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n711), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n701), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n207), .A2(new_n348), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G200), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G190), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n721), .A2(new_n295), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n723), .A2(new_n242), .B1(new_n725), .B2(new_n202), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n295), .A2(G200), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n207), .B1(new_n727), .B2(new_n348), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n463), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n726), .A2(new_n281), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n720), .B(KEYINPUT92), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n727), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n730), .B1(new_n314), .B2(new_n733), .C1(new_n253), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n207), .A2(G179), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n295), .A3(G200), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT93), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G107), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G87), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n737), .A2(new_n734), .ZN(new_n748));
  INV_X1    g0548(.A(G159), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT32), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OR3_X1    g0550(.A1(new_n748), .A2(KEYINPUT32), .A3(new_n749), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n744), .A2(new_n747), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n748), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n753), .A2(G329), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n287), .B(new_n754), .C1(G326), .C2(new_n724), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n755), .B1(new_n735), .B2(new_n756), .C1(new_n757), .C2(new_n733), .ZN(new_n758));
  INV_X1    g0558(.A(new_n728), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n759), .A2(G294), .B1(new_n746), .B2(G303), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n760), .B1(new_n723), .B2(new_n761), .C1(new_n742), .C2(new_n762), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n736), .A2(new_n752), .B1(new_n758), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n719), .B1(new_n764), .B2(new_n715), .ZN(new_n765));
  INV_X1    g0565(.A(new_n714), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n718), .B(new_n765), .C1(new_n649), .C2(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n703), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(G396));
  XNOR2_X1  g0569(.A(new_n300), .B(KEYINPUT96), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n296), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n619), .A2(new_n653), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n669), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n266), .A2(new_n646), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n770), .A2(new_n296), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n300), .B2(new_n653), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n773), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n701), .B1(new_n778), .B2(new_n694), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n694), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n715), .A2(new_n712), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n701), .B1(G77), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n735), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G116), .B1(G303), .B2(new_n724), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n723), .A2(KEYINPUT94), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n723), .A2(KEYINPUT94), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n762), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT95), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n287), .B(new_n729), .C1(G311), .C2(new_n753), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n542), .B2(new_n745), .ZN(new_n792));
  INV_X1    g0592(.A(new_n733), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(G294), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n493), .B2(new_n742), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G137), .A2(new_n724), .B1(new_n722), .B2(G150), .ZN(new_n796));
  INV_X1    g0596(.A(G143), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n735), .B2(new_n749), .C1(new_n797), .C2(new_n733), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT34), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n743), .A2(G68), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n728), .A2(new_n314), .B1(new_n745), .B2(new_n202), .ZN(new_n803));
  INV_X1    g0603(.A(new_n706), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(G132), .C2(new_n753), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n790), .A2(new_n795), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n783), .B1(new_n807), .B2(new_n715), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n777), .B2(new_n713), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n780), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G384));
  INV_X1    g0611(.A(new_n567), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n812), .A2(KEYINPUT35), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(KEYINPUT35), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n813), .A2(new_n814), .A3(new_n468), .A4(new_n215), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n816));
  XNOR2_X1  g0616(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OR3_X1    g0617(.A1(new_n219), .A2(new_n253), .A3(new_n393), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n206), .B(G13), .C1(new_n818), .C2(new_n241), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n360), .A2(new_n646), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT39), .ZN(new_n823));
  INV_X1    g0623(.A(new_n644), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n403), .A2(new_n249), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n395), .B1(new_n402), .B2(new_n242), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT16), .B1(new_n826), .B2(KEYINPUT100), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT100), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n395), .C1(new_n402), .C2(new_n242), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n825), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n412), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n433), .B2(new_n440), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n438), .B1(new_n830), .B2(new_n831), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n832), .A2(new_n835), .A3(new_n426), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n836), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n434), .A2(new_n824), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n439), .A2(new_n838), .A3(new_n839), .A4(new_n426), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n836), .A2(KEYINPUT37), .B1(KEYINPUT101), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n834), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n834), .B(KEYINPUT38), .C1(new_n841), .C2(new_n837), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n823), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT103), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n423), .A2(new_n621), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n849), .A2(KEYINPUT103), .A3(new_n839), .A4(new_n838), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n439), .A2(new_n838), .A3(new_n426), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n848), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT76), .B1(new_n426), .B2(KEYINPUT17), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n426), .A2(KEYINPUT76), .A3(KEYINPUT17), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n430), .A2(new_n431), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n430), .A2(new_n431), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n854), .A2(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n838), .B1(new_n858), .B2(new_n622), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n843), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n845), .A2(new_n860), .A3(new_n823), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n846), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n845), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n836), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n826), .A2(KEYINPUT100), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n404), .A3(new_n829), .ZN(new_n867));
  INV_X1    g0667(.A(new_n825), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n412), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n423), .B1(new_n870), .B2(new_n824), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n839), .B1(new_n871), .B2(new_n835), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n840), .A2(KEYINPUT101), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n865), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n874), .B2(new_n834), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT39), .B1(new_n864), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(KEYINPUT102), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT104), .B1(new_n863), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n845), .A2(new_n860), .A3(new_n823), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(KEYINPUT102), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n846), .A2(new_n862), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n822), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n622), .A2(new_n824), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n864), .A2(new_n875), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n358), .A2(new_n653), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n388), .B2(new_n389), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n360), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n349), .B1(new_n390), .B2(new_n387), .ZN(new_n892));
  INV_X1    g0692(.A(new_n889), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT98), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n646), .B(new_n771), .C1(new_n613), .C2(new_n618), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n770), .A2(new_n646), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n898), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n773), .A2(KEYINPUT98), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n895), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT99), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n888), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g0704(.A(KEYINPUT99), .B(new_n895), .C1(new_n899), .C2(new_n901), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n886), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n884), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT105), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n674), .A2(new_n442), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n638), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n908), .B(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n676), .A2(new_n689), .A3(new_n690), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n913), .A2(new_n777), .A3(new_n894), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n845), .A2(new_n860), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n913), .A2(new_n777), .A3(new_n912), .A4(new_n894), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n845), .B2(new_n844), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n442), .B2(new_n691), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n913), .A2(new_n777), .A3(new_n894), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n845), .B2(new_n860), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n922), .A2(new_n912), .B1(new_n887), .B2(new_n917), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n596), .A3(new_n913), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n920), .A2(new_n924), .A3(G330), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n911), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n206), .B2(new_n698), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n911), .A2(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n820), .B1(new_n927), .B2(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n707), .A2(new_n231), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n716), .C1(new_n210), .C2(new_n255), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n701), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT108), .Z(new_n933));
  INV_X1    g0733(.A(new_n788), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(G294), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n743), .A2(G97), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n706), .B1(G317), .B2(new_n753), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n724), .A2(G311), .B1(new_n759), .B2(G107), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n746), .A2(G116), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT46), .ZN(new_n941));
  INV_X1    g0741(.A(G303), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n941), .B1(new_n762), .B2(new_n735), .C1(new_n942), .C2(new_n733), .ZN(new_n943));
  INV_X1    g0743(.A(G137), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n287), .B1(new_n944), .B2(new_n748), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n728), .A2(new_n242), .B1(new_n745), .B2(new_n314), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(G143), .C2(new_n724), .ZN(new_n947));
  INV_X1    g0747(.A(G150), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n947), .B1(new_n202), .B2(new_n735), .C1(new_n948), .C2(new_n733), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n743), .A2(G77), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n788), .B2(new_n749), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n939), .A2(new_n943), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT47), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n715), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n952), .A2(new_n953), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n520), .A2(new_n653), .ZN(new_n957));
  MUX2_X1   g0757(.A(new_n604), .B(new_n611), .S(new_n957), .Z(new_n958));
  OAI221_X1 g0758(.A(new_n933), .B1(new_n955), .B2(new_n956), .C1(new_n958), .C2(new_n766), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n657), .A2(new_n655), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n659), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(new_n650), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n695), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n591), .A2(new_n653), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT106), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n588), .B(new_n591), .C1(new_n572), .C2(new_n653), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n660), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT45), .Z(new_n969));
  NOR2_X1   g0769(.A1(new_n660), .A2(new_n967), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n656), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n656), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n963), .B(new_n974), .C1(new_n975), .C2(new_n973), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n696), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n663), .B(KEYINPUT41), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n700), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n980));
  INV_X1    g0780(.A(new_n967), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n591), .B1(new_n981), .B2(new_n593), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n653), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n981), .A2(new_n658), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT42), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n984), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n980), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n989), .B(new_n990), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n656), .A2(new_n981), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n959), .B1(new_n979), .B2(new_n993), .ZN(G387));
  INV_X1    g0794(.A(new_n715), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n723), .A2(new_n316), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n804), .B(new_n996), .C1(G150), .C2(new_n753), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n784), .A2(G68), .B1(new_n793), .B2(G50), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n745), .A2(new_n253), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n728), .A2(new_n255), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G159), .C2(new_n724), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n997), .A2(new_n998), .A3(new_n936), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n706), .B1(G326), .B2(new_n753), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n728), .A2(new_n762), .B1(new_n745), .B2(new_n528), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n784), .A2(G303), .B1(G322), .B2(new_n724), .ZN(new_n1005));
  INV_X1    g0805(.A(G317), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n733), .C1(new_n756), .C2(new_n788), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT48), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT49), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1003), .B1(new_n468), .B2(new_n742), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1002), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT110), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n995), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n1015), .B2(new_n1014), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n250), .A2(G50), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT109), .ZN(new_n1020));
  AOI211_X1 g0820(.A(G45), .B(new_n666), .C1(G68), .C2(G77), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1021), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(KEYINPUT109), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n707), .B1(new_n1022), .B2(new_n1024), .C1(new_n273), .C2(new_n236), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n704), .A2(new_n666), .B1(new_n542), .B2(new_n662), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n719), .B1(new_n1027), .B2(new_n716), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1017), .B(new_n1028), .C1(new_n655), .C2(new_n766), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n962), .A2(new_n695), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n663), .B1(new_n962), .B2(new_n695), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1029), .B1(new_n699), .B2(new_n962), .C1(new_n1030), .C2(new_n1031), .ZN(G393));
  OAI211_X1 g0832(.A(new_n976), .B(new_n663), .C1(new_n975), .C2(new_n963), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n981), .A2(new_n714), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n707), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n716), .B1(new_n463), .B2(new_n210), .C1(new_n1035), .C2(new_n240), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n701), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n934), .A2(G50), .B1(G87), .B2(new_n743), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n728), .A2(new_n253), .B1(new_n745), .B2(new_n242), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1039), .B(new_n804), .C1(G143), .C2(new_n753), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(new_n250), .C2(new_n735), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n733), .A2(new_n749), .B1(new_n948), .B2(new_n725), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT51), .Z(new_n1043));
  OAI22_X1  g0843(.A1(new_n733), .A2(new_n756), .B1(new_n1006), .B2(new_n725), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT52), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n934), .A2(G303), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n784), .A2(G294), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n745), .A2(new_n762), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n281), .B1(new_n748), .B2(new_n757), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(G116), .C2(new_n759), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1046), .A2(new_n744), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1041), .A2(new_n1043), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1037), .B1(new_n1052), .B2(new_n715), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n975), .A2(new_n700), .B1(new_n1034), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1033), .A2(new_n1054), .ZN(G390));
  NAND3_X1  g0855(.A1(new_n693), .A2(new_n777), .A3(new_n894), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n902), .A2(new_n821), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n898), .B1(new_n673), .B2(new_n772), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(new_n895), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n821), .B(KEYINPUT111), .Z(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n915), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1057), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n897), .A2(new_n896), .A3(new_n898), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT98), .B1(new_n773), .B2(new_n900), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n894), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n822), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n878), .A2(new_n883), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n1056), .A3(new_n1065), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1067), .A2(new_n700), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n878), .A2(new_n712), .A3(new_n883), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n463), .A2(new_n735), .B1(new_n733), .B2(new_n468), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n747), .B(new_n281), .C1(new_n528), .C2(new_n748), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n725), .A2(new_n762), .B1(new_n253), .B2(new_n728), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1079), .B(new_n802), .C1(new_n542), .C2(new_n788), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n724), .A2(G128), .B1(new_n759), .B2(G159), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n746), .A2(G150), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT53), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n934), .B2(G137), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT54), .B(G143), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n784), .A2(new_n1087), .B1(new_n793), .B2(G132), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1085), .B(new_n1088), .C1(KEYINPUT53), .C2(new_n1082), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n281), .B1(new_n753), .B2(G125), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n742), .B2(new_n202), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT113), .Z(new_n1092));
  OAI21_X1  g0892(.A(new_n1080), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n995), .B1(new_n1093), .B2(KEYINPUT114), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(KEYINPUT114), .B2(new_n1093), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n316), .A2(new_n781), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1075), .A2(new_n701), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1074), .A2(KEYINPUT115), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT115), .B1(new_n1074), .B2(new_n1097), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n596), .A2(new_n693), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n909), .A2(new_n638), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n777), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n895), .B1(new_n694), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(new_n1056), .A3(new_n1062), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1106), .A2(new_n1056), .B1(new_n899), .B2(new_n901), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1104), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n664), .B1(new_n1101), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1112), .A2(new_n1103), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1067), .A2(new_n1073), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT112), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1072), .A2(new_n1056), .A3(new_n1065), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1056), .B1(new_n1072), .B2(new_n1065), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1110), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AND4_X1   g0918(.A1(KEYINPUT112), .A2(new_n1118), .A3(new_n663), .A4(new_n1114), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1100), .B1(new_n1115), .B2(new_n1119), .ZN(G378));
  INV_X1    g0920(.A(new_n326), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n634), .A2(new_n1121), .A3(new_n636), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n324), .A2(new_n824), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT118), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1127));
  NAND4_X1  g0927(.A1(new_n634), .A2(new_n1121), .A3(new_n636), .A4(new_n1124), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n923), .A2(G330), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1127), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1132), .A2(KEYINPUT119), .A3(new_n1129), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1139), .B(G330), .C1(new_n916), .C2(new_n918), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1133), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n884), .B2(new_n906), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n821), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n919), .A2(new_n692), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1140), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n887), .B1(new_n1070), .B2(KEYINPUT99), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n902), .A2(new_n903), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n885), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1144), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1143), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n700), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n701), .B1(G50), .B2(new_n782), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G41), .B1(new_n753), .B2(G283), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n804), .B(new_n1155), .C1(new_n733), .C2(new_n542), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n500), .B2(new_n784), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n743), .A2(G58), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n999), .B1(G68), .B2(new_n759), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G97), .A2(new_n722), .B1(new_n724), .B2(G116), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT58), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n272), .B1(new_n804), .B2(new_n277), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1161), .A2(new_n1162), .B1(new_n202), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT116), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n722), .A2(G132), .B1(new_n746), .B2(new_n1087), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1166), .B1(new_n733), .B2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n724), .A2(G125), .B1(new_n759), .B2(G150), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT117), .Z(new_n1170));
  AOI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(G137), .C2(new_n784), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT59), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1174), .B1(new_n749), .B2(new_n742), .C1(new_n1171), .C2(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1165), .B1(new_n1162), .B2(new_n1161), .C1(new_n1173), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1154), .B1(new_n1177), .B2(new_n715), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1139), .B2(new_n713), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1153), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1114), .A2(new_n1104), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1143), .A2(new_n1150), .A3(KEYINPUT57), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n664), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1116), .A2(new_n1117), .A3(new_n1110), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1152), .B1(new_n1186), .B2(new_n1103), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1184), .A2(KEYINPUT120), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1182), .B1(new_n1114), .B2(new_n1104), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n664), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1180), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(G375));
  XOR2_X1   g0993(.A(new_n699), .B(KEYINPUT121), .Z(new_n1194));
  OR2_X1    g0994(.A1(new_n1112), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT122), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n701), .B1(G68), .B2(new_n782), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n895), .A2(new_n712), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT123), .Z(new_n1201));
  NAND2_X1  g1001(.A1(new_n934), .A2(new_n1087), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n724), .A2(G132), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n759), .A2(G50), .B1(new_n746), .B2(G159), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1202), .A2(new_n1158), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n804), .B1(G128), .B2(new_n753), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n735), .B2(new_n948), .C1(new_n944), .C2(new_n733), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n784), .A2(G107), .B1(new_n793), .B2(G283), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n287), .B(new_n1000), .C1(G303), .C2(new_n753), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n724), .A2(G294), .B1(new_n746), .B2(G97), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n950), .B1(new_n788), .B2(new_n468), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1205), .A2(new_n1207), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1199), .B(new_n1201), .C1(new_n715), .C2(new_n1213), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1197), .A2(new_n1198), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1112), .A2(new_n1103), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n1110), .A3(new_n978), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(G381));
  OR4_X1    g1018(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1219), .A2(G387), .A3(G381), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1111), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1100), .B1(new_n1186), .B2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G375), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1220), .A2(new_n1223), .ZN(G407));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n1220), .B2(new_n645), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(G213), .ZN(G409));
  OAI21_X1  g1026(.A(new_n1179), .B1(new_n1151), .B2(new_n1194), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1187), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n978), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1222), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(KEYINPUT120), .A3(new_n663), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1187), .A2(new_n1185), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1191), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1180), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(G378), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT124), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1234), .A2(G378), .A3(new_n1238), .A4(new_n1235), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1230), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT62), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1216), .B1(new_n1113), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1112), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n663), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1215), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n810), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1215), .A2(G384), .A3(new_n1245), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n645), .A2(G213), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NOR4_X1   g1051(.A1(new_n1240), .A2(new_n1241), .A3(new_n1249), .A4(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1240), .B2(KEYINPUT125), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1255), .B(new_n1230), .C1(new_n1237), .C2(new_n1239), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1254), .A2(new_n1249), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1253), .B1(new_n1257), .B2(KEYINPUT62), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1240), .A2(new_n1251), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1251), .A2(G2897), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1249), .B(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1259), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1258), .A2(KEYINPUT126), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1230), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1238), .B1(new_n1192), .B2(G378), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1239), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1255), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1249), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1240), .A2(KEYINPUT125), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .A4(new_n1250), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1252), .B1(new_n1274), .B2(new_n1241), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1266), .B1(new_n1275), .B2(new_n1263), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(G393), .B(new_n768), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(G390), .B(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(G387), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(KEYINPUT127), .Z(new_n1280));
  NAND3_X1  g1080(.A1(new_n1265), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1272), .A2(KEYINPUT63), .ZN(new_n1282));
  AOI211_X1 g1082(.A(KEYINPUT61), .B(new_n1279), .C1(new_n1260), .C2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n1262), .C1(KEYINPUT63), .C2(new_n1257), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(G405));
  OAI22_X1  g1086(.A1(new_n1268), .A2(new_n1269), .B1(new_n1192), .B2(new_n1222), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(new_n1272), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1280), .B(new_n1288), .ZN(G402));
endmodule


