//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n451), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(G2106), .ZN(G319));
  INV_X1    g033(.A(G125), .ZN(new_n459));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n466), .A2(new_n473), .ZN(G160));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(KEYINPUT67), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n460), .A2(KEYINPUT67), .A3(new_n461), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n467), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(KEYINPUT69), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n490), .B(new_n492), .C1(new_n476), .C2(new_n475), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n467), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n460), .B2(new_n461), .ZN(new_n496));
  XOR2_X1   g071(.A(KEYINPUT69), .B(KEYINPUT4), .Z(new_n497));
  OAI211_X1 g072(.A(new_n493), .B(new_n494), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n467), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT68), .A4(G2104), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n498), .A2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  OR3_X1    g094(.A1(new_n515), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n515), .B2(new_n518), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n510), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n526), .A2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n511), .A2(new_n534), .B1(new_n513), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(G171));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n511), .A2(new_n540), .B1(new_n513), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n517), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT71), .B1(new_n542), .B2(new_n544), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND3_X1  g130(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n510), .A2(new_n558), .A3(G53), .A4(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n509), .A2(new_n510), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G91), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n563));
  OAI21_X1  g138(.A(G65), .B1(new_n527), .B2(new_n528), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n566), .B2(G651), .ZN(new_n567));
  AOI211_X1 g142(.A(KEYINPUT72), .B(new_n517), .C1(new_n564), .C2(new_n565), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n560), .B(new_n562), .C1(new_n567), .C2(new_n568), .ZN(G299));
  OR2_X1    g144(.A1(new_n536), .A2(new_n538), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  OAI21_X1  g147(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n573));
  INV_X1    g148(.A(G49), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n573), .B1(new_n513), .B2(new_n574), .C1(new_n575), .C2(new_n511), .ZN(G288));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n511), .A2(new_n577), .B1(new_n513), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g154(.A1(G73), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n509), .B2(G61), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n517), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  AND2_X1   g159(.A1(new_n510), .A2(G543), .ZN(new_n585));
  AOI22_X1  g160(.A1(G85), .A2(new_n561), .B1(new_n585), .B2(G47), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n517), .B2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n511), .A2(KEYINPUT73), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT73), .B1(new_n511), .B2(new_n590), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n529), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(G651), .A2(new_n599), .B1(new_n585), .B2(G54), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n589), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n589), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  OAI21_X1  g184(.A(KEYINPUT74), .B1(new_n550), .B2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n601), .B2(new_n608), .ZN(new_n612));
  MUX2_X1   g187(.A(new_n610), .B(KEYINPUT74), .S(new_n612), .Z(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n471), .A2(G2104), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n481), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n483), .A2(G123), .ZN(new_n620));
  OR2_X1    g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n621), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT75), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G14), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n636), .A2(new_n639), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n637), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(KEYINPUT76), .B(KEYINPUT18), .Z(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2096), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT77), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  INV_X1    g233(.A(new_n648), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(new_n651), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1981), .B(G1986), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n671), .A2(new_n676), .A3(new_n674), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n676), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT78), .B(KEYINPUT20), .Z(new_n679));
  AOI211_X1 g254(.A(new_n675), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n678), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(KEYINPUT79), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(KEYINPUT79), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n668), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n684), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n682), .A3(new_n667), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n687), .ZN(G229));
  NOR2_X1   g263(.A1(G6), .A2(G16), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n583), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT32), .ZN(new_n691));
  INV_X1    g266(.A(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n694), .A2(KEYINPUT81), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(KEYINPUT81), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n703), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(G1971), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n693), .B(new_n706), .C1(G1971), .C2(new_n705), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n481), .A2(G131), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n483), .A2(G119), .ZN(new_n713));
  OR2_X1    g288(.A1(G95), .A2(G2105), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n717), .B2(new_n710), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT80), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n703), .A2(G24), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT82), .Z(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G290), .B2(new_n702), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1986), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(KEYINPUT83), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n720), .B2(new_n721), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n708), .A2(new_n709), .A3(new_n722), .A4(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n727), .A2(KEYINPUT83), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n710), .A2(G33), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n481), .A2(G139), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n460), .A2(new_n461), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n739), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n735), .B(new_n738), .C1(new_n467), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2072), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  INV_X1    g321(.A(G34), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G160), .B2(new_n710), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2084), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n752), .A2(KEYINPUT86), .A3(G28), .ZN(new_n753));
  AOI21_X1  g328(.A(KEYINPUT86), .B1(new_n752), .B2(G28), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n710), .B1(new_n752), .B2(G28), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n745), .A2(new_n751), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G4), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n601), .B2(G16), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n744), .B(new_n757), .C1(G1348), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n702), .A2(G19), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n550), .B2(new_n702), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1341), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n710), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n710), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(new_n764), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n764), .ZN(new_n770));
  INV_X1    g345(.A(new_n759), .ZN(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n710), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n467), .A2(G116), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n483), .A2(G128), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n481), .A2(G140), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(new_n710), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n710), .A2(G32), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n481), .A2(G141), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n483), .A2(G129), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT26), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n467), .A2(G2104), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n790), .B1(G105), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n785), .A2(new_n786), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n784), .B1(new_n793), .B2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT27), .B(G1996), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n783), .A2(G2067), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n783), .A2(G2067), .ZN(new_n797));
  NAND2_X1  g372(.A1(G286), .A2(G16), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n694), .A2(G21), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT84), .B(G1966), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n800), .A2(new_n802), .B1(new_n623), .B2(new_n710), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n694), .A2(G5), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G171), .B2(new_n694), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n805), .A2(G1961), .B1(new_n750), .B2(G2084), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n796), .A2(new_n797), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n760), .A2(new_n769), .A3(new_n773), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n710), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n710), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT29), .Z(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G2090), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n703), .A2(G20), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT89), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT23), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n694), .B2(new_n605), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1956), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n800), .A2(new_n802), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT85), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n794), .B2(new_n795), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n805), .A2(G1961), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT87), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n817), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n808), .A2(new_n812), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n732), .A2(new_n733), .A3(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n511), .A2(new_n827), .B1(new_n513), .B2(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n517), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n545), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n832), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n834), .B1(new_n549), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n608), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT90), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n835), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  INV_X1    g423(.A(KEYINPUT40), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n781), .B(G164), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n616), .B(KEYINPUT94), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n483), .A2(G130), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n467), .A2(KEYINPUT93), .A3(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT93), .B1(new_n467), .B2(G118), .ZN(new_n858));
  OR2_X1    g433(.A1(G106), .A2(G2105), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n857), .A2(G2104), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n481), .A2(G142), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT91), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n481), .A2(new_n864), .A3(G142), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n861), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n856), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT95), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n856), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n716), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n741), .B(new_n793), .Z(new_n873));
  AOI21_X1  g448(.A(new_n716), .B1(new_n868), .B2(new_n870), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n868), .A2(new_n870), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n717), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n878), .B2(new_n871), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n853), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n871), .A3(new_n876), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n852), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n623), .B(G160), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G162), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n880), .B2(new_n883), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n849), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n887), .A4(new_n886), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(G395));
  NAND2_X1  g468(.A1(G299), .A2(KEYINPUT97), .ZN(new_n894));
  OR2_X1    g469(.A1(G299), .A2(KEYINPUT97), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n601), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n838), .A2(KEYINPUT97), .A3(G299), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT96), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n601), .A2(new_n900), .A3(new_n608), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT96), .B1(new_n838), .B2(G559), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n836), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n836), .B1(new_n901), .B2(new_n902), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n899), .B(KEYINPUT98), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n896), .A2(KEYINPUT41), .A3(new_n897), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n907), .A2(new_n909), .A3(new_n903), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n903), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT98), .B1(new_n913), .B2(new_n899), .ZN(new_n914));
  XNOR2_X1  g489(.A(G166), .B(G288), .ZN(new_n915));
  XNOR2_X1  g490(.A(G290), .B(new_n583), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(G303), .A2(G288), .ZN(new_n919));
  NOR2_X1   g494(.A1(G166), .A2(new_n696), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT42), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n918), .A2(new_n921), .A3(KEYINPUT42), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n912), .A2(new_n914), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT98), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n925), .A2(new_n928), .A3(new_n911), .A4(new_n906), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n924), .A2(new_n929), .A3(G868), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT99), .B1(new_n835), .B2(new_n611), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n924), .A2(new_n929), .A3(KEYINPUT99), .A4(G868), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n932), .A2(KEYINPUT100), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT100), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(G295));
  AND2_X1   g511(.A1(new_n932), .A2(new_n933), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n549), .A2(new_n835), .ZN(new_n939));
  NAND2_X1  g514(.A1(G301), .A2(KEYINPUT101), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n941));
  NAND2_X1  g516(.A1(G171), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(G286), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(G171), .A2(new_n941), .A3(G168), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n939), .A2(new_n943), .A3(new_n833), .A4(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(KEYINPUT103), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(KEYINPUT103), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n833), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n944), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(KEYINPUT102), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT102), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n946), .B(new_n947), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n909), .A2(new_n910), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n915), .A2(new_n917), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n919), .A2(new_n920), .A3(new_n916), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n948), .A2(new_n949), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n945), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n948), .A2(KEYINPUT104), .A3(new_n949), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n899), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n955), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n887), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n953), .A2(new_n954), .B1(new_n899), .B2(new_n963), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n958), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n938), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n943), .A2(new_n944), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n970), .B1(new_n971), .B2(new_n836), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n950), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n973), .A2(new_n899), .A3(new_n947), .A4(new_n946), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n961), .A2(new_n909), .A3(new_n910), .A4(new_n962), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n958), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n967), .B2(new_n958), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(KEYINPUT105), .A3(new_n977), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n969), .B1(new_n983), .B2(new_n938), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT44), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n980), .A2(new_n981), .A3(new_n938), .A4(new_n982), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT43), .B1(new_n966), .B2(new_n968), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n985), .A2(new_n990), .ZN(G397));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n498), .B2(new_n507), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n465), .A2(G40), .A3(new_n470), .A4(new_n472), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n781), .B(G2067), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n793), .B(G1996), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n716), .B(new_n719), .Z(new_n1001));
  OR2_X1    g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(G290), .B(G1986), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n997), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT122), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  OR3_X1    g581(.A1(G168), .A2(KEYINPUT120), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT120), .B1(G168), .B2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(KEYINPUT51), .ZN(new_n1010));
  INV_X1    g585(.A(new_n996), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n502), .A2(new_n506), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT69), .B(KEYINPUT4), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n477), .B2(new_n495), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1012), .A2(new_n1014), .A3(new_n494), .A4(new_n493), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n995), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n801), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n996), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(G2084), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT106), .ZN(new_n1021));
  NOR2_X1   g596(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1015), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1019), .B(new_n1020), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1006), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1010), .B1(new_n1026), .B2(KEYINPUT121), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1028), .B(new_n1006), .C1(new_n1018), .C2(new_n1025), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1005), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1018), .A2(new_n1025), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1028), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1026), .A2(KEYINPUT121), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(KEYINPUT122), .A3(new_n1034), .A4(new_n1010), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT51), .B1(new_n1026), .B2(new_n1009), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1031), .A2(new_n1009), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n1017), .B2(G2078), .ZN(new_n1041));
  INV_X1    g616(.A(G1961), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1011), .B(new_n1043), .C1(new_n1024), .C2(new_n1023), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1041), .A2(KEYINPUT123), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n1040), .C1(new_n1017), .C2(G2078), .ZN(new_n1047));
  XOR2_X1   g622(.A(new_n473), .B(KEYINPUT124), .Z(new_n1048));
  NAND3_X1  g623(.A1(new_n767), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1048), .A2(new_n466), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(new_n995), .A3(new_n1016), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1045), .A2(G301), .A3(new_n1047), .A4(new_n1051), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1052), .A2(KEYINPUT125), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1041), .A2(KEYINPUT123), .ZN(new_n1054));
  OR3_X1    g629(.A1(new_n1017), .A2(new_n1040), .A3(G2078), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1044), .A2(new_n1042), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1054), .A2(new_n1047), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G171), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(KEYINPUT125), .A3(new_n1052), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1053), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  OAI221_X1 g637(.A(G8), .B1(G288), .B2(new_n1062), .C1(new_n996), .C2(new_n993), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT52), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1011), .A2(new_n992), .A3(new_n1015), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n696), .A2(G1976), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(G8), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(G61), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n529), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(G651), .B1(new_n1072), .B2(new_n580), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n561), .A2(G86), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n585), .A2(G48), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT109), .B(G1981), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1077), .A2(KEYINPUT110), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(KEYINPUT110), .ZN(new_n1079));
  OAI22_X1  g654(.A1(new_n1078), .A2(new_n1079), .B1(new_n692), .B2(new_n583), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1070), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI221_X1 g657(.A(KEYINPUT49), .B1(new_n692), .B2(new_n583), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1069), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(G166), .B2(new_n1006), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n520), .A2(G8), .A3(new_n521), .A4(new_n1085), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1971), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1017), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT107), .B(G2090), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1044), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1094), .A3(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1019), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1019), .A2(KEYINPUT111), .A3(new_n1096), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n1092), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1006), .B1(new_n1101), .B2(new_n1091), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1084), .B(new_n1095), .C1(new_n1102), .C2(new_n1089), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1057), .A2(G171), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1045), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1060), .B1(new_n1105), .B2(G171), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1039), .A2(new_n1061), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT72), .B1(new_n1109), .B2(new_n517), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n566), .A2(new_n563), .A3(G651), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1110), .A2(new_n1111), .B1(G91), .B2(new_n561), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1112), .B(new_n560), .C1(KEYINPUT114), .C2(KEYINPUT57), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT114), .B(new_n562), .C1(new_n567), .C2(new_n568), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n1115));
  NAND3_X1  g690(.A1(G299), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(G2072), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n995), .A2(new_n1011), .A3(new_n1016), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT113), .B(G1956), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1019), .B2(new_n1096), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1113), .B(new_n1116), .C1(new_n1120), .C2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n993), .A2(new_n996), .A3(G2067), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1044), .B2(new_n772), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n838), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1097), .A2(new_n1121), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1119), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1130), .A3(KEYINPUT61), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  NAND3_X1  g709(.A1(new_n1065), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n993), .B2(new_n996), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT116), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1135), .B(new_n1137), .C1(G1996), .C2(new_n1017), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n550), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1141), .A3(new_n550), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT117), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1147), .B(KEYINPUT61), .C1(new_n1124), .C2(new_n1130), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1132), .B(new_n1143), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n1151), .B(new_n1125), .C1(new_n1044), .C2(new_n772), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n601), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(KEYINPUT118), .A3(new_n838), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1150), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1131), .B1(new_n1149), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT119), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1162), .B(new_n1131), .C1(new_n1149), .C2(new_n1159), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1108), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1039), .A2(KEYINPUT62), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1037), .A2(new_n1166), .A3(new_n1038), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1103), .A2(new_n1058), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1171));
  NOR2_X1   g746(.A1(G288), .A2(G1976), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1084), .ZN(new_n1174));
  OAI22_X1  g749(.A1(new_n1173), .A2(new_n1070), .B1(new_n1174), .B2(new_n1095), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT112), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1032), .A2(G286), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1103), .B2(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1084), .A2(new_n1095), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1089), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1182), .A2(new_n1100), .B1(new_n1090), .B2(new_n1017), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n1183), .B2(new_n1006), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1180), .A2(KEYINPUT112), .A3(new_n1184), .A4(new_n1177), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1179), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1094), .A2(G8), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1181), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1180), .A2(KEYINPUT63), .A3(new_n1177), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1175), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1169), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1004), .B1(new_n1164), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n997), .B1(new_n998), .B2(new_n793), .ZN(new_n1194));
  NOR3_X1   g769(.A1(new_n995), .A2(G1996), .A3(new_n996), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT46), .Z(new_n1196));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT126), .Z(new_n1198));
  OR2_X1    g773(.A1(new_n1198), .A2(KEYINPUT47), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(KEYINPUT47), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1002), .A2(new_n997), .ZN(new_n1201));
  NOR2_X1   g776(.A1(G290), .A2(G1986), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n997), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n717), .A2(new_n719), .ZN(new_n1205));
  OAI22_X1  g780(.A1(new_n1000), .A2(new_n1205), .B1(G2067), .B2(new_n781), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1201), .A2(new_n1204), .B1(new_n997), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g782(.A1(new_n1199), .A2(new_n1200), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1193), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g784(.A1(new_n685), .A2(new_n687), .A3(G319), .A4(new_n661), .ZN(new_n1211));
  AOI211_X1 g785(.A(KEYINPUT127), .B(new_n1211), .C1(new_n642), .C2(new_n645), .ZN(new_n1212));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1213));
  INV_X1    g787(.A(new_n1211), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n646), .B2(new_n1214), .ZN(new_n1215));
  OAI22_X1  g789(.A1(new_n888), .A2(new_n889), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1216), .B1(new_n987), .B2(new_n986), .ZN(G308));
  OAI221_X1 g791(.A(new_n988), .B1(new_n889), .B2(new_n888), .C1(new_n1215), .C2(new_n1212), .ZN(G225));
endmodule


