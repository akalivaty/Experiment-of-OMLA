//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1203,
    new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(new_n466), .ZN(new_n476));
  OR3_X1    g051(.A1(new_n476), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  OR3_X1    g054(.A1(new_n478), .A2(KEYINPUT68), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(new_n478), .B2(new_n479), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n476), .A2(new_n461), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n461), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n483), .A2(G124), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(KEYINPUT69), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT69), .B1(new_n482), .B2(new_n487), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n467), .A2(G126), .A3(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n461), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n461), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  OR2_X1    g074(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G50), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n502), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G88), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n506), .B2(new_n512), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(G62), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n516), .B1(new_n521), .B2(G651), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  AOI211_X1 g098(.A(KEYINPUT71), .B(new_n523), .C1(new_n519), .C2(new_n520), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n514), .A2(new_n515), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  OAI221_X1 g102(.A(new_n527), .B1(new_n522), .B2(new_n524), .C1(new_n514), .C2(new_n515), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(G166));
  AOI22_X1  g104(.A1(new_n503), .A2(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT73), .B(G89), .Z(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n505), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n532), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n530), .A2(G90), .B1(new_n505), .B2(G52), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  OAI21_X1  g115(.A(G64), .B1(new_n517), .B2(new_n518), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n540), .B1(new_n543), .B2(G651), .ZN(new_n544));
  AOI211_X1 g119(.A(KEYINPUT74), .B(new_n523), .C1(new_n541), .C2(new_n542), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n508), .B2(new_n509), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT75), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n517), .A2(new_n518), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n553), .B(new_n550), .C1(new_n554), .C2(new_n548), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(G651), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n530), .A2(G81), .B1(new_n505), .B2(G43), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n554), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(new_n530), .B2(G91), .ZN(new_n571));
  AND2_X1   g146(.A1(KEYINPUT6), .A2(G651), .ZN(new_n572));
  NOR2_X1   g147(.A1(KEYINPUT6), .A2(G651), .ZN(new_n573));
  OAI211_X1 g148(.A(G53), .B(G543), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n511), .A2(new_n576), .A3(G53), .A4(G543), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  AND3_X1   g153(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n578), .B1(new_n575), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n571), .B1(new_n579), .B2(new_n580), .ZN(G299));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g157(.A1(G166), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n526), .A2(KEYINPUT78), .A3(new_n528), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n530), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n505), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT79), .B1(new_n554), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n510), .A2(new_n592), .A3(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G48), .B2(new_n505), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n530), .A2(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n554), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n601), .A2(KEYINPUT80), .A3(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT81), .B(G47), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n530), .A2(G85), .B1(new_n505), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(G543), .B1(new_n572), .B2(new_n573), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(KEYINPUT82), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n611), .B2(KEYINPUT82), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n554), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n612), .A2(new_n614), .B1(new_n617), .B2(G651), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n510), .A2(new_n511), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n610), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n610), .B1(new_n625), .B2(G868), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  INV_X1    g203(.A(G299), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G280));
  XOR2_X1   g205(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n561), .ZN(G323));
  XOR2_X1   g211(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n637));
  XNOR2_X1  g212(.A(G323), .B(new_n637), .ZN(G282));
  AND2_X1   g213(.A1(new_n475), .A2(new_n477), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G135), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n461), .A2(G111), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(KEYINPUT85), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n641), .B2(KEYINPUT85), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n642), .A2(new_n644), .B1(new_n483), .B2(G123), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT12), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT13), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(G2100), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(G2100), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  OR2_X1    g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT88), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n675), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n671), .B2(new_n674), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n671), .A3(new_n674), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(KEYINPUT18), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(KEYINPUT18), .ZN(new_n685));
  OAI221_X1 g260(.A(new_n678), .B1(new_n679), .B2(new_n681), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G2096), .B(G2100), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n690));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT20), .Z(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n692), .A2(new_n695), .A3(new_n698), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n697), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1991), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1981), .B(G1986), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT91), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n704), .B(new_n708), .ZN(G229));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G27), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT103), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n498), .B(KEYINPUT4), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n483), .A2(G126), .B1(new_n493), .B2(new_n495), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n712), .B1(new_n715), .B2(G29), .ZN(new_n716));
  INV_X1    g291(.A(G2078), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G34), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n719), .A2(KEYINPUT24), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(KEYINPUT24), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n710), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G160), .B2(new_n710), .ZN(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n710), .A2(G33), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT99), .B(KEYINPUT25), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n461), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G139), .B2(new_n639), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n726), .B1(new_n732), .B2(new_n710), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n734), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n725), .B1(G2072), .B2(new_n733), .C1(new_n736), .C2(G1961), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n718), .B(new_n737), .C1(G2072), .C2(new_n733), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n734), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(G1966), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n646), .A2(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(G1966), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  OR2_X1    g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n744), .A2(new_n710), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n742), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n741), .B(new_n748), .C1(G1961), .C2(new_n736), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT102), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT101), .B(KEYINPUT26), .Z(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n754), .B(new_n755), .Z(new_n756));
  AOI211_X1 g331(.A(new_n753), .B(new_n756), .C1(G129), .C2(new_n483), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n475), .A2(G141), .A3(new_n477), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT100), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G32), .B(new_n760), .S(G29), .Z(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT27), .B(G1996), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n738), .A2(new_n751), .A3(new_n752), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT104), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n752), .A2(new_n763), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT104), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n766), .A2(new_n767), .A3(new_n751), .A4(new_n738), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n771), .B(new_n772), .Z(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n734), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT106), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n629), .B2(new_n734), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n710), .A2(G26), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  OAI21_X1  g358(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n784));
  INV_X1    g359(.A(G116), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G2105), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT98), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(KEYINPUT98), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n787), .A2(new_n788), .B1(G128), .B2(new_n483), .ZN(new_n789));
  INV_X1    g364(.A(G140), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n478), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n783), .B1(new_n791), .B2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2067), .ZN(new_n793));
  NOR2_X1   g368(.A1(G4), .A2(G16), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n625), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT97), .B(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n561), .A2(new_n734), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n734), .B2(G19), .ZN(new_n799));
  INV_X1    g374(.A(G1341), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n793), .B(new_n797), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n781), .B(new_n801), .C1(new_n800), .C2(new_n799), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n769), .A2(new_n775), .A3(new_n776), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G16), .A2(G22), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G166), .B2(G16), .ZN(new_n805));
  INV_X1    g380(.A(G1971), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G6), .B(G305), .S(G16), .Z(new_n808));
  XOR2_X1   g383(.A(KEYINPUT32), .B(G1981), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n734), .A2(G23), .ZN(new_n811));
  INV_X1    g386(.A(G288), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n734), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT33), .B(G1976), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n813), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n807), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n710), .A2(G25), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n475), .A2(G131), .A3(new_n477), .ZN(new_n821));
  NOR2_X1   g396(.A1(G95), .A2(G2105), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT92), .ZN(new_n823));
  INV_X1    g398(.A(G107), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n463), .B1(new_n824), .B2(G2105), .ZN(new_n825));
  AOI22_X1  g400(.A1(G119), .A2(new_n483), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n820), .B1(new_n828), .B2(new_n710), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT93), .Z(new_n830));
  XOR2_X1   g405(.A(KEYINPUT35), .B(G1991), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n734), .A2(G24), .ZN(new_n835));
  INV_X1    g410(.A(new_n608), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n604), .B2(new_n605), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n837), .B2(new_n734), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1986), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n833), .A2(new_n834), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n819), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT95), .B1(new_n819), .B2(new_n840), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n818), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT36), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n818), .B(new_n848), .C1(new_n843), .C2(new_n844), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n803), .B1(new_n847), .B2(new_n849), .ZN(G311));
  AND4_X1   g425(.A1(new_n769), .A2(new_n775), .A3(new_n776), .A4(new_n802), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n841), .B(new_n842), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n848), .B1(new_n852), .B2(new_n818), .ZN(new_n853));
  INV_X1    g428(.A(new_n849), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(G150));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n620), .A2(new_n856), .B1(new_n857), .B2(new_n611), .ZN(new_n858));
  INV_X1    g433(.A(G67), .ZN(new_n859));
  INV_X1    g434(.A(G80), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n554), .A2(new_n859), .B1(new_n860), .B2(new_n502), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n523), .B1(new_n861), .B2(KEYINPUT107), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT107), .ZN(new_n863));
  OAI221_X1 g438(.A(new_n863), .B1(new_n860), .B2(new_n502), .C1(new_n554), .C2(new_n859), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n858), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n556), .A2(new_n558), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT76), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n556), .A2(new_n558), .A3(new_n557), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n861), .A2(KEYINPUT107), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(G651), .A3(new_n864), .ZN(new_n874));
  INV_X1    g449(.A(new_n858), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(new_n869), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n618), .A2(new_n624), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(new_n632), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n879), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT108), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n885), .B(new_n866), .C1(new_n883), .C2(new_n882), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n884), .A2(KEYINPUT108), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n868), .B1(new_n886), .B2(new_n887), .ZN(G145));
  INV_X1    g463(.A(new_n646), .ZN(new_n889));
  XOR2_X1   g464(.A(G160), .B(KEYINPUT109), .Z(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n489), .B2(new_n490), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR3_X1   g467(.A1(new_n489), .A2(new_n490), .A3(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(G162), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n646), .A3(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n732), .B1(new_n757), .B2(new_n759), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n757), .A2(new_n759), .A3(new_n732), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n828), .A2(KEYINPUT110), .ZN(new_n902));
  INV_X1    g477(.A(new_n649), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n827), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n903), .B1(new_n902), .B2(new_n905), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n900), .B(new_n901), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  INV_X1    g485(.A(new_n901), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n910), .B(new_n906), .C1(new_n911), .C2(new_n899), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n791), .A2(new_n715), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n791), .A2(new_n715), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n639), .A2(G142), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n461), .A2(G118), .ZN(new_n916));
  OAI21_X1  g491(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n483), .A2(G130), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n913), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n914), .B2(new_n913), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n909), .A2(new_n912), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n909), .B2(new_n912), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n898), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n924), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n897), .B(new_n894), .C1(new_n928), .C2(new_n925), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g507(.A(new_n878), .B(new_n634), .Z(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  AND2_X1   g509(.A1(G299), .A2(new_n880), .ZN(new_n935));
  NOR2_X1   g510(.A1(G299), .A2(new_n880), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n629), .A2(new_n625), .ZN(new_n938));
  NAND2_X1  g513(.A1(G299), .A2(new_n880), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT41), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n933), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n878), .B(new_n634), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n935), .A2(new_n936), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT42), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n944), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n933), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n948), .B(new_n949), .C1(new_n941), .C2(new_n933), .ZN(new_n950));
  XNOR2_X1  g525(.A(G290), .B(G305), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n526), .A2(new_n528), .A3(G288), .ZN(new_n952));
  NAND2_X1  g527(.A1(G166), .A2(new_n812), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(G305), .B(new_n837), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n526), .A2(new_n528), .A3(G288), .ZN(new_n956));
  AOI21_X1  g531(.A(G288), .B1(new_n526), .B2(new_n528), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n946), .A2(new_n950), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n946), .B2(new_n950), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n865), .A2(G868), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(G331));
  NOR2_X1   g539(.A1(G331), .A2(KEYINPUT111), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n962), .B2(new_n963), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n967), .ZN(G295));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(G301), .A2(G168), .ZN(new_n970));
  OAI211_X1 g545(.A(G286), .B(new_n539), .C1(new_n544), .C2(new_n545), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n872), .A2(new_n972), .A3(new_n877), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n876), .B1(new_n559), .B2(new_n560), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n865), .A2(new_n556), .A3(new_n558), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n974), .A2(new_n975), .B1(new_n970), .B2(new_n971), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n944), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(new_n872), .B2(new_n877), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n974), .A2(new_n975), .A3(new_n970), .A4(new_n971), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n937), .A4(new_n940), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT113), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n973), .A2(new_n976), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n941), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n959), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(KEYINPUT114), .A3(new_n930), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n977), .A2(new_n980), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n980), .A2(KEYINPUT113), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n988), .A2(new_n954), .A3(new_n958), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT114), .B1(new_n985), .B2(new_n930), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT43), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n977), .A2(new_n980), .B1(new_n954), .B2(new_n958), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(KEYINPUT115), .ZN(new_n995));
  AOI21_X1  g570(.A(G37), .B1(new_n994), .B2(KEYINPUT115), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n990), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n969), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n985), .A2(new_n930), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n986), .A4(new_n990), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n997), .B2(KEYINPUT43), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT116), .B1(new_n999), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1002), .A2(new_n986), .A3(new_n990), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(KEYINPUT43), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1009), .B(new_n1010), .C1(new_n1013), .C2(new_n969), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1008), .A2(new_n1014), .ZN(G397));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(G164), .B2(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G160), .A2(G40), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n760), .B(G1996), .ZN(new_n1020));
  INV_X1    g595(.A(G2067), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n791), .B(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n827), .B(new_n831), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(G290), .A2(G1986), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1019), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G8), .ZN(new_n1031));
  INV_X1    g606(.A(G40), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n470), .A2(new_n473), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n713), .B2(new_n714), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n596), .A2(new_n1036), .A3(new_n597), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT118), .B(G86), .Z(new_n1038));
  NAND2_X1  g613(.A1(new_n530), .A2(new_n1038), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n596), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1037), .B1(new_n1040), .B2(new_n1036), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT49), .B(new_n1037), .C1(new_n1040), .C2(new_n1036), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n1035), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n812), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1037), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1035), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1033), .B1(KEYINPUT45), .B2(new_n1034), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1034), .A2(KEYINPUT45), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G1971), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1034), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1033), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G2090), .ZN(new_n1058));
  OAI21_X1  g633(.A(G8), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n812), .A2(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1035), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1067), .A2(KEYINPUT117), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n1035), .B2(new_n1065), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1067), .B1(new_n1070), .B2(KEYINPUT117), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1045), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1049), .B1(new_n1064), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1966), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1054), .A2(new_n724), .A3(new_n1033), .A4(new_n1056), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(G168), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1031), .B1(KEYINPUT125), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1078), .A2(KEYINPUT125), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1077), .B(new_n1079), .C1(KEYINPUT125), .C2(new_n1078), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(G8), .A3(G286), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G303), .A2(G8), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(new_n1061), .A3(new_n1059), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1072), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1064), .A2(new_n1086), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1050), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1034), .A2(KEYINPUT45), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1093), .A2(KEYINPUT53), .A3(new_n717), .A4(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1017), .A2(new_n717), .A3(new_n1033), .A4(new_n1094), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1961), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1057), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G171), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1095), .A2(new_n1098), .A3(new_n1100), .A4(G301), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1103), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1092), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1052), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT121), .B(G1956), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1057), .A2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n575), .A2(new_n577), .ZN(new_n1114));
  INV_X1    g689(.A(new_n571), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(KEYINPUT57), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1114), .A2(new_n1116), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT123), .Z(new_n1118));
  NOR2_X1   g693(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1110), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT122), .B1(new_n1121), .B2(G2067), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1033), .A2(new_n1123), .A3(new_n1021), .A4(new_n1034), .ZN(new_n1124));
  INV_X1    g699(.A(G1348), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1122), .A2(new_n1124), .B1(new_n1057), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(new_n880), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1119), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1057), .A2(new_n1125), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1129), .B(new_n880), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1130), .A2(new_n1131), .A3(KEYINPUT124), .A4(KEYINPUT60), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n625), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT124), .B1(new_n1126), .B2(KEYINPUT60), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1050), .A2(new_n1051), .A3(G1996), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT58), .B(G1341), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n561), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT59), .ZN(new_n1146));
  OAI211_X1 g721(.A(KEYINPUT61), .B(new_n1120), .C1(new_n1113), .C2(new_n1118), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1110), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1117), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1128), .B1(new_n1141), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1073), .B1(new_n1108), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1089), .A2(new_n1061), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1072), .B1(new_n1155), .B2(new_n1060), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1102), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1156), .A2(new_n1090), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1086), .A2(KEYINPUT62), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1086), .A2(KEYINPUT62), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1162), .A2(new_n1156), .A3(new_n1090), .A4(new_n1157), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT126), .B1(new_n1164), .B2(new_n1160), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1154), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1031), .B(G286), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1059), .A2(KEYINPUT120), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1169), .B(G8), .C1(new_n1053), .C2(new_n1058), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1168), .A2(new_n1089), .A3(new_n1061), .A4(new_n1170), .ZN(new_n1171));
  AND4_X1   g746(.A1(KEYINPUT63), .A2(new_n1156), .A3(new_n1167), .A4(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1156), .A2(new_n1090), .A3(new_n1167), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT119), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1156), .A2(KEYINPUT119), .A3(new_n1090), .A4(new_n1167), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1172), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1030), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1019), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1179), .A2(new_n1027), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT48), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n1026), .B2(new_n1019), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT46), .ZN(new_n1183));
  OR3_X1    g758(.A1(new_n1179), .A2(new_n1183), .A3(G1996), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1019), .B1(new_n1023), .B2(new_n760), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1179), .B2(G1996), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT47), .Z(new_n1188));
  NAND3_X1  g763(.A1(new_n1024), .A2(new_n831), .A3(new_n828), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1189), .B1(G2067), .B2(new_n791), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1182), .B(new_n1188), .C1(new_n1019), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1178), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n688), .A2(G319), .A3(new_n669), .ZN(new_n1195));
  NOR2_X1   g769(.A1(G229), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n931), .A2(new_n1196), .ZN(new_n1197));
  NOR3_X1   g771(.A1(new_n1013), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n993), .A2(new_n998), .ZN(new_n1199));
  AND2_X1   g773(.A1(new_n931), .A2(new_n1196), .ZN(new_n1200));
  AOI21_X1  g774(.A(KEYINPUT127), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n1198), .A2(new_n1201), .ZN(G308));
  OAI21_X1  g776(.A(new_n1194), .B1(new_n1013), .B2(new_n1197), .ZN(new_n1203));
  NAND3_X1  g777(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT127), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1204), .ZN(G225));
endmodule


