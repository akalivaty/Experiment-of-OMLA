

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803;

  NAND2_X1 U371 ( .A1(n437), .A2(n458), .ZN(n350) );
  AND2_X1 U372 ( .A1(n621), .A2(n359), .ZN(n352) );
  AND2_X1 U373 ( .A1(n698), .A2(n422), .ZN(n477) );
  AND2_X1 U374 ( .A1(n385), .A2(n353), .ZN(n405) );
  XNOR2_X1 U375 ( .A(n365), .B(G122), .ZN(n556) );
  XNOR2_X1 U376 ( .A(n496), .B(G119), .ZN(n540) );
  NAND2_X1 U377 ( .A1(n438), .A2(n350), .ZN(n416) );
  XNOR2_X2 U378 ( .A(n547), .B(G134), .ZN(n559) );
  NAND2_X2 U379 ( .A1(n467), .A2(n717), .ZN(n425) );
  XOR2_X1 U380 ( .A(n660), .B(KEYINPUT28), .Z(n351) );
  AND2_X2 U381 ( .A1(n384), .A2(n394), .ZN(n391) );
  AND2_X2 U382 ( .A1(n421), .A2(n424), .ZN(n420) );
  AND2_X2 U383 ( .A1(n715), .A2(n364), .ZN(n469) );
  XNOR2_X2 U384 ( .A(n386), .B(G113), .ZN(n563) );
  INV_X2 U385 ( .A(G104), .ZN(n386) );
  NOR2_X2 U386 ( .A1(n383), .A2(n642), .ZN(n428) );
  XNOR2_X2 U387 ( .A(n714), .B(n713), .ZN(n468) );
  NAND2_X2 U388 ( .A1(n379), .A2(n377), .ZN(n714) );
  XNOR2_X2 U389 ( .A(n477), .B(n361), .ZN(n621) );
  INV_X1 U390 ( .A(n633), .ZN(n371) );
  XNOR2_X1 U391 ( .A(n793), .B(n537), .ZN(n742) );
  INV_X2 U392 ( .A(G953), .ZN(n454) );
  OR2_X1 U393 ( .A1(n694), .A2(n771), .ZN(n380) );
  XNOR2_X1 U394 ( .A(n664), .B(KEYINPUT46), .ZN(n381) );
  NAND2_X1 U395 ( .A1(n391), .A2(n390), .ZN(n654) );
  XNOR2_X1 U396 ( .A(n663), .B(n662), .ZN(n803) );
  AND2_X1 U397 ( .A1(n401), .A2(n488), .ZN(n395) );
  XNOR2_X1 U398 ( .A(n609), .B(n608), .ZN(n633) );
  XNOR2_X1 U399 ( .A(n448), .B(KEYINPUT1), .ZN(n698) );
  OR2_X1 U400 ( .A1(n659), .A2(n656), .ZN(n636) );
  AND2_X1 U401 ( .A1(n407), .A2(n414), .ZN(n413) );
  XNOR2_X1 U402 ( .A(n444), .B(n561), .ZN(n622) );
  XNOR2_X1 U403 ( .A(n525), .B(n524), .ZN(n659) );
  XNOR2_X1 U404 ( .A(n734), .B(n736), .ZN(n737) );
  XNOR2_X1 U405 ( .A(n453), .B(n562), .ZN(n732) );
  XNOR2_X1 U406 ( .A(n387), .B(n487), .ZN(n781) );
  XNOR2_X1 U407 ( .A(n519), .B(n518), .ZN(n453) );
  XNOR2_X1 U408 ( .A(n501), .B(KEYINPUT73), .ZN(n567) );
  XNOR2_X1 U409 ( .A(n516), .B(n515), .ZN(n519) );
  XNOR2_X1 U410 ( .A(G116), .B(KEYINPUT3), .ZN(n496) );
  XNOR2_X1 U411 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n506) );
  AND2_X1 U412 ( .A1(n385), .A2(n647), .ZN(n404) );
  XNOR2_X1 U413 ( .A(n428), .B(n360), .ZN(n385) );
  NAND2_X1 U414 ( .A1(n405), .A2(n406), .ZN(n401) );
  XNOR2_X2 U415 ( .A(n559), .B(n491), .ZN(n529) );
  AND2_X1 U416 ( .A1(n378), .A2(n706), .ZN(n377) );
  XNOR2_X1 U417 ( .A(n368), .B(n549), .ZN(n702) );
  NAND2_X1 U418 ( .A1(n748), .A2(n716), .ZN(n368) );
  INV_X1 U419 ( .A(KEYINPUT72), .ZN(n713) );
  NAND2_X1 U420 ( .A1(n633), .A2(n359), .ZN(n465) );
  INV_X1 U421 ( .A(n625), .ZN(n463) );
  NOR2_X1 U422 ( .A1(n621), .A2(n464), .ZN(n439) );
  OR2_X1 U423 ( .A1(n633), .A2(n359), .ZN(n464) );
  NAND2_X1 U424 ( .A1(n412), .A2(n411), .ZN(n410) );
  BUF_X1 U425 ( .A(n617), .Z(n593) );
  XNOR2_X1 U426 ( .A(n593), .B(KEYINPUT6), .ZN(n666) );
  INV_X1 U427 ( .A(G107), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n531), .B(G101), .ZN(n539) );
  XNOR2_X1 U429 ( .A(G110), .B(KEYINPUT93), .ZN(n531) );
  XNOR2_X1 U430 ( .A(n781), .B(n369), .ZN(n748) );
  XNOR2_X1 U431 ( .A(n546), .B(n548), .ZN(n486) );
  XNOR2_X1 U432 ( .A(n545), .B(n485), .ZN(n484) );
  NAND2_X1 U433 ( .A1(n710), .A2(n429), .ZN(n476) );
  NAND2_X1 U434 ( .A1(n778), .A2(n411), .ZN(n444) );
  NAND2_X1 U435 ( .A1(n742), .A2(G469), .ZN(n407) );
  XNOR2_X1 U436 ( .A(n510), .B(n509), .ZN(n792) );
  NAND2_X1 U437 ( .A1(n454), .A2(n575), .ZN(n501) );
  AND2_X1 U438 ( .A1(n493), .A2(KEYINPUT82), .ZN(n492) );
  XNOR2_X1 U439 ( .A(KEYINPUT68), .B(G131), .ZN(n507) );
  NAND2_X1 U440 ( .A1(n465), .A2(n689), .ZN(n389) );
  NOR2_X1 U441 ( .A1(n675), .A2(n607), .ZN(n609) );
  XOR2_X1 U442 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n554) );
  XNOR2_X1 U443 ( .A(n792), .B(n511), .ZN(n562) );
  INV_X1 U444 ( .A(G146), .ZN(n511) );
  XNOR2_X1 U445 ( .A(n475), .B(n473), .ZN(n472) );
  XNOR2_X1 U446 ( .A(n474), .B(G122), .ZN(n473) );
  XNOR2_X1 U447 ( .A(n563), .B(n564), .ZN(n475) );
  XNOR2_X1 U448 ( .A(G143), .B(KEYINPUT100), .ZN(n474) );
  XNOR2_X1 U449 ( .A(n529), .B(n530), .ZN(n793) );
  AND2_X1 U450 ( .A1(n666), .A2(n408), .ZN(n422) );
  AND2_X1 U451 ( .A1(n398), .A2(n396), .ZN(n390) );
  NAND2_X1 U452 ( .A1(n471), .A2(n623), .ZN(n665) );
  XNOR2_X1 U453 ( .A(n539), .B(n538), .ZN(n487) );
  XNOR2_X1 U454 ( .A(n388), .B(n540), .ZN(n387) );
  INV_X1 U455 ( .A(KEYINPUT16), .ZN(n538) );
  XNOR2_X1 U456 ( .A(n480), .B(n479), .ZN(n478) );
  INV_X1 U457 ( .A(KEYINPUT78), .ZN(n479) );
  NAND2_X1 U458 ( .A1(n481), .A2(n708), .ZN(n480) );
  INV_X1 U459 ( .A(KEYINPUT83), .ZN(n711) );
  NAND2_X1 U460 ( .A1(n460), .A2(n461), .ZN(n434) );
  INV_X1 U461 ( .A(n694), .ZN(n375) );
  NAND2_X1 U462 ( .A1(n374), .A2(n695), .ZN(n373) );
  XNOR2_X1 U463 ( .A(n456), .B(n550), .ZN(n650) );
  AND2_X1 U464 ( .A1(n650), .A2(n652), .ZN(n400) );
  NAND2_X1 U465 ( .A1(G469), .A2(G902), .ZN(n414) );
  XNOR2_X1 U466 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n497) );
  XNOR2_X1 U467 ( .A(G137), .B(G113), .ZN(n498) );
  XOR2_X1 U468 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n564) );
  XNOR2_X1 U469 ( .A(G902), .B(KEYINPUT15), .ZN(n716) );
  AND2_X1 U470 ( .A1(n492), .A2(n452), .ZN(n450) );
  XNOR2_X1 U471 ( .A(n543), .B(KEYINPUT17), .ZN(n545) );
  XNOR2_X1 U472 ( .A(G125), .B(KEYINPUT91), .ZN(n541) );
  XOR2_X1 U473 ( .A(KEYINPUT94), .B(KEYINPUT18), .Z(n542) );
  INV_X1 U474 ( .A(n650), .ZN(n397) );
  XNOR2_X1 U475 ( .A(n648), .B(n455), .ZN(n406) );
  INV_X1 U476 ( .A(KEYINPUT110), .ZN(n455) );
  INV_X1 U477 ( .A(n636), .ZN(n408) );
  XNOR2_X1 U478 ( .A(n366), .B(n556), .ZN(n388) );
  XNOR2_X1 U479 ( .A(n530), .B(n512), .ZN(n516) );
  NOR2_X1 U480 ( .A1(n440), .A2(G953), .ZN(n517) );
  INV_X1 U481 ( .A(G234), .ZN(n440) );
  AND2_X1 U482 ( .A1(n476), .A2(KEYINPUT64), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n641), .B(n482), .ZN(n481) );
  INV_X1 U484 ( .A(KEYINPUT81), .ZN(n482) );
  INV_X1 U485 ( .A(n707), .ZN(n367) );
  OR2_X1 U486 ( .A1(n766), .A2(n470), .ZN(n667) );
  NAND2_X1 U487 ( .A1(n666), .A2(n355), .ZN(n470) );
  NAND2_X1 U488 ( .A1(n462), .A2(n625), .ZN(n461) );
  NOR2_X1 U489 ( .A1(n352), .A2(n389), .ZN(n433) );
  INV_X1 U490 ( .A(n460), .ZN(n435) );
  BUF_X1 U491 ( .A(n702), .Z(n456) );
  XNOR2_X1 U492 ( .A(n668), .B(n602), .ZN(n675) );
  NAND2_X1 U493 ( .A1(n382), .A2(n355), .ZN(n660) );
  INV_X1 U494 ( .A(n795), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n558), .B(n445), .ZN(n778) );
  XNOR2_X1 U496 ( .A(n562), .B(n472), .ZN(n570) );
  XOR2_X1 U497 ( .A(G107), .B(G104), .Z(n535) );
  XNOR2_X1 U498 ( .A(n748), .B(n747), .ZN(n749) );
  NAND2_X1 U499 ( .A1(n654), .A2(n653), .ZN(n392) );
  XNOR2_X1 U500 ( .A(n615), .B(KEYINPUT32), .ZN(n370) );
  XNOR2_X1 U501 ( .A(n665), .B(KEYINPUT108), .ZN(n766) );
  AND2_X1 U502 ( .A1(n446), .A2(n358), .ZN(n483) );
  INV_X1 U503 ( .A(G122), .ZN(n415) );
  AND2_X1 U504 ( .A1(n647), .A2(KEYINPUT74), .ZN(n353) );
  OR2_X1 U505 ( .A1(n603), .A2(n601), .ZN(n354) );
  AND2_X1 U506 ( .A1(n659), .A2(n658), .ZN(n355) );
  AND2_X1 U507 ( .A1(n729), .A2(n640), .ZN(n356) );
  NAND2_X1 U508 ( .A1(n376), .A2(n375), .ZN(n357) );
  INV_X1 U509 ( .A(G902), .ZN(n411) );
  INV_X1 U510 ( .A(G237), .ZN(n575) );
  AND2_X1 U511 ( .A1(n354), .A2(n712), .ZN(n358) );
  XOR2_X1 U512 ( .A(KEYINPUT34), .B(KEYINPUT76), .Z(n359) );
  XOR2_X1 U513 ( .A(KEYINPUT111), .B(KEYINPUT30), .Z(n360) );
  XNOR2_X1 U514 ( .A(KEYINPUT90), .B(KEYINPUT33), .ZN(n361) );
  XNOR2_X1 U515 ( .A(n570), .B(n569), .ZN(n734) );
  NOR2_X1 U516 ( .A1(n716), .A2(KEYINPUT82), .ZN(n362) );
  XNOR2_X1 U517 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n363) );
  AND2_X1 U518 ( .A1(n362), .A2(n493), .ZN(n364) );
  INV_X1 U519 ( .A(KEYINPUT64), .ZN(n452) );
  INV_X1 U520 ( .A(n563), .ZN(n366) );
  AND2_X1 U521 ( .A1(n715), .A2(KEYINPUT2), .ZN(n710) );
  OR2_X1 U522 ( .A1(n715), .A2(n367), .ZN(n641) );
  AND2_X1 U523 ( .A1(n715), .A2(n454), .ZN(n783) );
  XNOR2_X2 U524 ( .A(n441), .B(n363), .ZN(n715) );
  XNOR2_X1 U525 ( .A(n486), .B(n484), .ZN(n369) );
  NAND2_X1 U526 ( .A1(n627), .A2(n370), .ZN(n443) );
  XNOR2_X1 U527 ( .A(n370), .B(G119), .ZN(G21) );
  NAND2_X1 U528 ( .A1(n371), .A2(n612), .ZN(n613) );
  NAND2_X1 U529 ( .A1(n371), .A2(n638), .ZN(n756) );
  NAND2_X1 U530 ( .A1(n373), .A2(n372), .ZN(n379) );
  NAND2_X1 U531 ( .A1(n357), .A2(n381), .ZN(n372) );
  INV_X1 U532 ( .A(n381), .ZN(n374) );
  NOR2_X1 U533 ( .A1(n771), .A2(KEYINPUT48), .ZN(n376) );
  NAND2_X1 U534 ( .A1(n380), .A2(KEYINPUT48), .ZN(n378) );
  INV_X1 U535 ( .A(n383), .ZN(n382) );
  NAND2_X1 U536 ( .A1(n383), .A2(n659), .ZN(n618) );
  XNOR2_X2 U537 ( .A(n617), .B(KEYINPUT106), .ZN(n383) );
  NAND2_X1 U538 ( .A1(n393), .A2(n400), .ZN(n384) );
  XNOR2_X2 U539 ( .A(n392), .B(n655), .ZN(n730) );
  INV_X1 U540 ( .A(n402), .ZN(n393) );
  NAND2_X1 U541 ( .A1(n395), .A2(n402), .ZN(n394) );
  NAND2_X1 U542 ( .A1(n402), .A2(n401), .ZN(n690) );
  NAND2_X1 U543 ( .A1(n397), .A2(n488), .ZN(n396) );
  NAND2_X1 U544 ( .A1(n399), .A2(n400), .ZN(n398) );
  INV_X1 U545 ( .A(n401), .ZN(n399) );
  NAND2_X2 U546 ( .A1(n403), .A2(n649), .ZN(n402) );
  NAND2_X1 U547 ( .A1(n404), .A2(n406), .ZN(n403) );
  NAND2_X1 U548 ( .A1(n408), .A2(n448), .ZN(n648) );
  AND2_X2 U549 ( .A1(n425), .A2(n452), .ZN(n418) );
  NAND2_X2 U550 ( .A1(n413), .A2(n409), .ZN(n448) );
  OR2_X1 U551 ( .A1(n742), .A2(n410), .ZN(n409) );
  INV_X1 U552 ( .A(G469), .ZN(n412) );
  NOR2_X1 U553 ( .A1(n416), .A2(n626), .ZN(n627) );
  XNOR2_X1 U554 ( .A(n416), .B(n415), .ZN(n802) );
  INV_X1 U555 ( .A(n425), .ZN(n421) );
  NAND2_X2 U556 ( .A1(n419), .A2(n417), .ZN(n776) );
  NOR2_X2 U557 ( .A1(n418), .A2(n426), .ZN(n417) );
  NAND2_X1 U558 ( .A1(n420), .A2(n423), .ZN(n419) );
  NAND2_X1 U559 ( .A1(n466), .A2(n492), .ZN(n424) );
  NAND2_X1 U560 ( .A1(n451), .A2(n427), .ZN(n426) );
  NAND2_X1 U561 ( .A1(n466), .A2(n450), .ZN(n427) );
  XNOR2_X2 U562 ( .A(n457), .B(n508), .ZN(n617) );
  NOR2_X1 U563 ( .A1(n709), .A2(KEYINPUT64), .ZN(n449) );
  INV_X1 U564 ( .A(n709), .ZN(n429) );
  XNOR2_X1 U565 ( .A(n709), .B(n430), .ZN(n794) );
  NAND2_X1 U566 ( .A1(n431), .A2(n434), .ZN(n438) );
  NAND2_X1 U567 ( .A1(n433), .A2(n432), .ZN(n431) );
  NAND2_X1 U568 ( .A1(n435), .A2(n439), .ZN(n432) );
  NOR2_X1 U569 ( .A1(n439), .A2(n352), .ZN(n437) );
  NAND2_X1 U570 ( .A1(n442), .A2(n356), .ZN(n441) );
  XNOR2_X1 U571 ( .A(n443), .B(n628), .ZN(n442) );
  XNOR2_X1 U572 ( .A(n559), .B(n557), .ZN(n445) );
  XNOR2_X1 U573 ( .A(n447), .B(n711), .ZN(n446) );
  NAND2_X1 U574 ( .A1(n478), .A2(n476), .ZN(n447) );
  NAND2_X1 U575 ( .A1(n351), .A2(n448), .ZN(n676) );
  NAND2_X1 U576 ( .A1(n449), .A2(n710), .ZN(n451) );
  NAND2_X1 U577 ( .A1(n719), .A2(n411), .ZN(n457) );
  XNOR2_X2 U578 ( .A(n529), .B(n489), .ZN(n719) );
  XNOR2_X1 U579 ( .A(n483), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U580 ( .A1(n459), .A2(n463), .ZN(n458) );
  INV_X1 U581 ( .A(n465), .ZN(n459) );
  NAND2_X1 U582 ( .A1(n689), .A2(n463), .ZN(n460) );
  INV_X1 U583 ( .A(n689), .ZN(n462) );
  NAND2_X1 U584 ( .A1(n468), .A2(n715), .ZN(n466) );
  NAND2_X1 U585 ( .A1(n469), .A2(n468), .ZN(n467) );
  INV_X1 U586 ( .A(n622), .ZN(n471) );
  INV_X1 U587 ( .A(n544), .ZN(n485) );
  INV_X1 U588 ( .A(n652), .ZN(n488) );
  XNOR2_X2 U589 ( .A(n490), .B(n503), .ZN(n489) );
  XNOR2_X2 U590 ( .A(n502), .B(n540), .ZN(n490) );
  XNOR2_X1 U591 ( .A(n544), .B(n507), .ZN(n491) );
  INV_X1 U592 ( .A(KEYINPUT2), .ZN(n493) );
  AND2_X1 U593 ( .A1(n686), .A2(n685), .ZN(n494) );
  XOR2_X1 U594 ( .A(n566), .B(n565), .Z(n495) );
  NOR2_X1 U595 ( .A1(n692), .A2(n763), .ZN(n693) );
  INV_X1 U596 ( .A(KEYINPUT44), .ZN(n628) );
  XNOR2_X1 U597 ( .A(n495), .B(n568), .ZN(n569) );
  INV_X1 U598 ( .A(n547), .ZN(n548) );
  INV_X1 U599 ( .A(KEYINPUT88), .ZN(n670) );
  XNOR2_X1 U600 ( .A(n670), .B(KEYINPUT36), .ZN(n671) );
  XNOR2_X1 U601 ( .A(n672), .B(n671), .ZN(n674) );
  INV_X1 U602 ( .A(KEYINPUT63), .ZN(n724) );
  XNOR2_X1 U603 ( .A(n498), .B(n497), .ZN(n500) );
  XOR2_X1 U604 ( .A(KEYINPUT99), .B(G101), .Z(n499) );
  XNOR2_X1 U605 ( .A(n500), .B(n499), .ZN(n503) );
  NAND2_X1 U606 ( .A1(n567), .A2(G210), .ZN(n502) );
  XNOR2_X2 U607 ( .A(KEYINPUT77), .B(G143), .ZN(n505) );
  INV_X1 U608 ( .A(G128), .ZN(n504) );
  XNOR2_X2 U609 ( .A(n505), .B(n504), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n506), .B(G146), .ZN(n544) );
  INV_X1 U611 ( .A(G472), .ZN(n508) );
  XNOR2_X1 U612 ( .A(G140), .B(G125), .ZN(n510) );
  XNOR2_X1 U613 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n509) );
  XNOR2_X2 U614 ( .A(KEYINPUT67), .B(G137), .ZN(n530) );
  XNOR2_X1 U615 ( .A(KEYINPUT69), .B(KEYINPUT23), .ZN(n512) );
  XNOR2_X1 U616 ( .A(G110), .B(G128), .ZN(n514) );
  XNOR2_X1 U617 ( .A(G119), .B(KEYINPUT24), .ZN(n513) );
  XNOR2_X1 U618 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U619 ( .A(KEYINPUT8), .B(n517), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n552), .A2(G221), .ZN(n518) );
  NAND2_X1 U621 ( .A1(n732), .A2(n411), .ZN(n525) );
  NAND2_X1 U622 ( .A1(n716), .A2(G234), .ZN(n521) );
  INV_X1 U623 ( .A(KEYINPUT20), .ZN(n520) );
  XNOR2_X1 U624 ( .A(n521), .B(n520), .ZN(n527) );
  INV_X1 U625 ( .A(n527), .ZN(n522) );
  NAND2_X1 U626 ( .A1(n522), .A2(G217), .ZN(n523) );
  XNOR2_X1 U627 ( .A(n523), .B(KEYINPUT25), .ZN(n524) );
  INV_X1 U628 ( .A(G221), .ZN(n526) );
  OR2_X1 U629 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U630 ( .A(n528), .B(KEYINPUT21), .ZN(n656) );
  NAND2_X1 U631 ( .A1(G227), .A2(n454), .ZN(n532) );
  XNOR2_X1 U632 ( .A(KEYINPUT97), .B(n532), .ZN(n533) );
  XNOR2_X1 U633 ( .A(n533), .B(G140), .ZN(n534) );
  XNOR2_X1 U634 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U635 ( .A(n539), .B(n536), .ZN(n537) );
  XNOR2_X1 U636 ( .A(n542), .B(n541), .ZN(n546) );
  AND2_X1 U637 ( .A1(G224), .A2(n454), .ZN(n543) );
  NAND2_X1 U638 ( .A1(n411), .A2(n575), .ZN(n551) );
  AND2_X1 U639 ( .A1(n551), .A2(G210), .ZN(n549) );
  INV_X1 U640 ( .A(KEYINPUT38), .ZN(n550) );
  NAND2_X1 U641 ( .A1(n551), .A2(G214), .ZN(n697) );
  NAND2_X1 U642 ( .A1(n650), .A2(n697), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G217), .A2(n552), .ZN(n553) );
  XNOR2_X1 U644 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U645 ( .A(n555), .B(KEYINPUT104), .Z(n558) );
  XNOR2_X1 U646 ( .A(G116), .B(n556), .ZN(n557) );
  INV_X1 U647 ( .A(KEYINPUT105), .ZN(n560) );
  XNOR2_X1 U648 ( .A(n560), .B(G478), .ZN(n561) );
  XOR2_X1 U649 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n566) );
  XNOR2_X1 U650 ( .A(G131), .B(KEYINPUT103), .ZN(n565) );
  NAND2_X1 U651 ( .A1(G214), .A2(n567), .ZN(n568) );
  NOR2_X1 U652 ( .A1(G902), .A2(n734), .ZN(n572) );
  XNOR2_X1 U653 ( .A(KEYINPUT13), .B(G475), .ZN(n571) );
  XNOR2_X1 U654 ( .A(n572), .B(n571), .ZN(n623) );
  NOR2_X1 U655 ( .A1(n622), .A2(n623), .ZN(n610) );
  INV_X1 U656 ( .A(n610), .ZN(n579) );
  NOR2_X1 U657 ( .A1(n581), .A2(n579), .ZN(n573) );
  XNOR2_X1 U658 ( .A(n573), .B(KEYINPUT41), .ZN(n661) );
  NOR2_X1 U659 ( .A1(n621), .A2(n661), .ZN(n574) );
  NOR2_X1 U660 ( .A1(G953), .A2(n574), .ZN(n712) );
  XOR2_X1 U661 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n577) );
  NAND2_X1 U662 ( .A1(G234), .A2(G237), .ZN(n576) );
  XNOR2_X1 U663 ( .A(n577), .B(n576), .ZN(n604) );
  NAND2_X1 U664 ( .A1(G952), .A2(n604), .ZN(n603) );
  NOR2_X1 U665 ( .A1(n650), .A2(n697), .ZN(n578) );
  NOR2_X1 U666 ( .A1(n579), .A2(n578), .ZN(n584) );
  INV_X1 U667 ( .A(n623), .ZN(n580) );
  NAND2_X1 U668 ( .A1(n622), .A2(n580), .ZN(n769) );
  NAND2_X1 U669 ( .A1(n665), .A2(n769), .ZN(n683) );
  INV_X1 U670 ( .A(n683), .ZN(n582) );
  NOR2_X1 U671 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U672 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U673 ( .A(KEYINPUT119), .B(n585), .Z(n586) );
  NOR2_X1 U674 ( .A1(n621), .A2(n586), .ZN(n599) );
  XOR2_X1 U675 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n588) );
  INV_X1 U676 ( .A(n698), .ZN(n673) );
  NAND2_X1 U677 ( .A1(n673), .A2(n636), .ZN(n587) );
  XOR2_X1 U678 ( .A(n588), .B(n587), .Z(n592) );
  INV_X1 U679 ( .A(n593), .ZN(n637) );
  NAND2_X1 U680 ( .A1(n659), .A2(n656), .ZN(n589) );
  XNOR2_X1 U681 ( .A(n589), .B(KEYINPUT49), .ZN(n590) );
  NOR2_X1 U682 ( .A1(n637), .A2(n590), .ZN(n591) );
  NAND2_X1 U683 ( .A1(n592), .A2(n591), .ZN(n595) );
  OR2_X1 U684 ( .A1(n593), .A2(n636), .ZN(n594) );
  OR2_X1 U685 ( .A1(n673), .A2(n594), .ZN(n634) );
  NAND2_X1 U686 ( .A1(n595), .A2(n634), .ZN(n596) );
  XNOR2_X1 U687 ( .A(KEYINPUT51), .B(n596), .ZN(n597) );
  NOR2_X1 U688 ( .A1(n661), .A2(n597), .ZN(n598) );
  NOR2_X1 U689 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U690 ( .A(n600), .B(KEYINPUT52), .ZN(n601) );
  NAND2_X1 U691 ( .A1(n702), .A2(n697), .ZN(n668) );
  INV_X1 U692 ( .A(KEYINPUT19), .ZN(n602) );
  NOR2_X1 U693 ( .A1(n603), .A2(G953), .ZN(n646) );
  XNOR2_X1 U694 ( .A(KEYINPUT95), .B(G898), .ZN(n786) );
  NAND2_X1 U695 ( .A1(G953), .A2(n786), .ZN(n782) );
  NAND2_X1 U696 ( .A1(G902), .A2(n604), .ZN(n643) );
  NOR2_X1 U697 ( .A1(n782), .A2(n643), .ZN(n605) );
  NOR2_X1 U698 ( .A1(n646), .A2(n605), .ZN(n606) );
  XNOR2_X1 U699 ( .A(n606), .B(KEYINPUT96), .ZN(n607) );
  INV_X1 U700 ( .A(KEYINPUT0), .ZN(n608) );
  INV_X1 U701 ( .A(n656), .ZN(n611) );
  AND2_X1 U702 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U703 ( .A(n613), .B(KEYINPUT22), .ZN(n616) );
  NOR2_X1 U704 ( .A1(n616), .A2(n666), .ZN(n629) );
  INV_X1 U705 ( .A(n659), .ZN(n631) );
  NOR2_X1 U706 ( .A1(n673), .A2(n631), .ZN(n614) );
  NAND2_X1 U707 ( .A1(n629), .A2(n614), .ZN(n615) );
  INV_X1 U708 ( .A(n616), .ZN(n620) );
  NOR2_X1 U709 ( .A1(n698), .A2(n618), .ZN(n619) );
  NAND2_X1 U710 ( .A1(n620), .A2(n619), .ZN(n728) );
  INV_X1 U711 ( .A(n728), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U713 ( .A(n624), .B(KEYINPUT107), .ZN(n689) );
  XOR2_X1 U714 ( .A(KEYINPUT35), .B(KEYINPUT75), .Z(n625) );
  NAND2_X1 U715 ( .A1(n629), .A2(n673), .ZN(n630) );
  XNOR2_X1 U716 ( .A(n630), .B(KEYINPUT87), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n729) );
  NOR2_X1 U718 ( .A1(n633), .A2(n634), .ZN(n635) );
  XNOR2_X1 U719 ( .A(n635), .B(KEYINPUT31), .ZN(n768) );
  NOR2_X1 U720 ( .A1(n648), .A2(n637), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n768), .A2(n756), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n639), .A2(n683), .ZN(n640) );
  XNOR2_X1 U723 ( .A(KEYINPUT2), .B(KEYINPUT79), .ZN(n707) );
  INV_X1 U724 ( .A(n697), .ZN(n642) );
  OR2_X1 U725 ( .A1(n454), .A2(n643), .ZN(n644) );
  NOR2_X1 U726 ( .A1(n644), .A2(G900), .ZN(n645) );
  NOR2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n657) );
  INV_X1 U728 ( .A(n657), .ZN(n647) );
  INV_X1 U729 ( .A(KEYINPUT74), .ZN(n649) );
  INV_X1 U730 ( .A(KEYINPUT86), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n651), .B(KEYINPUT39), .ZN(n652) );
  INV_X1 U732 ( .A(n665), .ZN(n653) );
  INV_X1 U733 ( .A(KEYINPUT40), .ZN(n655) );
  NOR2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n658) );
  OR2_X1 U735 ( .A1(n661), .A2(n676), .ZN(n663) );
  INV_X1 U736 ( .A(KEYINPUT42), .ZN(n662) );
  NOR2_X2 U737 ( .A1(n730), .A2(n803), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n667), .B(KEYINPUT109), .ZN(n696) );
  INV_X1 U739 ( .A(n668), .ZN(n669) );
  AND2_X1 U740 ( .A1(n696), .A2(n669), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n771) );
  INV_X1 U742 ( .A(n675), .ZN(n678) );
  INV_X1 U743 ( .A(n676), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n681) );
  NOR2_X1 U745 ( .A1(KEYINPUT47), .A2(n681), .ZN(n679) );
  NAND2_X1 U746 ( .A1(n683), .A2(n679), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT70), .ZN(n686) );
  NAND2_X1 U748 ( .A1(KEYINPUT80), .A2(n681), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n684), .A2(KEYINPUT47), .ZN(n685) );
  NAND2_X1 U751 ( .A1(n681), .A2(KEYINPUT47), .ZN(n688) );
  INV_X1 U752 ( .A(KEYINPUT80), .ZN(n687) );
  AND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n692) );
  AND2_X1 U754 ( .A1(n456), .A2(n689), .ZN(n691) );
  AND2_X1 U755 ( .A1(n690), .A2(n691), .ZN(n763) );
  NAND2_X1 U756 ( .A1(n494), .A2(n693), .ZN(n694) );
  INV_X1 U757 ( .A(KEYINPUT48), .ZN(n695) );
  NAND2_X1 U758 ( .A1(n696), .A2(n697), .ZN(n699) );
  NOR2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n701) );
  INV_X1 U760 ( .A(KEYINPUT43), .ZN(n700) );
  XNOR2_X1 U761 ( .A(n701), .B(n700), .ZN(n704) );
  INV_X1 U762 ( .A(n456), .ZN(n703) );
  AND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n774) );
  INV_X1 U764 ( .A(n769), .ZN(n705) );
  AND2_X1 U765 ( .A1(n654), .A2(n705), .ZN(n726) );
  NOR2_X1 U766 ( .A1(n774), .A2(n726), .ZN(n706) );
  BUF_X1 U767 ( .A(n714), .Z(n709) );
  NAND2_X1 U768 ( .A1(n709), .A2(n707), .ZN(n708) );
  NAND2_X1 U769 ( .A1(n716), .A2(KEYINPUT82), .ZN(n717) );
  NAND2_X1 U770 ( .A1(n776), .A2(G472), .ZN(n721) );
  XOR2_X1 U771 ( .A(KEYINPUT112), .B(KEYINPUT62), .Z(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n723) );
  INV_X1 U774 ( .A(G952), .ZN(n722) );
  AND2_X1 U775 ( .A1(n722), .A2(G953), .ZN(n780) );
  NOR2_X2 U776 ( .A1(n723), .A2(n780), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n725), .B(n724), .ZN(G57) );
  XOR2_X1 U778 ( .A(G134), .B(n726), .Z(G36) );
  XOR2_X1 U779 ( .A(G110), .B(KEYINPUT113), .Z(n727) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(G12) );
  XNOR2_X1 U781 ( .A(n729), .B(G101), .ZN(G3) );
  XOR2_X1 U782 ( .A(n730), .B(G131), .Z(G33) );
  NAND2_X1 U783 ( .A1(n776), .A2(G217), .ZN(n731) );
  XOR2_X1 U784 ( .A(n732), .B(n731), .Z(n733) );
  NOR2_X1 U785 ( .A1(n733), .A2(n780), .ZN(G66) );
  NAND2_X1 U786 ( .A1(n776), .A2(G475), .ZN(n738) );
  XNOR2_X1 U787 ( .A(KEYINPUT92), .B(KEYINPUT121), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n735), .B(KEYINPUT59), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X2 U790 ( .A1(n739), .A2(n780), .ZN(n740) );
  XNOR2_X1 U791 ( .A(n740), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U792 ( .A1(n776), .A2(G469), .ZN(n744) );
  XOR2_X1 U793 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n741) );
  XNOR2_X1 U794 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U795 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U796 ( .A1(n745), .A2(n780), .ZN(G54) );
  NAND2_X1 U797 ( .A1(n776), .A2(G210), .ZN(n750) );
  XOR2_X1 U798 ( .A(KEYINPUT89), .B(KEYINPUT54), .Z(n746) );
  XNOR2_X1 U799 ( .A(n746), .B(KEYINPUT55), .ZN(n747) );
  XNOR2_X1 U800 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X2 U801 ( .A1(n751), .A2(n780), .ZN(n754) );
  XNOR2_X1 U802 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n752) );
  XOR2_X1 U803 ( .A(n752), .B(KEYINPUT85), .Z(n753) );
  XNOR2_X1 U804 ( .A(n754), .B(n753), .ZN(G51) );
  NOR2_X1 U805 ( .A1(n756), .A2(n766), .ZN(n755) );
  XOR2_X1 U806 ( .A(G104), .B(n755), .Z(G6) );
  NOR2_X1 U807 ( .A1(n756), .A2(n769), .ZN(n758) );
  XNOR2_X1 U808 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n757) );
  XNOR2_X1 U809 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U810 ( .A(G107), .B(n759), .ZN(G9) );
  NOR2_X1 U811 ( .A1(n769), .A2(n681), .ZN(n761) );
  XNOR2_X1 U812 ( .A(KEYINPUT29), .B(KEYINPUT114), .ZN(n760) );
  XNOR2_X1 U813 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U814 ( .A(G128), .B(n762), .ZN(G30) );
  XOR2_X1 U815 ( .A(G143), .B(n763), .Z(G45) );
  NOR2_X1 U816 ( .A1(n766), .A2(n681), .ZN(n765) );
  XNOR2_X1 U817 ( .A(G146), .B(KEYINPUT115), .ZN(n764) );
  XNOR2_X1 U818 ( .A(n765), .B(n764), .ZN(G48) );
  NOR2_X1 U819 ( .A1(n766), .A2(n768), .ZN(n767) );
  XOR2_X1 U820 ( .A(G113), .B(n767), .Z(G15) );
  NOR2_X1 U821 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U822 ( .A(G116), .B(n770), .Z(G18) );
  XNOR2_X1 U823 ( .A(n771), .B(KEYINPUT116), .ZN(n772) );
  XNOR2_X1 U824 ( .A(n772), .B(KEYINPUT37), .ZN(n773) );
  XNOR2_X1 U825 ( .A(G125), .B(n773), .ZN(G27) );
  XNOR2_X1 U826 ( .A(G140), .B(n774), .ZN(n775) );
  XNOR2_X1 U827 ( .A(n775), .B(KEYINPUT117), .ZN(G42) );
  NAND2_X1 U828 ( .A1(n776), .A2(G478), .ZN(n777) );
  XOR2_X1 U829 ( .A(n778), .B(n777), .Z(n779) );
  NOR2_X1 U830 ( .A1(n780), .A2(n779), .ZN(G63) );
  NAND2_X1 U831 ( .A1(n782), .A2(n781), .ZN(n791) );
  XOR2_X1 U832 ( .A(KEYINPUT123), .B(n783), .Z(n789) );
  NAND2_X1 U833 ( .A1(G953), .A2(G224), .ZN(n784) );
  XOR2_X1 U834 ( .A(KEYINPUT61), .B(n784), .Z(n785) );
  NOR2_X1 U835 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U836 ( .A(KEYINPUT122), .B(n787), .ZN(n788) );
  NOR2_X1 U837 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U838 ( .A(n791), .B(n790), .ZN(G69) );
  XNOR2_X1 U839 ( .A(n793), .B(n792), .ZN(n795) );
  NAND2_X1 U840 ( .A1(n794), .A2(n454), .ZN(n801) );
  XOR2_X1 U841 ( .A(G227), .B(n795), .Z(n796) );
  XNOR2_X1 U842 ( .A(n796), .B(KEYINPUT124), .ZN(n797) );
  NAND2_X1 U843 ( .A1(n797), .A2(G900), .ZN(n798) );
  XOR2_X1 U844 ( .A(KEYINPUT125), .B(n798), .Z(n799) );
  NAND2_X1 U845 ( .A1(G953), .A2(n799), .ZN(n800) );
  NAND2_X1 U846 ( .A1(n801), .A2(n800), .ZN(G72) );
  XNOR2_X1 U847 ( .A(KEYINPUT126), .B(n802), .ZN(G24) );
  XOR2_X1 U848 ( .A(G137), .B(n803), .Z(G39) );
endmodule

