//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT21), .B(G898), .Z(new_n190));
  NAND3_X1  g004(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT82), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT3), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G107), .ZN(new_n201));
  OR3_X1    g015(.A1(new_n193), .A2(KEYINPUT3), .A3(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G101), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n199), .A2(new_n201), .A3(new_n205), .A4(new_n202), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n207));
  XOR2_X1   g021(.A(G116), .B(G119), .Z(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT2), .B(G113), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT2), .B(G113), .Z(new_n211));
  XNOR2_X1  g025(.A(G116), .B(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT4), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n203), .A2(new_n215), .A3(G101), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n198), .B1(G104), .B2(new_n197), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n206), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT5), .ZN(new_n221));
  INV_X1    g035(.A(G119), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G116), .ZN(new_n223));
  OAI211_X1 g037(.A(G113), .B(new_n223), .C1(new_n208), .C2(new_n221), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n213), .ZN(new_n225));
  OR3_X1    g039(.A1(new_n220), .A2(KEYINPUT84), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT84), .B1(new_n220), .B2(new_n225), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n217), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(G110), .B(G122), .Z(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT85), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT6), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n229), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n217), .A2(new_n226), .A3(new_n234), .A4(new_n227), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n228), .A2(new_n231), .A3(KEYINPUT6), .A4(new_n229), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT65), .B1(new_n238), .B2(G146), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT64), .B(G146), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n240), .B(new_n243), .C1(new_n244), .C2(new_n238), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n238), .A2(G146), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n244), .B2(new_n238), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI22_X1  g063(.A1(new_n245), .A2(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G125), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n238), .A2(KEYINPUT65), .A3(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(G143), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT1), .B1(new_n244), .B2(new_n238), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G128), .A4(new_n240), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n253), .A2(new_n255), .A3(new_n238), .ZN(new_n260));
  INV_X1    g074(.A(new_n247), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n256), .B2(G143), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n251), .B1(new_n267), .B2(G125), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n188), .A2(G224), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(KEYINPUT7), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n251), .B(new_n271), .C1(new_n267), .C2(G125), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n220), .A2(KEYINPUT86), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n225), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n229), .B(KEYINPUT8), .Z(new_n278));
  OAI211_X1 g092(.A(new_n213), .B(new_n224), .C1(new_n220), .C2(KEYINPUT86), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n275), .A2(new_n235), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n281), .B2(new_n283), .ZN(new_n285));
  OAI22_X1  g099(.A1(new_n237), .A2(new_n270), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(KEYINPUT88), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n291));
  INV_X1    g105(.A(new_n270), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n293), .B(new_n287), .C1(new_n285), .C2(new_n284), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G475), .ZN(new_n299));
  XNOR2_X1  g113(.A(G125), .B(G140), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n256), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT76), .B1(new_n256), .B2(new_n300), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n303), .A2(new_n304), .B1(new_n241), .B2(new_n300), .ZN(new_n305));
  OR2_X1    g119(.A1(KEYINPUT70), .A2(G237), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT70), .A2(G237), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(G214), .A3(new_n188), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n238), .ZN(new_n310));
  AOI21_X1  g124(.A(G953), .B1(new_n306), .B2(new_n307), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(G143), .A3(G214), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT18), .A2(G131), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT18), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n316), .B(new_n317), .C1(new_n310), .C2(new_n312), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT89), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n310), .A2(new_n312), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT18), .A3(G131), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT89), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n314), .A4(new_n305), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G113), .B(G122), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(new_n193), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(G131), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT17), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n310), .A2(new_n317), .A3(new_n312), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n331), .A2(KEYINPUT16), .A3(G140), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n300), .B2(KEYINPUT16), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n333), .A2(G146), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(G146), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT90), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n320), .A2(KEYINPUT17), .A3(G131), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n335), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT90), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n330), .A2(new_n336), .A3(new_n337), .A4(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n324), .A2(new_n326), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n327), .A2(new_n329), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n300), .B(KEYINPUT19), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n256), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n335), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n326), .B1(new_n324), .B2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n299), .B(new_n283), .C1(new_n343), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT20), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(new_n347), .ZN(new_n351));
  INV_X1    g165(.A(new_n326), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n342), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n299), .A4(new_n283), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n326), .B1(new_n324), .B2(new_n341), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n283), .B1(new_n343), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G475), .ZN(new_n360));
  XNOR2_X1  g174(.A(G116), .B(G122), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n197), .ZN(new_n362));
  INV_X1    g176(.A(G116), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT14), .A3(G122), .ZN(new_n364));
  INV_X1    g178(.A(new_n361), .ZN(new_n365));
  OAI211_X1 g179(.A(G107), .B(new_n364), .C1(new_n365), .C2(KEYINPUT14), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n265), .B2(G143), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n238), .A2(KEYINPUT91), .A3(G128), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n265), .A2(G143), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT92), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(KEYINPUT92), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G134), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n376), .A2(new_n377), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n362), .B(new_n366), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n365), .A2(G107), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n376), .A2(new_n377), .B1(new_n382), .B2(new_n362), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n370), .A2(new_n384), .B1(new_n265), .B2(G143), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n384), .B2(new_n370), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G134), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(KEYINPUT93), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT93), .B1(new_n383), .B2(new_n387), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n381), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT73), .B(G217), .Z(new_n392));
  XOR2_X1   g206(.A(KEYINPUT9), .B(G234), .Z(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(new_n188), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n390), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n388), .ZN(new_n397));
  INV_X1    g211(.A(new_n394), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n381), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n283), .ZN(new_n401));
  INV_X1    g215(.A(G478), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT15), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n400), .B(new_n283), .C1(KEYINPUT15), .C2(new_n402), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n357), .A2(new_n360), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n393), .A2(new_n283), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n408), .A2(G221), .ZN(new_n409));
  INV_X1    g223(.A(G469), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(new_n283), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n188), .A2(G227), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(G140), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT81), .B(G110), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n238), .B1(new_n253), .B2(new_n255), .ZN(new_n416));
  OAI21_X1  g230(.A(G128), .B1(new_n416), .B2(new_n263), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(new_n245), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n265), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n257), .B2(new_n240), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n206), .B(new_n219), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n249), .B1(new_n260), .B2(new_n261), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n416), .A2(new_n239), .A3(new_n252), .ZN(new_n425));
  INV_X1    g239(.A(new_n246), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n207), .A2(new_n427), .A3(new_n216), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n267), .A2(KEYINPUT10), .A3(new_n206), .A4(new_n219), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G137), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(G134), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(G134), .ZN(new_n433));
  NAND2_X1  g247(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n431), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n435), .A2(new_n317), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n434), .B1(new_n377), .B2(G137), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n377), .A2(G137), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n439), .A2(new_n437), .A3(new_n436), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G131), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n430), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n441), .B(new_n317), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n423), .A2(new_n428), .A3(new_n445), .A4(new_n429), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n415), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n220), .A2(new_n266), .A3(new_n259), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n421), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n445), .B2(KEYINPUT83), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n450), .A2(new_n443), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n452), .B1(new_n450), .B2(new_n443), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n446), .B(new_n415), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n411), .B1(new_n456), .B2(new_n410), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n446), .A2(new_n415), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n446), .B1(new_n453), .B2(new_n454), .ZN(new_n460));
  INV_X1    g274(.A(new_n415), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n459), .A2(new_n444), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G469), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n409), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  AND4_X1   g278(.A1(new_n192), .A2(new_n298), .A3(new_n407), .A4(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G472), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n433), .A2(new_n440), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G131), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n441), .B2(G131), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n258), .A2(G128), .B1(new_n261), .B2(new_n260), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n418), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n425), .A2(new_n426), .ZN(new_n473));
  INV_X1    g287(.A(new_n424), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n443), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n210), .A2(new_n213), .A3(KEYINPUT68), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT68), .B1(new_n210), .B2(new_n213), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n472), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT28), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n472), .A2(new_n475), .B1(new_n210), .B2(new_n213), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n267), .A2(new_n470), .B1(new_n427), .B2(new_n443), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT69), .B1(new_n485), .B2(new_n478), .ZN(new_n486));
  AND4_X1   g300(.A1(KEYINPUT69), .A2(new_n472), .A3(new_n475), .A4(new_n478), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n482), .B1(new_n488), .B2(KEYINPUT28), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n311), .A2(G210), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(G101), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT29), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n445), .A2(new_n250), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n469), .B1(new_n259), .B2(new_n266), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n498));
  OR2_X1    g312(.A1(KEYINPUT67), .A2(KEYINPUT30), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n472), .A2(new_n475), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n479), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n485), .A2(KEYINPUT69), .A3(new_n478), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n501), .A2(new_n214), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n494), .B1(new_n505), .B2(new_n493), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n504), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n485), .B2(new_n478), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n482), .B1(new_n508), .B2(KEYINPUT28), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n493), .A2(KEYINPUT29), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n466), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT71), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n489), .B2(new_n493), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT31), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n505), .A2(new_n516), .A3(new_n493), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n505), .A2(new_n493), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT31), .ZN(new_n519));
  INV_X1    g333(.A(new_n493), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n480), .B1(new_n507), .B2(new_n484), .ZN(new_n521));
  OAI211_X1 g335(.A(KEYINPUT71), .B(new_n520), .C1(new_n521), .C2(new_n482), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n515), .A2(new_n517), .A3(new_n519), .A4(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(G472), .A2(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT32), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT32), .ZN(new_n528));
  AOI211_X1 g342(.A(KEYINPUT72), .B(new_n528), .C1(new_n523), .C2(new_n524), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n513), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT80), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT22), .B(G137), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n222), .A2(G128), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n535), .A2(KEYINPUT23), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n265), .A2(G119), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n536), .A2(new_n539), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G110), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n535), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT24), .B(G110), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n338), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n301), .B(new_n302), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n544), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT75), .B(G110), .Z(new_n549));
  OAI21_X1  g363(.A(new_n548), .B1(new_n541), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n550), .A3(new_n335), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT77), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n534), .B(new_n546), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n546), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n551), .A2(new_n552), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n552), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n534), .B(KEYINPUT78), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n555), .B(new_n283), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT79), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n392), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(G234), .B2(new_n283), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT25), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n567), .A2(G902), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n555), .B(new_n570), .C1(new_n559), .C2(new_n560), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n530), .A2(new_n531), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n531), .B1(new_n530), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n465), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  AOI21_X1  g392(.A(new_n466), .B1(new_n523), .B2(new_n283), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n580), .A2(new_n525), .A3(new_n464), .ZN(new_n581));
  INV_X1    g395(.A(new_n287), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n286), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n294), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n296), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n581), .A2(new_n573), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n357), .A2(new_n360), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n192), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n391), .A2(new_n394), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n398), .B1(new_n397), .B2(new_n381), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT33), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n395), .A2(new_n399), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(G478), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(G478), .A2(G902), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n400), .A2(new_n402), .A3(new_n283), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n589), .A2(new_n590), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n587), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT34), .B(G104), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n404), .A2(new_n405), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n350), .A2(new_n356), .A3(KEYINPUT94), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n349), .A2(new_n608), .A3(KEYINPUT20), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n606), .A2(new_n607), .A3(new_n360), .A4(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n605), .B1(new_n610), .B2(new_n590), .ZN(new_n611));
  INV_X1    g425(.A(new_n610), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(KEYINPUT95), .A3(new_n192), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n587), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT35), .B(G107), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  INV_X1    g430(.A(KEYINPUT36), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n560), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n559), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n570), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n569), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n622), .A2(new_n406), .A3(new_n590), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n581), .A2(new_n298), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT37), .B(G110), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G12));
  NAND4_X1  g440(.A1(new_n530), .A2(new_n464), .A3(new_n586), .A4(new_n621), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n189), .B(KEYINPUT96), .ZN(new_n628));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  INV_X1    g443(.A(new_n191), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n610), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n265), .ZN(G30));
  INV_X1    g449(.A(new_n524), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n489), .A2(new_n514), .A3(new_n493), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n483), .B1(new_n503), .B2(new_n504), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n481), .B1(new_n638), .B2(new_n480), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT71), .B1(new_n639), .B2(new_n520), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n517), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n516), .B1(new_n505), .B2(new_n493), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n636), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n528), .B1(new_n645), .B2(KEYINPUT72), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT32), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n283), .B1(new_n508), .B2(new_n493), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n505), .A2(new_n520), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n648), .A2(KEYINPUT97), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT97), .B1(new_n648), .B2(new_n651), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n631), .B(KEYINPUT39), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n464), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n295), .B(KEYINPUT38), .Z(new_n662));
  AOI22_X1  g476(.A1(new_n357), .A2(new_n360), .B1(new_n404), .B2(new_n405), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n296), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n621), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n656), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(new_n238), .ZN(G45));
  AND3_X1   g483(.A1(new_n530), .A2(new_n464), .A3(new_n586), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n589), .A2(new_n599), .A3(new_n631), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n670), .A2(new_n671), .A3(new_n621), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n672), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT99), .B1(new_n627), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  INV_X1    g491(.A(new_n455), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n447), .ZN(new_n679));
  OAI21_X1  g493(.A(G469), .B1(new_n679), .B2(G902), .ZN(new_n680));
  INV_X1    g494(.A(new_n409), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n410), .B(new_n283), .C1(new_n678), .C2(new_n447), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n585), .A2(new_n683), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n530), .A2(new_n573), .A3(new_n684), .A4(new_n600), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT100), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G15));
  NAND2_X1  g502(.A1(new_n613), .A2(new_n611), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n530), .A3(new_n573), .A4(new_n684), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  NAND3_X1  g505(.A1(new_n530), .A2(new_n623), .A3(new_n684), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  OR2_X1    g507(.A1(new_n509), .A2(new_n493), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n636), .B1(new_n694), .B2(new_n644), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n579), .A2(new_n683), .A3(new_n572), .A4(new_n695), .ZN(new_n696));
  AND4_X1   g510(.A1(new_n192), .A2(new_n584), .A3(new_n663), .A4(new_n296), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n683), .ZN(new_n700));
  INV_X1    g514(.A(new_n695), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n580), .A2(new_n700), .A3(new_n573), .A4(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n584), .A2(new_n663), .A3(new_n192), .A4(new_n296), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT101), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NOR3_X1   g520(.A1(new_n622), .A2(new_n579), .A3(new_n695), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n684), .A2(new_n672), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  XNOR2_X1  g523(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n409), .A2(new_n666), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n463), .A2(KEYINPUT102), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n459), .A2(new_n444), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n460), .A2(new_n461), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .A4(G469), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n457), .A2(new_n713), .A3(KEYINPUT103), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  INV_X1    g533(.A(new_n411), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n682), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n716), .B1(new_n462), .B2(G469), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n712), .B(new_n295), .C1(new_n718), .C2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n530), .A3(new_n573), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n710), .B1(new_n725), .B2(new_n674), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT32), .B1(new_n523), .B2(new_n524), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n512), .B1(new_n727), .B2(KEYINPUT105), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n645), .B2(KEYINPUT32), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n645), .A2(KEYINPUT32), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n589), .A2(new_n599), .A3(new_n733), .A4(new_n631), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n724), .A2(new_n732), .A3(new_n573), .A4(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(KEYINPUT106), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(KEYINPUT106), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n726), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  AND2_X1   g553(.A1(new_n632), .A2(KEYINPUT107), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n632), .A2(KEYINPUT107), .ZN(new_n741));
  OR3_X1    g555(.A1(new_n725), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  NOR2_X1   g557(.A1(new_n588), .A2(new_n599), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(KEYINPUT43), .Z(new_n745));
  OAI21_X1  g559(.A(new_n621), .B1(new_n579), .B2(new_n645), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT108), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n295), .A2(new_n666), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n462), .B(KEYINPUT45), .Z(new_n756));
  OAI211_X1 g570(.A(new_n755), .B(G469), .C1(new_n756), .C2(G902), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(G469), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(KEYINPUT46), .A3(new_n720), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n682), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n681), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n657), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n750), .A2(new_n754), .A3(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT109), .B(G137), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G39));
  NAND2_X1  g579(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n760), .B2(new_n681), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n761), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(new_n766), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n512), .B1(new_n646), .B2(new_n647), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n674), .A2(new_n753), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n572), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  INV_X1    g587(.A(new_n628), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n752), .A2(new_n700), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n745), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n732), .A2(new_n573), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT115), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(KEYINPUT48), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n782), .A2(KEYINPUT48), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n188), .A2(G952), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n655), .A2(new_n573), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n189), .A3(new_n775), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n589), .A2(new_n599), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n783), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n580), .A2(new_n573), .A3(new_n701), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n745), .A2(new_n774), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n684), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n708), .B1(new_n627), .B2(new_n633), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n631), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n622), .A2(KEYINPUT112), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n621), .B2(new_n631), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n585), .A2(new_n664), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n718), .A2(new_n723), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n681), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n804), .B1(new_n653), .B2(new_n654), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n530), .A2(new_n464), .A3(new_n586), .A4(new_n621), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n671), .B1(new_n806), .B2(new_n672), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n627), .A2(KEYINPUT99), .A3(new_n674), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n796), .B(new_n805), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n795), .B1(new_n673), .B2(new_n675), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(KEYINPUT52), .A3(new_n805), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n724), .A2(new_n672), .A3(new_n707), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n607), .A2(new_n360), .A3(new_n609), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n753), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n622), .A2(new_n606), .A3(new_n631), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n530), .A3(new_n464), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n530), .A2(new_n464), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(KEYINPUT111), .A3(new_n817), .A4(new_n818), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n815), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n738), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT80), .B1(new_n770), .B2(new_n572), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n574), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n685), .B1(new_n827), .B2(new_n465), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n588), .A2(new_n599), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n192), .A3(new_n406), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n297), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n573), .A3(new_n581), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n692), .A3(new_n624), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n702), .A2(new_n703), .A3(KEYINPUT101), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n828), .A2(new_n837), .A3(new_n690), .A4(new_n742), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n825), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n814), .A2(new_n839), .A3(KEYINPUT53), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT53), .B1(new_n814), .B2(new_n839), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT54), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  AND4_X1   g658(.A1(KEYINPUT52), .A2(new_n676), .A3(new_n796), .A4(new_n805), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(new_n812), .B2(new_n805), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n685), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n577), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n692), .A2(new_n624), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n690), .A3(new_n705), .A4(new_n832), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n738), .A3(new_n742), .A4(new_n824), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n844), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n814), .A2(new_n839), .A3(KEYINPUT53), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n843), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n794), .B1(new_n842), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT51), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n787), .A2(new_n589), .A3(new_n599), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n776), .A2(new_n707), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n680), .A2(new_n682), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n681), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n752), .B(new_n792), .C1(new_n769), .C2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n792), .A2(new_n666), .A3(new_n662), .A4(new_n700), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT50), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n859), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n858), .A2(KEYINPUT51), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT54), .B1(new_n840), .B2(new_n841), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n854), .A2(new_n843), .A3(new_n855), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT113), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n793), .A2(new_n857), .A3(new_n870), .A4(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(G952), .B2(G953), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n862), .B(KEYINPUT49), .Z(new_n876));
  NAND3_X1  g690(.A1(new_n662), .A2(new_n744), .A3(new_n876), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n786), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n712), .B2(new_n878), .ZN(G75));
  NOR2_X1   g693(.A1(new_n188), .A2(G952), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n291), .B(new_n270), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n840), .A2(new_n841), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n283), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(G210), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n854), .A2(new_n855), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(G902), .A3(new_n289), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n882), .A2(new_n886), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n888), .A2(KEYINPUT117), .A3(G902), .A4(new_n289), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n891), .A2(KEYINPUT118), .A3(new_n892), .A4(new_n893), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n880), .B(new_n887), .C1(new_n896), .C2(new_n897), .ZN(G51));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n872), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n854), .A2(KEYINPUT119), .A3(new_n843), .A4(new_n855), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n871), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n411), .B(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n679), .B(KEYINPUT120), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n884), .A2(G469), .A3(new_n756), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n880), .B1(new_n906), .B2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  INV_X1    g723(.A(new_n354), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n911), .A2(new_n912), .A3(new_n880), .ZN(G60));
  NAND2_X1  g727(.A1(new_n593), .A2(new_n595), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n597), .B(KEYINPUT59), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n902), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n880), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT121), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n920), .B(new_n880), .C1(new_n902), .C2(new_n916), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n857), .A2(new_n873), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n914), .B1(new_n922), .B2(new_n915), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n919), .A2(new_n921), .A3(new_n923), .ZN(G63));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT60), .Z(new_n926));
  NAND3_X1  g740(.A1(new_n888), .A2(new_n619), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n888), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n555), .B1(new_n559), .B2(new_n560), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n888), .A2(new_n932), .A3(new_n619), .A4(new_n926), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n928), .A2(new_n931), .A3(new_n918), .A4(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g749(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G66));
  NAND2_X1  g753(.A1(new_n190), .A2(G224), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n852), .B2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n237), .B1(G898), .B2(new_n188), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  AND2_X1   g758(.A1(new_n829), .A2(new_n406), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n659), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n827), .A2(new_n752), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n763), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n668), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n812), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n772), .A3(new_n955), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n345), .B(KEYINPUT124), .Z(new_n957));
  XNOR2_X1  g771(.A(new_n501), .B(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n188), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(G227), .ZN(new_n961));
  OAI21_X1  g775(.A(G953), .B1(new_n961), .B2(new_n629), .ZN(new_n962));
  NAND2_X1  g776(.A1(G900), .A2(G953), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n762), .A2(new_n802), .A3(new_n777), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n763), .A2(new_n772), .A3(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n965), .A2(new_n738), .A3(new_n742), .A4(new_n812), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n963), .B1(new_n966), .B2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n958), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n960), .A2(new_n962), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(new_n960), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G72));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT63), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n505), .A2(new_n520), .ZN(new_n974));
  OR4_X1    g788(.A1(new_n650), .A2(new_n883), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n973), .B(KEYINPUT127), .Z(new_n976));
  INV_X1    g790(.A(new_n852), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n966), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n974), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n975), .A2(new_n979), .A3(new_n918), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n976), .B1(new_n956), .B2(new_n977), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n650), .B2(new_n981), .ZN(G57));
endmodule


