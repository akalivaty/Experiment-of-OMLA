//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n197), .A3(new_n200), .A4(new_n195), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT81), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(KEYINPUT81), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n205), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n211), .A2(G107), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n209), .A2(new_n210), .A3(new_n212), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n212), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT66), .A3(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT65), .A2(G146), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT65), .A2(G146), .ZN(new_n227));
  OAI21_X1  g041(.A(G143), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n225), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT1), .B1(new_n223), .B2(G146), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n225), .A2(new_n228), .B1(G128), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n217), .B(new_n219), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(KEYINPUT82), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT82), .B1(new_n234), .B2(new_n235), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT65), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT65), .A2(G146), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n223), .A3(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT64), .B1(new_n223), .B2(G146), .ZN(new_n243));
  OR3_X1    g057(.A1(new_n223), .A2(KEYINPUT64), .A3(G146), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT65), .B(G146), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n249), .A2(G143), .B1(new_n222), .B2(new_n224), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT0), .A3(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n214), .B1(new_n215), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n212), .B1(new_n205), .B2(new_n208), .ZN(new_n256));
  OAI21_X1  g070(.A(G101), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n259), .B(G101), .C1(new_n255), .C2(new_n256), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n217), .A2(new_n219), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT83), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n217), .A2(new_n264), .A3(new_n219), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n249), .B2(G143), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n245), .B1(new_n268), .B2(new_n229), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n250), .A2(new_n230), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n235), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n253), .A2(new_n261), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n203), .B1(new_n239), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n231), .A2(new_n233), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n235), .B1(new_n274), .B2(new_n262), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n236), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n258), .A2(new_n251), .A3(new_n248), .A4(new_n260), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n217), .A2(new_n264), .A3(new_n219), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n264), .B1(new_n217), .B2(new_n219), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n269), .A2(new_n270), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT10), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n279), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n278), .A2(new_n285), .A3(new_n202), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n191), .B1(new_n273), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT85), .ZN(new_n288));
  INV_X1    g102(.A(new_n262), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n234), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n202), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT12), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT12), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n293), .A3(new_n202), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n271), .B1(new_n281), .B2(new_n280), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n277), .A2(new_n295), .A3(new_n279), .A4(new_n236), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n292), .B(new_n294), .C1(new_n296), .C2(new_n202), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n297), .A2(new_n191), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n299), .B(new_n191), .C1(new_n273), .C2(new_n286), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n288), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G469), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(G469), .A2(G902), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n191), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n239), .A2(new_n272), .A3(new_n203), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n296), .A2(new_n202), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n190), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n306), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n307), .B1(new_n306), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g126(.A(G469), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n304), .A2(new_n305), .A3(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT9), .B(G234), .Z(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G221), .B1(new_n316), .B2(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT86), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n320), .A3(new_n317), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G217), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(G234), .B2(new_n303), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n331), .B2(new_n325), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n221), .ZN(new_n333));
  OAI211_X1 g147(.A(G146), .B(new_n327), .C1(new_n331), .C2(new_n325), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(KEYINPUT75), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n336), .A3(new_n221), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n229), .A2(KEYINPUT74), .A3(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n229), .A2(G119), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT74), .B1(new_n229), .B2(G119), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT24), .B(G110), .Z(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n229), .A2(KEYINPUT23), .A3(G119), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n345), .B(new_n346), .C1(G119), .C2(new_n229), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G110), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n335), .A2(new_n337), .A3(new_n343), .A4(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT76), .B(G110), .ZN(new_n350));
  OAI22_X1  g164(.A1(new_n347), .A2(new_n350), .B1(new_n341), .B2(new_n342), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n249), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT77), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n249), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n351), .A2(new_n334), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT79), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n349), .A2(new_n361), .A3(new_n358), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT78), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n364), .A2(KEYINPUT22), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(KEYINPUT22), .ZN(new_n366));
  OR3_X1    g180(.A1(new_n365), .A2(new_n366), .A3(new_n196), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n196), .B1(new_n365), .B2(new_n366), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n359), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(new_n361), .A3(new_n367), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT25), .B1(new_n373), .B2(new_n303), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n375));
  AOI211_X1 g189(.A(new_n375), .B(G902), .C1(new_n370), .C2(new_n372), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n324), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n324), .A2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n377), .A2(KEYINPUT80), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT80), .B1(new_n377), .B2(new_n379), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n248), .A2(new_n251), .A3(new_n202), .ZN(new_n384));
  INV_X1    g198(.A(new_n195), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n193), .A2(G137), .ZN(new_n386));
  OAI21_X1  g200(.A(G131), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n201), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n269), .B2(new_n270), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n383), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT2), .A2(G113), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n393));
  INV_X1    g207(.A(G113), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT67), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT67), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(KEYINPUT2), .B2(G113), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n392), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G116), .B(G119), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT68), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n248), .A2(new_n251), .A3(new_n202), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G128), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n231), .B1(new_n245), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n403), .B(KEYINPUT30), .C1(new_n406), .C2(new_n388), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n390), .A2(new_n402), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n388), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n283), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n395), .A2(new_n397), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n391), .ZN(new_n412));
  INV_X1    g226(.A(new_n399), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n400), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(KEYINPUT68), .A3(new_n413), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n410), .A2(new_n403), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(G237), .A2(G953), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G210), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT70), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT26), .B(G101), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT29), .B1(new_n419), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n402), .B1(new_n384), .B2(new_n389), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n431), .A2(new_n418), .A3(KEYINPUT71), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT28), .B1(new_n431), .B2(KEYINPUT71), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(new_n426), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n428), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n435), .B1(new_n428), .B2(new_n434), .ZN(new_n437));
  INV_X1    g251(.A(new_n418), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n417), .B1(new_n410), .B2(new_n403), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT28), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n430), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n426), .A2(KEYINPUT29), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n303), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n436), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G472), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT73), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n428), .A2(new_n434), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT72), .ZN(new_n448));
  INV_X1    g262(.A(new_n443), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n428), .A2(new_n434), .A3(new_n435), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT73), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(G472), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT31), .B1(new_n419), .B2(new_n427), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT31), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n408), .A2(new_n426), .A3(new_n456), .A4(new_n418), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT71), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n429), .B1(new_n439), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n431), .A2(new_n418), .A3(KEYINPUT71), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n459), .A2(new_n460), .B1(new_n429), .B2(new_n418), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n455), .B(new_n457), .C1(new_n461), .C2(new_n426), .ZN(new_n462));
  NOR2_X1   g276(.A1(G472), .A2(G902), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT32), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(KEYINPUT32), .A3(new_n463), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n382), .B1(new_n454), .B2(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(G110), .B(G122), .Z(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT87), .B(KEYINPUT5), .ZN(new_n471));
  INV_X1    g285(.A(G119), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G116), .ZN(new_n473));
  OAI21_X1  g287(.A(G113), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G116), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G119), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT87), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT5), .ZN(new_n480));
  AND4_X1   g294(.A1(new_n473), .A2(new_n476), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT88), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n480), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(G116), .A3(new_n472), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n399), .A2(new_n471), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(G113), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n398), .A2(new_n399), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n263), .B2(new_n265), .ZN(new_n490));
  AND4_X1   g304(.A1(new_n416), .A2(new_n258), .A3(new_n415), .A4(new_n260), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n470), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n470), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n258), .A2(new_n415), .A3(new_n416), .A4(new_n260), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n493), .B(new_n494), .C1(new_n282), .C2(new_n489), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n406), .A2(new_n329), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n252), .A2(G125), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G224), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(G953), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n499), .B(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n470), .C1(new_n490), .C2(new_n491), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n496), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT89), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n496), .A2(new_n502), .A3(new_n507), .A4(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n499), .B1(new_n510), .B2(new_n501), .ZN(new_n511));
  INV_X1    g325(.A(new_n501), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT7), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n474), .B1(KEYINPUT5), .B2(new_n399), .ZN(new_n514));
  INV_X1    g328(.A(new_n488), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n514), .A2(new_n262), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n262), .B2(new_n489), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT90), .B(KEYINPUT8), .Z(new_n518));
  XNOR2_X1  g332(.A(new_n470), .B(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n511), .B(new_n513), .C1(new_n517), .C2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n495), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G210), .B1(G237), .B2(G902), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n509), .A2(new_n303), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  AOI211_X1 g339(.A(G902), .B(new_n522), .C1(new_n506), .C2(new_n508), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n524), .B(KEYINPUT91), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n188), .A2(G952), .ZN(new_n529));
  NAND2_X1  g343(.A1(G234), .A2(G237), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT21), .B(G898), .Z(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(G902), .A3(G953), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G214), .B1(G237), .B2(G902), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n528), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n335), .A2(new_n337), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n420), .A2(G143), .A3(G214), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G143), .B1(new_n420), .B2(G214), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n540), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n200), .A3(new_n538), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n541), .A2(new_n544), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n541), .A2(new_n543), .A3(KEYINPUT93), .A4(new_n544), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n537), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n354), .A2(new_n356), .B1(G146), .B2(new_n331), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n540), .B(new_n539), .C1(KEYINPUT18), .C2(G131), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n541), .A2(new_n553), .ZN(new_n554));
  OR3_X1    g368(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G113), .B(G122), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(new_n211), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n550), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n557), .B1(new_n550), .B2(new_n555), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n303), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G475), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT20), .ZN(new_n563));
  INV_X1    g377(.A(new_n557), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n331), .B(KEYINPUT19), .ZN(new_n566));
  INV_X1    g380(.A(new_n249), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n334), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n541), .A2(new_n543), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n564), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n558), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G475), .ZN(new_n573));
  AND4_X1   g387(.A1(new_n563), .A2(new_n572), .A3(new_n573), .A4(new_n303), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(G475), .B1(new_n558), .B2(new_n571), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(new_n303), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n562), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(new_n562), .C1(new_n574), .C2(new_n578), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n229), .A2(G143), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT96), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n229), .A2(G143), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n193), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(G116), .B(G122), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(new_n207), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n591), .A2(new_n586), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n586), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n595), .A3(new_n586), .ZN(new_n596));
  AND4_X1   g410(.A1(new_n592), .A2(new_n594), .A3(new_n596), .A4(new_n585), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n588), .B(new_n590), .C1(new_n597), .C2(new_n193), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n585), .A2(new_n587), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G134), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n588), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n475), .A2(G122), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n207), .B1(new_n602), .B2(KEYINPUT14), .ZN(new_n603));
  INV_X1    g417(.A(new_n589), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n316), .A2(new_n323), .A3(G953), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n598), .A2(new_n607), .A3(new_n609), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(KEYINPUT15), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n613), .B(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n583), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n322), .A2(new_n469), .A3(new_n536), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  OR2_X1    g434(.A1(new_n380), .A2(new_n381), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n462), .A2(new_n303), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n623), .A2(new_n464), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n314), .A2(new_n320), .A3(new_n317), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n320), .B1(new_n314), .B2(new_n317), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n621), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n535), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n509), .A2(new_n303), .A3(new_n523), .ZN(new_n629));
  INV_X1    g443(.A(new_n524), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n628), .B1(new_n631), .B2(new_n525), .ZN(new_n632));
  INV_X1    g446(.A(new_n613), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT98), .A3(new_n614), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n613), .B2(G478), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n611), .A2(KEYINPUT33), .A3(new_n612), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT33), .B1(new_n611), .B2(new_n612), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n614), .A2(G902), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n634), .A2(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n580), .B2(new_n582), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n632), .A2(new_n534), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n627), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  AND3_X1   g460(.A1(new_n577), .A2(new_n303), .A3(new_n576), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n578), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(KEYINPUT99), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n649), .A2(new_n650), .B1(G475), .B2(new_n561), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n632), .A2(new_n534), .A3(new_n617), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n627), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  OAI211_X1 g469(.A(new_n536), .B(new_n618), .C1(new_n625), .C2(new_n626), .ZN(new_n656));
  INV_X1    g470(.A(new_n624), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT36), .B1(new_n367), .B2(new_n368), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n359), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n378), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n377), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n656), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT37), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G110), .ZN(G12));
  OAI21_X1  g479(.A(new_n531), .B1(G900), .B2(new_n533), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT100), .Z(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n651), .A2(new_n617), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n662), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n451), .A2(new_n452), .A3(G472), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n452), .B1(new_n451), .B2(G472), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n468), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n322), .A2(new_n670), .A3(new_n673), .A4(new_n632), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XOR2_X1   g489(.A(new_n667), .B(KEYINPUT39), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n322), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n528), .B(KEYINPUT38), .Z(new_n679));
  INV_X1    g493(.A(new_n419), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n427), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n438), .A2(new_n439), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n303), .B1(new_n683), .B2(new_n426), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n466), .A2(new_n467), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n583), .A2(new_n617), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n679), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n661), .A2(new_n628), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n322), .A2(new_n691), .A3(new_n676), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n678), .A2(new_n689), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  NAND2_X1  g508(.A1(new_n642), .A2(new_n668), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n662), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n322), .A2(new_n673), .A3(new_n632), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  AND3_X1   g512(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n302), .B1(new_n301), .B2(new_n303), .ZN(new_n700));
  INV_X1    g514(.A(new_n317), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n673), .A2(new_n621), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n643), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT41), .B(G113), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT101), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n704), .B(new_n706), .ZN(G15));
  NOR2_X1   g521(.A1(new_n703), .A2(new_n652), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n475), .ZN(G18));
  NAND2_X1  g523(.A1(new_n301), .A2(new_n303), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n317), .A3(new_n304), .ZN(new_n712));
  INV_X1    g526(.A(new_n525), .ZN(new_n713));
  AOI21_X1  g527(.A(G902), .B1(new_n506), .B2(new_n508), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n524), .B1(new_n714), .B2(new_n523), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n535), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n712), .A2(new_n716), .A3(new_n662), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n466), .A2(new_n467), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n446), .B2(new_n453), .ZN(new_n719));
  INV_X1    g533(.A(new_n583), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n534), .A3(new_n616), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND3_X1  g538(.A1(new_n702), .A2(new_n534), .A3(new_n632), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n441), .A2(new_n427), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n455), .A3(new_n457), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n463), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n623), .A2(new_n377), .A3(new_n379), .A4(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT102), .B1(new_n583), .B2(new_n617), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n732), .B(new_n616), .C1(new_n580), .C2(new_n582), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n730), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n725), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(G122), .Z(G24));
  INV_X1    g550(.A(new_n695), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n623), .A2(new_n661), .A3(new_n728), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n702), .A3(new_n632), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  NAND2_X1  g554(.A1(new_n377), .A2(new_n379), .ZN(new_n741));
  AOI22_X1  g555(.A1(KEYINPUT106), .A2(new_n468), .B1(new_n446), .B2(new_n453), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n468), .A2(KEYINPUT106), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n310), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT104), .A4(new_n190), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT103), .B1(new_n297), .B2(new_n191), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n297), .A2(KEYINPUT103), .A3(new_n191), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n748), .B(G469), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n304), .A2(new_n305), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n317), .ZN(new_n753));
  INV_X1    g567(.A(new_n527), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n629), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n525), .A3(new_n535), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n753), .A2(new_n695), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n753), .A2(new_n756), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n469), .A2(new_n759), .A3(new_n737), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n758), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  OR2_X1    g580(.A1(new_n669), .A2(KEYINPUT107), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n669), .A2(KEYINPUT107), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n469), .A3(new_n759), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NOR2_X1   g584(.A1(new_n583), .A2(new_n641), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT43), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n583), .B2(new_n641), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n657), .A3(new_n661), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n756), .ZN(new_n779));
  OR3_X1    g593(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT45), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n748), .B(KEYINPUT45), .C1(new_n749), .C2(new_n750), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(G469), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n305), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n305), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n304), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n317), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n776), .A2(new_n777), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n779), .A2(new_n789), .A3(new_n676), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  OR2_X1    g606(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n673), .A2(new_n621), .A3(new_n756), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n793), .A2(new_n737), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n753), .A2(new_n687), .A3(new_n661), .A4(new_n667), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n688), .A2(new_n732), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n583), .A2(KEYINPUT102), .A3(new_n617), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n716), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n674), .A2(new_n697), .A3(new_n739), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(KEYINPUT111), .A3(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT111), .B(KEYINPUT112), .Z(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n719), .B1(new_n319), .B2(new_n321), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n809), .B(new_n632), .C1(new_n670), .C2(new_n696), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(KEYINPUT52), .A3(new_n739), .A4(new_n803), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n806), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n808), .B1(new_n806), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n469), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n528), .A2(new_n642), .A3(new_n534), .A4(new_n535), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT108), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n628), .B1(new_n755), .B2(new_n525), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT108), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n819), .A3(new_n534), .A4(new_n642), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  OAI22_X1  g635(.A1(new_n815), .A2(new_n656), .B1(new_n627), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n663), .B1(new_n822), .B2(KEYINPUT109), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n673), .A2(new_n534), .A3(new_n618), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n702), .A2(new_n632), .A3(new_n661), .ZN(new_n825));
  OAI22_X1  g639(.A1(new_n703), .A2(new_n652), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI22_X1  g640(.A1(new_n703), .A2(new_n643), .B1(new_n725), .B2(new_n734), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n627), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n616), .B(KEYINPUT110), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n536), .A3(new_n720), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT109), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n619), .B(new_n832), .C1(new_n627), .C2(new_n821), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n823), .A2(new_n828), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n651), .A2(new_n668), .ZN(new_n835));
  INV_X1    g649(.A(new_n756), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n662), .A2(new_n830), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n809), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n757), .A2(new_n738), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n769), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n765), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n834), .A2(new_n842), .A3(KEYINPUT53), .ZN(new_n843));
  INV_X1    g657(.A(new_n663), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n822), .A2(KEYINPUT109), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n844), .A2(new_n845), .A3(new_n831), .A4(new_n833), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n804), .A2(new_n805), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n811), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n760), .A2(new_n762), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT105), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n840), .B1(new_n852), .B2(new_n758), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n846), .A2(new_n828), .A3(new_n848), .A4(new_n853), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n814), .A2(new_n843), .B1(new_n854), .B2(KEYINPUT53), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n798), .B1(new_n855), .B2(KEYINPUT54), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n834), .A2(new_n842), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n806), .A2(new_n811), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n807), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n806), .A2(new_n808), .A3(new_n811), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n857), .A2(new_n858), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n854), .A2(KEYINPUT53), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n798), .A2(new_n862), .A3(new_n863), .A4(KEYINPUT54), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n856), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n719), .A2(new_n382), .A3(new_n712), .ZN(new_n867));
  INV_X1    g681(.A(new_n643), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n702), .A2(new_n534), .A3(new_n632), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n729), .B1(new_n800), .B2(new_n801), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n867), .A2(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n652), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n867), .A2(new_n872), .B1(new_n717), .B2(new_n722), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT114), .B1(new_n826), .B2(new_n827), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n765), .A3(KEYINPUT115), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n841), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT115), .B1(new_n877), .B2(new_n765), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n823), .A2(new_n831), .A3(new_n833), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n858), .B1(new_n882), .B2(new_n814), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n857), .A2(new_n858), .A3(new_n848), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n866), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n531), .B1(new_n772), .B2(new_n774), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n712), .A2(new_n756), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n744), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT48), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n686), .A2(new_n531), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n621), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n642), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n529), .A3(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n887), .A2(new_n730), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n793), .A2(new_n795), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n711), .A2(new_n304), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n317), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n836), .B(new_n897), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n628), .A3(new_n702), .ZN(new_n903));
  INV_X1    g717(.A(new_n679), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n903), .A2(KEYINPUT50), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT50), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n894), .A2(new_n720), .A3(new_n641), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT51), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n889), .A2(new_n738), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n902), .A2(new_n912), .A3(new_n908), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n911), .ZN(new_n915));
  NAND2_X1  g729(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n896), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n865), .A2(new_n886), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n897), .A2(new_n632), .A3(new_n702), .ZN(new_n920));
  OAI22_X1  g734(.A1(new_n919), .A2(new_n920), .B1(G952), .B2(G953), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n900), .A2(KEYINPUT49), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n900), .A2(KEYINPUT49), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n741), .A2(new_n701), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n922), .A2(new_n535), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n679), .A2(new_n687), .A3(new_n771), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(G75));
  NOR2_X1   g741(.A1(new_n188), .A2(G952), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n877), .A2(new_n765), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT115), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(new_n846), .A3(new_n878), .A4(new_n841), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n860), .A2(new_n861), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT53), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n884), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(G210), .A3(G902), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n496), .A2(new_n504), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n502), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT55), .Z(new_n941));
  AOI21_X1  g755(.A(new_n928), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n935), .A2(G902), .A3(new_n754), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT117), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n941), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n883), .A2(new_n303), .A3(new_n885), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(KEYINPUT117), .A3(new_n754), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n945), .A2(new_n937), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n942), .A2(new_n949), .ZN(G51));
  NAND3_X1  g764(.A1(new_n934), .A2(KEYINPUT54), .A3(new_n884), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n886), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n305), .B(KEYINPUT57), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n301), .ZN(new_n955));
  INV_X1    g769(.A(new_n782), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n934), .A2(G902), .A3(new_n956), .A4(new_n884), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT118), .Z(new_n958));
  AOI21_X1  g772(.A(new_n928), .B1(new_n955), .B2(new_n958), .ZN(G54));
  NAND2_X1  g773(.A1(KEYINPUT58), .A2(G475), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT119), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n960), .A2(KEYINPUT119), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n947), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n571), .A3(new_n558), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n947), .A2(new_n572), .A3(new_n961), .A4(new_n962), .ZN(new_n965));
  INV_X1    g779(.A(new_n928), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G60));
  NAND2_X1  g781(.A1(G478), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT59), .Z(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n865), .B2(new_n886), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n966), .B1(new_n970), .B2(new_n639), .ZN(new_n971));
  INV_X1    g785(.A(new_n969), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n934), .A2(KEYINPUT54), .A3(new_n884), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT54), .B1(new_n934), .B2(new_n884), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n639), .B(new_n972), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT120), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n952), .A2(KEYINPUT120), .A3(new_n639), .A4(new_n972), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n971), .A2(new_n979), .ZN(G63));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT60), .Z(new_n982));
  NAND2_X1  g796(.A1(new_n935), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n373), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n935), .A2(new_n659), .A3(new_n982), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n966), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n985), .A2(KEYINPUT61), .A3(new_n966), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G66));
  NAND2_X1  g805(.A1(new_n834), .A2(new_n188), .ZN(new_n992));
  INV_X1    g806(.A(new_n532), .ZN(new_n993));
  OAI21_X1  g807(.A(G953), .B1(new_n993), .B2(new_n500), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(KEYINPUT121), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(KEYINPUT121), .B2(new_n992), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n939), .B1(G898), .B2(new_n188), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n996), .B(new_n997), .Z(G69));
  AND2_X1   g812(.A1(new_n390), .A2(new_n407), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(new_n566), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n674), .A2(new_n697), .A3(new_n739), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n693), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n642), .B1(new_n720), .B2(new_n830), .ZN(new_n1005));
  OR4_X1    g819(.A1(new_n815), .A2(new_n677), .A3(new_n756), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n796), .A2(new_n791), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1000), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n765), .A2(new_n769), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT123), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n789), .A2(new_n676), .A3(new_n744), .A4(new_n802), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1012), .A2(new_n1001), .A3(new_n1007), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1000), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1014), .A2(new_n188), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT122), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n188), .A2(G900), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1010), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(G72));
  INV_X1    g835(.A(KEYINPUT127), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1014), .B2(new_n834), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1025), .A2(new_n427), .A3(new_n680), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1024), .B1(new_n1008), .B2(new_n834), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT124), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1027), .A2(new_n1028), .A3(new_n681), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1028), .B1(new_n1027), .B2(new_n681), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1026), .B(new_n966), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n855), .ZN(new_n1033));
  OAI21_X1  g847(.A(KEYINPUT125), .B1(new_n419), .B2(new_n427), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n419), .A2(new_n427), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n1024), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT126), .Z(new_n1038));
  NOR2_X1   g852(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1022), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1027), .A2(new_n681), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(KEYINPUT124), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n928), .B1(new_n1042), .B2(new_n1029), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1039), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1043), .A2(KEYINPUT127), .A3(new_n1026), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1040), .A2(new_n1045), .ZN(G57));
endmodule


