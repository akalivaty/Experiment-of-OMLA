

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U546 ( .A1(n744), .A2(n997), .ZN(n746) );
  AND2_X1 U547 ( .A1(n989), .A2(n814), .ZN(n511) );
  INV_X1 U548 ( .A(n765), .ZN(n745) );
  NOR2_X1 U549 ( .A1(G651), .A2(G543), .ZN(n638) );
  NOR2_X1 U550 ( .A1(n800), .A2(n511), .ZN(n801) );
  XOR2_X1 U551 ( .A(KEYINPUT1), .B(n531), .Z(n639) );
  NOR2_X1 U552 ( .A1(n522), .A2(n521), .ZN(G160) );
  INV_X1 U553 ( .A(G2105), .ZN(n513) );
  NOR2_X4 U554 ( .A1(G2104), .A2(n513), .ZN(n887) );
  NAND2_X1 U555 ( .A1(G125), .A2(n887), .ZN(n512) );
  XNOR2_X1 U556 ( .A(n512), .B(KEYINPUT64), .ZN(n516) );
  AND2_X4 U557 ( .A1(n513), .A2(G2104), .ZN(n883) );
  NAND2_X1 U558 ( .A1(G101), .A2(n883), .ZN(n514) );
  XOR2_X1 U559 ( .A(KEYINPUT23), .B(n514), .Z(n515) );
  NAND2_X1 U560 ( .A1(n516), .A2(n515), .ZN(n522) );
  NAND2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XNOR2_X1 U562 ( .A(n517), .B(KEYINPUT65), .ZN(n888) );
  NAND2_X1 U563 ( .A1(G113), .A2(n888), .ZN(n520) );
  NOR2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n518), .Z(n884) );
  NAND2_X1 U566 ( .A1(G137), .A2(n884), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U568 ( .A1(G138), .A2(n884), .ZN(n523) );
  XNOR2_X1 U569 ( .A(n523), .B(KEYINPUT90), .ZN(n529) );
  AND2_X1 U570 ( .A1(n888), .A2(G114), .ZN(n527) );
  NAND2_X1 U571 ( .A1(G102), .A2(n883), .ZN(n525) );
  NAND2_X1 U572 ( .A1(G126), .A2(n887), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n528) );
  AND2_X1 U575 ( .A1(n529), .A2(n528), .ZN(G164) );
  INV_X1 U576 ( .A(G57), .ZN(G237) );
  INV_X1 U577 ( .A(G132), .ZN(G219) );
  INV_X1 U578 ( .A(G82), .ZN(G220) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n619) );
  NOR2_X2 U580 ( .A1(G651), .A2(n619), .ZN(n637) );
  NAND2_X1 U581 ( .A1(n637), .A2(G52), .ZN(n530) );
  XOR2_X1 U582 ( .A(KEYINPUT67), .B(n530), .Z(n533) );
  INV_X1 U583 ( .A(G651), .ZN(n535) );
  NOR2_X1 U584 ( .A1(G543), .A2(n535), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n639), .A2(G64), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U587 ( .A(KEYINPUT68), .B(n534), .ZN(n540) );
  NAND2_X1 U588 ( .A1(G90), .A2(n638), .ZN(n537) );
  NOR2_X1 U589 ( .A1(n619), .A2(n535), .ZN(n642) );
  NAND2_X1 U590 ( .A1(G77), .A2(n642), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U592 ( .A(KEYINPUT9), .B(n538), .Z(n539) );
  NOR2_X1 U593 ( .A1(n540), .A2(n539), .ZN(G171) );
  NAND2_X1 U594 ( .A1(G89), .A2(n638), .ZN(n541) );
  XNOR2_X1 U595 ( .A(n541), .B(KEYINPUT74), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n542), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G76), .A2(n642), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT5), .ZN(n550) );
  NAND2_X1 U600 ( .A1(G63), .A2(n639), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G51), .A2(n637), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n548), .Z(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U605 ( .A(n551), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U607 ( .A1(G94), .A2(G452), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U609 ( .A1(G7), .A2(G661), .ZN(n553) );
  XOR2_X1 U610 ( .A(n553), .B(KEYINPUT10), .Z(n829) );
  NAND2_X1 U611 ( .A1(n829), .A2(G567), .ZN(n554) );
  XOR2_X1 U612 ( .A(KEYINPUT11), .B(n554), .Z(G234) );
  NAND2_X1 U613 ( .A1(G81), .A2(n638), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT12), .B(n555), .Z(n556) );
  XNOR2_X1 U615 ( .A(n556), .B(KEYINPUT71), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G68), .A2(n642), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U618 ( .A(KEYINPUT13), .B(n559), .ZN(n566) );
  NAND2_X1 U619 ( .A1(G56), .A2(n639), .ZN(n560) );
  XNOR2_X1 U620 ( .A(KEYINPUT14), .B(n560), .ZN(n561) );
  INV_X1 U621 ( .A(n561), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n637), .A2(G43), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT72), .B(n562), .Z(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n992) );
  INV_X1 U626 ( .A(G860), .ZN(n586) );
  OR2_X1 U627 ( .A1(n992), .A2(n586), .ZN(G153) );
  INV_X1 U628 ( .A(G171), .ZN(G301) );
  NAND2_X1 U629 ( .A1(G868), .A2(G301), .ZN(n576) );
  NAND2_X1 U630 ( .A1(G54), .A2(n637), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G79), .A2(n642), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G66), .A2(n639), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G92), .A2(n638), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT73), .B(n569), .ZN(n570) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X2 U638 ( .A(n574), .B(KEYINPUT15), .ZN(n1005) );
  OR2_X1 U639 ( .A1(n1005), .A2(G868), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(G284) );
  NAND2_X1 U641 ( .A1(G91), .A2(n638), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G78), .A2(n642), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(KEYINPUT70), .B(n579), .Z(n583) );
  NAND2_X1 U645 ( .A1(G65), .A2(n639), .ZN(n581) );
  NAND2_X1 U646 ( .A1(G53), .A2(n637), .ZN(n580) );
  AND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(G299) );
  INV_X1 U649 ( .A(G868), .ZN(n658) );
  NOR2_X1 U650 ( .A1(G286), .A2(n658), .ZN(n585) );
  NOR2_X1 U651 ( .A1(G868), .A2(G299), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(G297) );
  NAND2_X1 U653 ( .A1(n586), .A2(G559), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n587), .A2(n1005), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n588), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U656 ( .A1(G559), .A2(n658), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n1005), .A2(n589), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT75), .ZN(n592) );
  NOR2_X1 U659 ( .A1(n992), .A2(G868), .ZN(n591) );
  NOR2_X1 U660 ( .A1(n592), .A2(n591), .ZN(G282) );
  NAND2_X1 U661 ( .A1(G135), .A2(n884), .ZN(n593) );
  XNOR2_X1 U662 ( .A(n593), .B(KEYINPUT76), .ZN(n600) );
  NAND2_X1 U663 ( .A1(G99), .A2(n883), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G111), .A2(n888), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n887), .A2(G123), .ZN(n596) );
  XOR2_X1 U667 ( .A(KEYINPUT18), .B(n596), .Z(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U670 ( .A(KEYINPUT77), .B(n601), .Z(n960) );
  XNOR2_X1 U671 ( .A(G2096), .B(n960), .ZN(n602) );
  NOR2_X1 U672 ( .A1(G2100), .A2(n602), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT78), .B(n603), .Z(G156) );
  NAND2_X1 U674 ( .A1(G559), .A2(n1005), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(n992), .ZN(n655) );
  NOR2_X1 U676 ( .A1(n655), .A2(G860), .ZN(n613) );
  NAND2_X1 U677 ( .A1(n639), .A2(G67), .ZN(n605) );
  XOR2_X1 U678 ( .A(KEYINPUT79), .B(n605), .Z(n607) );
  NAND2_X1 U679 ( .A1(n637), .A2(G55), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U681 ( .A(KEYINPUT80), .B(n608), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G93), .A2(n638), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G80), .A2(n642), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  OR2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n657) );
  XOR2_X1 U686 ( .A(n613), .B(n657), .Z(G145) );
  NAND2_X1 U687 ( .A1(n637), .A2(G49), .ZN(n614) );
  XOR2_X1 U688 ( .A(KEYINPUT81), .B(n614), .Z(n616) );
  NAND2_X1 U689 ( .A1(G651), .A2(G74), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U691 ( .A(KEYINPUT82), .B(n617), .ZN(n618) );
  NOR2_X1 U692 ( .A1(n639), .A2(n618), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n619), .A2(G87), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(G288) );
  NAND2_X1 U695 ( .A1(G60), .A2(n639), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G47), .A2(n637), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G85), .A2(n638), .ZN(n624) );
  XOR2_X1 U699 ( .A(KEYINPUT66), .B(n624), .Z(n625) );
  NOR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n642), .A2(G72), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(G290) );
  NAND2_X1 U703 ( .A1(n637), .A2(G48), .ZN(n635) );
  NAND2_X1 U704 ( .A1(G86), .A2(n638), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G61), .A2(n639), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n642), .A2(G73), .ZN(n631) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n631), .Z(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U711 ( .A(KEYINPUT83), .B(n636), .Z(G305) );
  NAND2_X1 U712 ( .A1(G50), .A2(n637), .ZN(n647) );
  NAND2_X1 U713 ( .A1(G88), .A2(n638), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G62), .A2(n639), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n642), .A2(G75), .ZN(n643) );
  XOR2_X1 U717 ( .A(KEYINPUT84), .B(n643), .Z(n644) );
  NOR2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n648), .B(KEYINPUT85), .ZN(G166) );
  XNOR2_X1 U721 ( .A(KEYINPUT86), .B(G290), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n649), .B(G299), .ZN(n650) );
  XNOR2_X1 U723 ( .A(KEYINPUT19), .B(n650), .ZN(n652) );
  XNOR2_X1 U724 ( .A(G305), .B(G166), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n657), .B(n653), .ZN(n654) );
  XNOR2_X1 U727 ( .A(G288), .B(n654), .ZN(n898) );
  XNOR2_X1 U728 ( .A(n655), .B(n898), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n661) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n662), .ZN(n664) );
  XOR2_X1 U735 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n663) );
  XNOR2_X1 U736 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U737 ( .A1(G2072), .A2(n665), .ZN(G158) );
  XNOR2_X1 U738 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U739 ( .A1(G661), .A2(G483), .ZN(n666) );
  XNOR2_X1 U740 ( .A(KEYINPUT89), .B(n666), .ZN(n675) );
  NOR2_X1 U741 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U742 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U743 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U744 ( .A1(G96), .A2(n669), .ZN(n834) );
  NAND2_X1 U745 ( .A1(G2106), .A2(n834), .ZN(n673) );
  NAND2_X1 U746 ( .A1(G120), .A2(G69), .ZN(n670) );
  NOR2_X1 U747 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U748 ( .A1(G108), .A2(n671), .ZN(n833) );
  NAND2_X1 U749 ( .A1(G567), .A2(n833), .ZN(n672) );
  NAND2_X1 U750 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT88), .B(n674), .Z(n836) );
  AND2_X1 U752 ( .A1(n675), .A2(n836), .ZN(n832) );
  NAND2_X1 U753 ( .A1(n832), .A2(G36), .ZN(G176) );
  XNOR2_X1 U754 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  NOR2_X2 U755 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NAND2_X1 U756 ( .A1(G160), .A2(G40), .ZN(n770) );
  XNOR2_X1 U757 ( .A(n770), .B(KEYINPUT97), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n769), .A2(n676), .ZN(n714) );
  XNOR2_X1 U759 ( .A(G1996), .B(KEYINPUT99), .ZN(n937) );
  NOR2_X1 U760 ( .A1(n714), .A2(n937), .ZN(n680) );
  INV_X1 U761 ( .A(n680), .ZN(n678) );
  XOR2_X1 U762 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n679) );
  INV_X1 U763 ( .A(n679), .ZN(n677) );
  NAND2_X1 U764 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U766 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U767 ( .A1(n714), .A2(G1341), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n684), .A2(n683), .ZN(n692) );
  INV_X1 U769 ( .A(n1005), .ZN(n685) );
  OR2_X1 U770 ( .A1(n685), .A2(n992), .ZN(n686) );
  OR2_X1 U771 ( .A1(n692), .A2(n686), .ZN(n690) );
  INV_X1 U772 ( .A(n714), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n709), .A2(G1348), .ZN(n688) );
  NOR2_X1 U774 ( .A1(G2067), .A2(n714), .ZN(n687) );
  NOR2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U777 ( .A(n691), .B(KEYINPUT101), .ZN(n695) );
  NOR2_X1 U778 ( .A1(n992), .A2(n692), .ZN(n693) );
  NOR2_X1 U779 ( .A1(n1005), .A2(n693), .ZN(n694) );
  NOR2_X1 U780 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U781 ( .A(n696), .B(KEYINPUT102), .ZN(n702) );
  NAND2_X1 U782 ( .A1(n709), .A2(G2072), .ZN(n697) );
  XOR2_X1 U783 ( .A(KEYINPUT27), .B(n697), .Z(n699) );
  INV_X1 U784 ( .A(n709), .ZN(n722) );
  NAND2_X1 U785 ( .A1(G1956), .A2(n722), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U787 ( .A1(G299), .A2(n703), .ZN(n700) );
  XOR2_X1 U788 ( .A(KEYINPUT103), .B(n700), .Z(n701) );
  NOR2_X1 U789 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U790 ( .A1(G299), .A2(n703), .ZN(n704) );
  XOR2_X1 U791 ( .A(KEYINPUT28), .B(n704), .Z(n705) );
  NOR2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U793 ( .A(n707), .B(KEYINPUT29), .ZN(n713) );
  NOR2_X1 U794 ( .A1(n709), .A2(G1961), .ZN(n708) );
  XOR2_X1 U795 ( .A(KEYINPUT98), .B(n708), .Z(n711) );
  XNOR2_X1 U796 ( .A(KEYINPUT25), .B(G2078), .ZN(n939) );
  NAND2_X1 U797 ( .A1(n709), .A2(n939), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n718) );
  NAND2_X1 U799 ( .A1(G171), .A2(n718), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n713), .A2(n712), .ZN(n734) );
  NAND2_X1 U801 ( .A1(G8), .A2(n714), .ZN(n765) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n765), .ZN(n737) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n714), .ZN(n733) );
  NOR2_X1 U804 ( .A1(n737), .A2(n733), .ZN(n715) );
  NAND2_X1 U805 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U806 ( .A(KEYINPUT30), .B(n716), .ZN(n717) );
  NOR2_X1 U807 ( .A1(G168), .A2(n717), .ZN(n720) );
  NOR2_X1 U808 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U810 ( .A(KEYINPUT31), .B(n721), .Z(n735) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n765), .ZN(n724) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n722), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U814 ( .A1(n725), .A2(G303), .ZN(n727) );
  AND2_X1 U815 ( .A1(n735), .A2(n727), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n734), .A2(n726), .ZN(n730) );
  INV_X1 U817 ( .A(n727), .ZN(n728) );
  OR2_X1 U818 ( .A1(n728), .A2(G286), .ZN(n729) );
  AND2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U821 ( .A(n732), .B(KEYINPUT32), .ZN(n741) );
  NAND2_X1 U822 ( .A1(G8), .A2(n733), .ZN(n739) );
  AND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U824 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U826 ( .A1(n741), .A2(n740), .ZN(n757) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n742) );
  NOR2_X1 U829 ( .A1(n749), .A2(n742), .ZN(n996) );
  NAND2_X1 U830 ( .A1(n757), .A2(n996), .ZN(n744) );
  NAND2_X1 U831 ( .A1(G288), .A2(G1976), .ZN(n743) );
  XNOR2_X1 U832 ( .A(n743), .B(KEYINPUT104), .ZN(n997) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n748) );
  INV_X1 U834 ( .A(KEYINPUT33), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n754) );
  NAND2_X1 U836 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U837 ( .A1(n765), .A2(n750), .ZN(n752) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n998) );
  INV_X1 U839 ( .A(n998), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n761) );
  NOR2_X1 U842 ( .A1(G2090), .A2(G303), .ZN(n755) );
  XOR2_X1 U843 ( .A(KEYINPUT105), .B(n755), .Z(n756) );
  NAND2_X1 U844 ( .A1(G8), .A2(n756), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n759), .A2(n765), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U848 ( .A(n762), .B(KEYINPUT106), .ZN(n767) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U850 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n768) );
  INV_X1 U853 ( .A(n768), .ZN(n802) );
  NOR2_X1 U854 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U855 ( .A(n771), .B(KEYINPUT92), .ZN(n814) );
  XOR2_X1 U856 ( .A(KEYINPUT96), .B(G1991), .Z(n938) );
  NAND2_X1 U857 ( .A1(G95), .A2(n883), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G131), .A2(n884), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n777) );
  NAND2_X1 U860 ( .A1(G119), .A2(n887), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G107), .A2(n888), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n866) );
  NOR2_X1 U864 ( .A1(n938), .A2(n866), .ZN(n786) );
  NAND2_X1 U865 ( .A1(G129), .A2(n887), .ZN(n779) );
  NAND2_X1 U866 ( .A1(G117), .A2(n888), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n883), .A2(G105), .ZN(n780) );
  XOR2_X1 U869 ( .A(KEYINPUT38), .B(n780), .Z(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n884), .A2(G141), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n867) );
  AND2_X1 U873 ( .A1(G1996), .A2(n867), .ZN(n785) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n961) );
  INV_X1 U875 ( .A(n961), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n814), .A2(n787), .ZN(n803) );
  NAND2_X1 U877 ( .A1(G104), .A2(n883), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G140), .A2(n884), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U880 ( .A(KEYINPUT34), .B(n790), .Z(n797) );
  NAND2_X1 U881 ( .A1(n887), .A2(G128), .ZN(n791) );
  XOR2_X1 U882 ( .A(KEYINPUT93), .B(n791), .Z(n793) );
  NAND2_X1 U883 ( .A1(n888), .A2(G116), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n795) );
  XNOR2_X1 U885 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n794) );
  XNOR2_X1 U886 ( .A(n795), .B(n794), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U888 ( .A(KEYINPUT36), .B(n798), .Z(n894) );
  XNOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  OR2_X1 U890 ( .A1(n894), .A2(n812), .ZN(n799) );
  XNOR2_X1 U891 ( .A(n799), .B(KEYINPUT95), .ZN(n972) );
  NAND2_X1 U892 ( .A1(n972), .A2(n814), .ZN(n810) );
  NAND2_X1 U893 ( .A1(n803), .A2(n810), .ZN(n800) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n989) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n817) );
  XOR2_X1 U896 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n809) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n867), .ZN(n963) );
  INV_X1 U898 ( .A(n803), .ZN(n806) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n804) );
  AND2_X1 U900 ( .A1(n938), .A2(n866), .ZN(n959) );
  NOR2_X1 U901 ( .A1(n804), .A2(n959), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n963), .A2(n807), .ZN(n808) );
  XNOR2_X1 U904 ( .A(n809), .B(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n812), .A2(n894), .ZN(n974) );
  NAND2_X1 U907 ( .A1(n813), .A2(n974), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U911 ( .A(KEYINPUT108), .B(G2454), .ZN(n827) );
  XNOR2_X1 U912 ( .A(G2430), .B(G2435), .ZN(n825) );
  XOR2_X1 U913 ( .A(G2451), .B(G2427), .Z(n820) );
  XNOR2_X1 U914 ( .A(G2438), .B(G2446), .ZN(n819) );
  XNOR2_X1 U915 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U916 ( .A(n821), .B(G2443), .Z(n823) );
  XNOR2_X1 U917 ( .A(G1341), .B(G1348), .ZN(n822) );
  XNOR2_X1 U918 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n828), .A2(G14), .ZN(n903) );
  XNOR2_X1 U922 ( .A(KEYINPUT109), .B(n903), .ZN(G401) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n829), .ZN(G217) );
  INV_X1 U924 ( .A(n829), .ZN(G223) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U926 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G188) );
  XOR2_X1 U929 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U934 ( .A(n835), .B(KEYINPUT111), .Z(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U936 ( .A(KEYINPUT112), .B(n836), .ZN(G319) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n838) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2072), .Z(n840) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2090), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U943 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1966), .B(G1981), .Z(n846) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1986), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U949 ( .A(G1976), .B(G1971), .Z(n848) );
  XNOR2_X1 U950 ( .A(G1961), .B(G1956), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U952 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U953 ( .A(KEYINPUT113), .B(G2474), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n854) );
  XOR2_X1 U955 ( .A(G1991), .B(KEYINPUT41), .Z(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G124), .A2(n887), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G100), .A2(n883), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n856), .B(KEYINPUT114), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G112), .A2(n888), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G136), .A2(n884), .ZN(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U965 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n864) );
  XNOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U969 ( .A(n865), .B(G162), .Z(n869) );
  XOR2_X1 U970 ( .A(n867), .B(n866), .Z(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n960), .B(n870), .ZN(n872) );
  XNOR2_X1 U973 ( .A(G164), .B(G160), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n882) );
  NAND2_X1 U975 ( .A1(G130), .A2(n887), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G118), .A2(n888), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n883), .A2(G106), .ZN(n875) );
  XOR2_X1 U979 ( .A(KEYINPUT115), .B(n875), .Z(n877) );
  NAND2_X1 U980 ( .A1(n884), .A2(G142), .ZN(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n878), .Z(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(n882), .B(n881), .Z(n896) );
  NAND2_X1 U985 ( .A1(G103), .A2(n883), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G139), .A2(n884), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G127), .A2(n887), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G115), .A2(n888), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n976) );
  XOR2_X1 U993 ( .A(n894), .B(n976), .Z(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U996 ( .A(n992), .B(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(G301), .B(n1005), .Z(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U999 ( .A(G286), .B(n901), .Z(n902) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n902), .ZN(G397) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n903), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1009 ( .A(G1961), .B(G5), .Z(n924) );
  XOR2_X1 U1010 ( .A(G1956), .B(G20), .Z(n911) );
  XNOR2_X1 U1011 ( .A(G1981), .B(KEYINPUT123), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(n909), .B(G6), .ZN(n910) );
  NAND2_X1 U1013 ( .A1(n911), .A2(n910), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(G19), .B(G1341), .ZN(n912) );
  NOR2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1016 ( .A(KEYINPUT124), .B(n914), .Z(n918) );
  XNOR2_X1 U1017 ( .A(KEYINPUT59), .B(G4), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(n915), .B(KEYINPUT125), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(G1348), .B(n916), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1021 ( .A(KEYINPUT60), .B(n919), .Z(n921) );
  XNOR2_X1 U1022 ( .A(G1966), .B(G21), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(KEYINPUT126), .B(n922), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(G1971), .B(G22), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(G23), .B(G1976), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n928) );
  XOR2_X1 U1029 ( .A(G1986), .B(G24), .Z(n927) );
  NAND2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(KEYINPUT58), .B(n929), .ZN(n930) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1033 ( .A(KEYINPUT61), .B(n932), .Z(n933) );
  NOR2_X1 U1034 ( .A1(G16), .A2(n933), .ZN(n957) );
  XNOR2_X1 U1035 ( .A(G2090), .B(G35), .ZN(n948) );
  XNOR2_X1 U1036 ( .A(G2067), .B(G26), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(G2072), .B(G33), .ZN(n934) );
  NOR2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1039 ( .A1(G28), .A2(n936), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(G32), .B(n937), .ZN(n943) );
  XOR2_X1 U1041 ( .A(n938), .B(G25), .Z(n941) );
  XOR2_X1 U1042 ( .A(n939), .B(G27), .Z(n940) );
  NOR2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(KEYINPUT53), .B(n946), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1048 ( .A(G2084), .B(G34), .Z(n949) );
  XNOR2_X1 U1049 ( .A(KEYINPUT54), .B(n949), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1051 ( .A(KEYINPUT55), .B(n952), .Z(n954) );
  INV_X1 U1052 ( .A(G29), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n955), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n987) );
  XOR2_X1 U1056 ( .A(G160), .B(G2084), .Z(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n970) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n968) );
  XOR2_X1 U1059 ( .A(G2090), .B(G162), .Z(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1061 ( .A(KEYINPUT51), .B(n964), .Z(n966) );
  XNOR2_X1 U1062 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(n966), .B(n965), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(KEYINPUT120), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n981) );
  XOR2_X1 U1069 ( .A(G2072), .B(n976), .Z(n978) );
  XOR2_X1 U1070 ( .A(G164), .B(G2078), .Z(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT50), .B(n979), .Z(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(KEYINPUT52), .B(n982), .ZN(n984) );
  INV_X1 U1075 ( .A(KEYINPUT55), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n985), .A2(G29), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n1014) );
  XNOR2_X1 U1079 ( .A(G1956), .B(G299), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(G1971), .A2(G303), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G1341), .B(n992), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT122), .B(n993), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1004) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G168), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(KEYINPUT57), .B(n1000), .Z(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1010) );
  XOR2_X1 U1092 ( .A(n1005), .B(G1348), .Z(n1007) );
  XNOR2_X1 U1093 ( .A(G301), .B(G1961), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(n1008), .B(KEYINPUT121), .ZN(n1009) );
  NOR2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(KEYINPUT56), .B(G16), .Z(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(n1015), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1101 ( .A(G150), .ZN(G311) );
endmodule

