//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT70), .B1(new_n195), .B2(G116), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT70), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n193), .A3(G119), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n194), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT2), .B(G113), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n199), .B(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT68), .A3(G134), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n203), .B2(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n205), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT71), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .A4(G128), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n226), .A2(KEYINPUT69), .A3(new_n222), .A4(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n220), .B2(G146), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n218), .A2(KEYINPUT65), .A3(G143), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n219), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n220), .A2(G146), .ZN(new_n233));
  OAI21_X1  g047(.A(G128), .B1(new_n233), .B2(new_n222), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n209), .A2(KEYINPUT71), .A3(new_n214), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n217), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n217), .A2(new_n236), .A3(KEYINPUT72), .A4(new_n237), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n211), .A2(new_n212), .A3(new_n205), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n211), .A2(new_n212), .A3(new_n244), .A4(new_n205), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(G131), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n214), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n226), .A2(KEYINPUT0), .A3(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n229), .A2(new_n220), .A3(G146), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n233), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT0), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n257), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n251), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n213), .B1(new_n242), .B2(KEYINPUT66), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT67), .A3(new_n245), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n250), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n240), .A2(new_n241), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT30), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n236), .A2(new_n214), .A3(new_n209), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n201), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n240), .A2(new_n201), .A3(new_n241), .A4(new_n266), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n192), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT29), .ZN(new_n276));
  INV_X1    g090(.A(new_n201), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n266), .A2(new_n238), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n266), .A2(new_n238), .A3(KEYINPUT74), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT28), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(new_n270), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n277), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n273), .B2(new_n285), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n275), .B(new_n276), .C1(new_n287), .C2(new_n192), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n267), .A2(new_n277), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n283), .B1(new_n289), .B2(new_n273), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(new_n282), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n192), .A2(new_n276), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G472), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n273), .A2(new_n191), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT73), .B1(new_n272), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n273), .A2(new_n191), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n300));
  INV_X1    g114(.A(new_n271), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(new_n267), .B2(KEYINPUT30), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n299), .B(new_n300), .C1(new_n302), .C2(new_n201), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(KEYINPUT31), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n299), .B(new_n305), .C1(new_n302), .C2(new_n201), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n192), .B1(new_n282), .B2(new_n286), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n296), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n310), .ZN(new_n312));
  AOI211_X1 g126(.A(KEYINPUT32), .B(new_n312), .C1(new_n304), .C2(new_n308), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n295), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G237), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G214), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n220), .A2(KEYINPUT89), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT89), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G143), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT18), .A2(G131), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n220), .A2(KEYINPUT89), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(G214), .A3(new_n187), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(KEYINPUT78), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(G125), .A3(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(G146), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n327), .A2(G140), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n218), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n325), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT91), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT90), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n319), .A2(G143), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n340), .A2(new_n323), .B1(new_n187), .B2(G214), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n317), .A2(new_n320), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT89), .B(G143), .ZN(new_n344));
  INV_X1    g158(.A(G214), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n345), .A2(G237), .A3(G953), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n324), .B(KEYINPUT90), .C1(new_n344), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n322), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n338), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI211_X1 g164(.A(KEYINPUT91), .B(new_n322), .C1(new_n343), .C2(new_n347), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n337), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G113), .B(G122), .ZN(new_n353));
  INV_X1    g167(.A(G104), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n332), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G146), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n218), .B1(new_n356), .B2(new_n358), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n324), .B1(new_n344), .B2(new_n346), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT17), .A3(G131), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT92), .B1(new_n363), .B2(G131), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(G131), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n321), .A2(new_n367), .A3(new_n213), .A4(new_n324), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n362), .B(new_n364), .C1(new_n369), .C2(KEYINPUT17), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n352), .A2(new_n355), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n359), .A2(G146), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT93), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n328), .A2(KEYINPUT19), .A3(new_n330), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT19), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n332), .A2(new_n333), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n372), .B(new_n373), .C1(G146), .C2(new_n377), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n374), .A2(new_n218), .A3(new_n376), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT93), .B1(new_n379), .B2(new_n361), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n369), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n352), .A2(KEYINPUT94), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n355), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT94), .B1(new_n352), .B2(new_n381), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n371), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(G475), .A2(G902), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n387), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT94), .ZN(new_n392));
  INV_X1    g206(.A(new_n347), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT90), .B1(new_n321), .B2(new_n324), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n349), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT91), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n348), .A2(new_n338), .A3(new_n349), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n336), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n378), .A2(new_n369), .A3(new_n380), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n392), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n383), .A3(new_n382), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n391), .B1(new_n401), .B2(new_n371), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT20), .ZN(new_n403));
  INV_X1    g217(.A(G902), .ZN(new_n404));
  INV_X1    g218(.A(new_n371), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n355), .B1(new_n352), .B2(new_n370), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G475), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n390), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G952), .ZN(new_n410));
  AOI211_X1 g224(.A(G953), .B(new_n410), .C1(G234), .C2(G237), .ZN(new_n411));
  INV_X1    g225(.A(G234), .ZN(new_n412));
  OAI211_X1 g226(.A(G902), .B(G953), .C1(new_n412), .C2(new_n315), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT99), .Z(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G478), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT15), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n220), .A2(G128), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n260), .A2(G143), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n420), .A3(new_n203), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT13), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n260), .B2(G143), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n220), .A2(KEYINPUT13), .A3(G128), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT96), .A4(new_n420), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT96), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n426), .A2(new_n220), .A3(KEYINPUT13), .A4(G128), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(G134), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT95), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n193), .B2(G122), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT95), .A3(G116), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G107), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n193), .A2(G122), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n421), .B(new_n428), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n430), .A2(new_n432), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT14), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n193), .A3(G122), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G107), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n419), .A2(new_n420), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G134), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n421), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT9), .B(G234), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(G217), .A3(new_n316), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n438), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT97), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT97), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n438), .A2(new_n449), .A3(new_n456), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n438), .A2(new_n449), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n452), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n460), .A2(KEYINPUT98), .A3(new_n404), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT98), .B1(new_n460), .B2(new_n404), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n418), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n418), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n460), .A2(new_n404), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n464), .B1(new_n465), .B2(KEYINPUT98), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n409), .A2(new_n416), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n314), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G221), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n451), .B2(new_n404), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n265), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n248), .B1(new_n264), .B2(new_n245), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n473), .A2(KEYINPUT82), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT3), .B1(new_n354), .B2(G107), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n434), .A3(G104), .ZN(new_n478));
  INV_X1    g292(.A(G101), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n354), .A2(G107), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n476), .A2(new_n478), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n354), .A2(G107), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n434), .A2(G104), .ZN(new_n483));
  OAI21_X1  g297(.A(G101), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n228), .A2(new_n235), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT83), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n225), .A2(new_n227), .B1(new_n232), .B2(new_n234), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT83), .A3(new_n485), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n219), .A2(new_n221), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n234), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n228), .B2(KEYINPUT81), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT81), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n225), .A2(new_n227), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n485), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n475), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT12), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n500), .B(new_n475), .C1(new_n491), .C2(new_n497), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n481), .A2(new_n484), .A3(KEYINPUT10), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n228), .B2(new_n235), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G101), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(KEYINPUT4), .A3(new_n481), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n507), .A3(G101), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n503), .B1(new_n510), .B2(new_n263), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n473), .A2(new_n474), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n511), .B(new_n513), .C1(KEYINPUT10), .C2(new_n497), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n499), .A2(new_n501), .A3(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G110), .B(G140), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n316), .A2(G227), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n228), .A2(KEYINPUT81), .ZN(new_n520));
  INV_X1    g334(.A(new_n493), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n496), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n485), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT10), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g338(.A1(new_n509), .A2(new_n262), .B1(new_n489), .B2(new_n502), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n518), .B1(new_n526), .B2(new_n513), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n512), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n519), .A2(new_n529), .A3(G469), .ZN(new_n530));
  INV_X1    g344(.A(G469), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n404), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n514), .A2(new_n528), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n518), .ZN(new_n536));
  INV_X1    g350(.A(new_n518), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n499), .A2(new_n501), .A3(new_n514), .A4(new_n537), .ZN(new_n538));
  AOI211_X1 g352(.A(G469), .B(G902), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n472), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT25), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n372), .A2(new_n334), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT79), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT23), .B1(new_n260), .B2(G119), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n544), .A2(KEYINPUT77), .B1(G119), .B2(new_n260), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n195), .A2(G128), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT77), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT23), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT76), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT23), .A2(G119), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(G128), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n260), .A2(KEYINPUT76), .A3(KEYINPUT23), .A4(G119), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n545), .A2(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G110), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n543), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n544), .A2(KEYINPUT77), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n260), .A2(G119), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n548), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n552), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n543), .A3(new_n554), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n546), .A2(new_n557), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT24), .B(G110), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n542), .B1(new_n555), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  OAI221_X1 g380(.A(new_n566), .B1(new_n553), .B2(new_n554), .C1(new_n360), .C2(new_n361), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT22), .B(G137), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n470), .A2(new_n412), .A3(G953), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n565), .B2(new_n567), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n541), .B1(new_n575), .B2(new_n404), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n565), .A2(new_n567), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n570), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n541), .A3(new_n404), .A4(new_n572), .ZN(new_n579));
  OAI21_X1  g393(.A(G217), .B1(new_n412), .B2(G902), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT75), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n575), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(G902), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI22_X1  g400(.A1(new_n576), .A2(new_n583), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT80), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI221_X1 g403(.A(KEYINPUT80), .B1(new_n584), .B2(new_n586), .C1(new_n576), .C2(new_n583), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G210), .B1(G237), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G122), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n199), .A2(KEYINPUT5), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n195), .A2(G116), .ZN(new_n599));
  OAI21_X1  g413(.A(G113), .B1(new_n599), .B2(KEYINPUT5), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT2), .B(G113), .Z(new_n603));
  NAND2_X1  g417(.A1(new_n199), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n523), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n600), .B1(new_n199), .B2(KEYINPUT5), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n196), .A2(new_n198), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n603), .A2(new_n607), .A3(new_n599), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n485), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n597), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT87), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n262), .A2(G125), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n228), .A2(new_n327), .A3(new_n235), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT7), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT85), .B(G224), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(G953), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n614), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n615), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT88), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n605), .B(new_n594), .C1(new_n509), .C2(new_n201), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n612), .A2(new_n613), .A3(KEYINPUT88), .A4(new_n619), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n618), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n404), .B1(new_n611), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n605), .B1(new_n509), .B2(new_n201), .ZN(new_n627));
  INV_X1    g441(.A(new_n594), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(KEYINPUT6), .A3(new_n623), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n617), .B(KEYINPUT84), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n614), .B(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT6), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n627), .A2(new_n633), .A3(new_n628), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n630), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n593), .B1(new_n626), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n625), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT87), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n610), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n630), .A2(new_n632), .A3(new_n634), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n404), .A3(new_n592), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(G214), .B1(G237), .B2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n540), .A2(new_n591), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n469), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G101), .ZN(G3));
  OR2_X1    g462(.A1(new_n465), .A2(G478), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n458), .B2(new_n452), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n460), .A2(new_n650), .B1(new_n454), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(G478), .A3(new_n404), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n409), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  INV_X1    g470(.A(G472), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n309), .B2(new_n404), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n312), .B1(new_n304), .B2(new_n308), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n416), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n643), .A2(new_n661), .A3(new_n644), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n540), .A2(new_n591), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n656), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  INV_X1    g480(.A(new_n409), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n467), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n663), .A2(new_n660), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NOR2_X1   g486(.A1(new_n570), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n577), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n585), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n576), .B2(new_n583), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n540), .A2(new_n645), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n660), .A2(new_n678), .A3(new_n468), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT37), .B(G110), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT101), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n679), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n411), .B1(new_n414), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n668), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n314), .A2(new_n678), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  NAND2_X1  g501(.A1(new_n298), .A2(new_n303), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n191), .B1(new_n289), .B2(new_n273), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n404), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G472), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n311), .B2(new_n313), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT102), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n539), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n515), .A2(new_n518), .B1(new_n527), .B2(new_n528), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n532), .B1(new_n696), .B2(G469), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n471), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n684), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n643), .B(KEYINPUT38), .Z(new_n703));
  INV_X1    g517(.A(new_n644), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n463), .B2(new_n466), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n409), .A2(new_n677), .A3(new_n705), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n701), .A2(new_n702), .A3(new_n703), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n694), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  INV_X1    g523(.A(new_n684), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n408), .B1(new_n402), .B2(KEYINPUT20), .ZN(new_n711));
  AOI211_X1 g525(.A(new_n389), .B(new_n391), .C1(new_n401), .C2(new_n371), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n654), .B(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n314), .A2(new_n678), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  XNOR2_X1  g530(.A(new_n659), .B(new_n296), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n591), .B1(new_n717), .B2(new_n295), .ZN(new_n718));
  AOI21_X1  g532(.A(G902), .B1(new_n536), .B2(new_n538), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT103), .B1(new_n719), .B2(new_n531), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n537), .B1(new_n514), .B2(new_n528), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n499), .A2(new_n501), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(new_n527), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n723), .B2(G902), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g539(.A(KEYINPUT103), .B(G469), .C1(new_n723), .C2(G902), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n472), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n662), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n718), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n656), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT41), .B(G113), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT104), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n731), .B(new_n733), .ZN(G15));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n669), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT105), .B(G116), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G18));
  NOR3_X1   g551(.A1(new_n728), .A2(new_n645), .A3(new_n677), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n469), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  AOI211_X1 g554(.A(new_n416), .B(new_n471), .C1(new_n725), .C2(new_n726), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n290), .A2(new_n282), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n272), .A2(new_n297), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n742), .A2(new_n192), .B1(new_n743), .B2(new_n305), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n312), .B1(new_n744), .B2(new_n304), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n658), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n643), .B(new_n705), .C1(new_n711), .C2(new_n712), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n409), .A2(KEYINPUT106), .A3(new_n643), .A4(new_n705), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n587), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n741), .A2(new_n746), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  NOR3_X1   g568(.A1(new_n658), .A2(new_n745), .A3(new_n677), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n471), .B(new_n645), .C1(new_n725), .C2(new_n726), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n714), .ZN(new_n758));
  INV_X1    g572(.A(new_n645), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n727), .A2(new_n714), .A3(new_n759), .A4(new_n472), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n298), .A2(KEYINPUT31), .A3(new_n303), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n306), .B1(new_n291), .B2(new_n191), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n310), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(G902), .B1(new_n304), .B2(new_n308), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n763), .B(new_n676), .C1(new_n657), .C2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT107), .B1(new_n760), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT108), .B(G125), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G27));
  NOR2_X1   g583(.A1(new_n643), .A2(new_n704), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n771), .A2(new_n540), .A3(new_n713), .ZN(new_n772));
  INV_X1    g586(.A(new_n591), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n314), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT42), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n314), .A2(new_n772), .A3(KEYINPUT42), .A4(new_n752), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  NOR2_X1   g593(.A1(new_n771), .A2(new_n540), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n314), .A2(new_n685), .A3(new_n773), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  AOI21_X1  g596(.A(KEYINPUT43), .B1(new_n667), .B2(new_n654), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n667), .A2(KEYINPUT43), .A3(new_n654), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n660), .A2(new_n677), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(KEYINPUT110), .A3(new_n785), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n696), .A2(KEYINPUT45), .ZN(new_n794));
  OAI21_X1  g608(.A(G469), .B1(new_n696), .B2(KEYINPUT45), .ZN(new_n795));
  OAI211_X1 g609(.A(KEYINPUT46), .B(new_n533), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT109), .A3(new_n695), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n794), .A2(new_n795), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n532), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(KEYINPUT46), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT109), .B1(new_n796), .B2(new_n695), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n472), .B(new_n699), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n788), .A2(KEYINPUT44), .A3(new_n789), .A4(new_n790), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n793), .A2(new_n770), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  OAI21_X1  g620(.A(new_n472), .B1(new_n800), .B2(new_n801), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n314), .A2(new_n773), .A3(new_n713), .A4(new_n771), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  XNOR2_X1  g626(.A(new_n727), .B(KEYINPUT49), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n704), .B(new_n471), .C1(new_n649), .C2(new_n653), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n667), .A2(new_n703), .A3(new_n752), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n693), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n767), .A2(new_n686), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n675), .B(new_n710), .C1(new_n576), .C2(new_n583), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n472), .C1(new_n534), .C2(new_n539), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n749), .B2(new_n750), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n692), .A2(new_n822), .A3(KEYINPUT113), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT113), .B1(new_n692), .B2(new_n822), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n715), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n817), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n698), .A2(new_n759), .A3(new_n676), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n717), .B2(new_n295), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n758), .A2(new_n766), .B1(new_n828), .B2(new_n685), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n692), .A2(new_n822), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n692), .A2(new_n822), .A3(KEYINPUT113), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n829), .A2(KEYINPUT52), .A3(new_n715), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n826), .A2(new_n835), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n409), .A2(new_n677), .A3(new_n467), .A4(new_n684), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n314), .A2(new_n780), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT111), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n314), .A2(new_n840), .A3(new_n780), .A4(new_n837), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n755), .A2(new_n772), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n781), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n778), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n718), .B(new_n729), .C1(new_n656), .C2(new_n669), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n668), .A2(new_n655), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n663), .A2(new_n660), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n753), .A2(new_n679), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n469), .B1(new_n646), .B2(new_n738), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n836), .A2(new_n852), .A3(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n818), .A2(KEYINPUT112), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n767), .A2(new_n855), .A3(new_n686), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n817), .B1(new_n832), .B2(new_n833), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n854), .A2(new_n715), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n818), .B2(new_n825), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(new_n852), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n853), .B1(new_n862), .B2(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n852), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n836), .A2(new_n852), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n472), .B1(new_n725), .B2(new_n726), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n809), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n786), .A2(new_n411), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n746), .A2(new_n752), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n876), .A3(new_n771), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n875), .A2(new_n876), .ZN(new_n879));
  INV_X1    g693(.A(new_n728), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n704), .A3(new_n703), .A4(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT50), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n880), .A2(new_n411), .A3(new_n773), .A4(new_n770), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n694), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n667), .A3(new_n649), .A4(new_n653), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n875), .A2(new_n728), .A3(new_n771), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n755), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT51), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n314), .A3(new_n752), .ZN(new_n892));
  NAND2_X1  g706(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n893));
  OR2_X1    g707(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n410), .B(G953), .C1(new_n879), .C2(new_n757), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n895), .B(new_n896), .C1(new_n892), .C2(new_n893), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n656), .B2(new_n885), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n878), .A2(new_n882), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n889), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n886), .A2(KEYINPUT115), .A3(new_n888), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(KEYINPUT51), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n898), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n872), .A2(new_n891), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n816), .B1(new_n905), .B2(new_n906), .ZN(G75));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n316), .A2(G952), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n404), .B1(new_n865), .B2(new_n868), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT56), .B1(new_n911), .B2(G210), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n630), .A2(new_n634), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(new_n632), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n910), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(G210), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n918), .B(new_n404), .C1(new_n865), .C2(new_n868), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n919), .A2(KEYINPUT56), .A3(new_n915), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n908), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n912), .A2(new_n916), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n915), .B1(new_n919), .B2(KEYINPUT56), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT117), .A4(new_n910), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n924), .ZN(G51));
  INV_X1    g739(.A(new_n723), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n865), .A2(new_n868), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n870), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n532), .B(KEYINPUT57), .Z(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n911), .A2(new_n798), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n909), .B1(new_n930), .B2(new_n931), .ZN(G54));
  NAND2_X1  g746(.A1(new_n927), .A2(G902), .ZN(new_n933));
  NAND2_X1  g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n371), .B(new_n401), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .A4(new_n386), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n910), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT118), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT118), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n935), .A2(new_n939), .A3(new_n910), .A4(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(G60));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT59), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n652), .B1(new_n872), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n652), .A2(new_n943), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n910), .B1(new_n928), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n946), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n584), .B1(new_n869), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n949), .B1(new_n865), .B2(new_n868), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n909), .B1(new_n951), .B2(new_n674), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n674), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(KEYINPUT119), .A3(new_n910), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n950), .B(new_n952), .C1(KEYINPUT119), .C2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(G66));
  OAI21_X1  g773(.A(G953), .B1(new_n415), .B2(new_n616), .ZN(new_n960));
  INV_X1    g774(.A(new_n851), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n913), .B1(G898), .B2(new_n316), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT120), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  AOI21_X1  g779(.A(new_n316), .B1(G227), .B2(G900), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT123), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT124), .Z(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n302), .B(new_n377), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n316), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n854), .A2(new_n708), .A3(new_n715), .A4(new_n856), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n811), .A2(new_n805), .ZN(new_n976));
  AOI211_X1 g790(.A(new_n771), .B(new_n700), .C1(new_n655), .C2(new_n668), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(new_n718), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n972), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n975), .A2(new_n978), .A3(new_n972), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n971), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n966), .A2(KEYINPUT123), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n854), .A2(new_n715), .A3(new_n856), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n314), .A2(new_n752), .A3(new_n751), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n778), .B(new_n781), .C1(new_n802), .C2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n805), .A3(new_n811), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n316), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n683), .A2(G953), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT122), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n970), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n983), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n969), .B1(new_n982), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n981), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(new_n979), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n993), .B(new_n968), .C1(new_n997), .C2(new_n971), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(G72));
  XOR2_X1   g813(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1000));
  NOR2_X1   g814(.A1(new_n657), .A2(new_n404), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n275), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n863), .B(new_n1002), .C1(new_n688), .C2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n272), .A2(new_n274), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT126), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(new_n191), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n987), .A2(new_n805), .A3(new_n811), .A4(new_n961), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(new_n1002), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1010), .A2(new_n909), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1011), .A2(KEYINPUT127), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1010), .A2(new_n1013), .A3(new_n909), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1004), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1006), .A2(new_n191), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n980), .A2(new_n961), .A3(new_n981), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(new_n1002), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1015), .A2(new_n1018), .ZN(G57));
endmodule


