//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202));
  INV_X1    g001(.A(G64gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G57gat), .ZN(new_n204));
  OR2_X1    g003(.A1(KEYINPUT91), .A2(G57gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT91), .A2(G57gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(G64gat), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n202), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT92), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n204), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n203), .A2(G57gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT9), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n208), .A2(new_n211), .B1(new_n202), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT94), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n207), .A2(new_n204), .ZN(new_n218));
  INV_X1    g017(.A(new_n202), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n211), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n202), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT94), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n217), .A2(new_n223), .A3(KEYINPUT21), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G1gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G1gat), .B2(new_n225), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G8gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT95), .ZN(new_n232));
  NAND2_X1  g031(.A1(G231gat), .A2(G233gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT93), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n232), .B(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n215), .A2(KEYINPUT21), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G155gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g039(.A(G183gat), .B(G211gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n237), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT10), .ZN(new_n245));
  NAND2_X1  g044(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(G85gat), .A3(G92gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(G85gat), .A2(G92gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT96), .A3(KEYINPUT7), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT97), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(KEYINPUT97), .A2(G99gat), .A3(G106gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(KEYINPUT8), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G85gat), .ZN(new_n256));
  INV_X1    g055(.A(G92gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(G99gat), .B(G106gat), .Z(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT98), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n247), .A2(new_n249), .B1(new_n256), .B2(new_n257), .ZN(new_n263));
  INV_X1    g062(.A(new_n260), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n255), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n263), .B2(new_n255), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT98), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n215), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n222), .B1(new_n261), .B2(new_n265), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n245), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n268), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n272), .A2(KEYINPUT10), .A3(new_n223), .A4(new_n217), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G230gat), .A2(G233gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n269), .A2(new_n270), .A3(new_n275), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G176gat), .B(G204gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  NAND3_X1  g080(.A1(new_n276), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  INV_X1    g082(.A(new_n275), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n284), .B1(new_n271), .B2(new_n273), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n285), .B2(new_n277), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT101), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n282), .A2(KEYINPUT101), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT15), .ZN(new_n292));
  INV_X1    g091(.A(G29gat), .ZN(new_n293));
  OR2_X1    g092(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G36gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n297), .A3(KEYINPUT14), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT14), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(G29gat), .B2(G36gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n292), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(KEYINPUT87), .A2(G36gat), .ZN(new_n304));
  OAI21_X1  g103(.A(G29gat), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n305), .A2(KEYINPUT15), .A3(new_n300), .A4(new_n298), .ZN(new_n306));
  XNOR2_X1  g105(.A(G43gat), .B(G50gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n296), .A2(new_n301), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(KEYINPUT15), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT88), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(KEYINPUT88), .A3(new_n311), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT17), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(KEYINPUT17), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n268), .B(new_n266), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n308), .A2(KEYINPUT88), .A3(new_n311), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT88), .B1(new_n308), .B2(new_n311), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n272), .ZN(new_n323));
  NAND3_X1  g122(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n323), .A2(KEYINPUT99), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT99), .B1(new_n323), .B2(new_n324), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n319), .B(new_n330), .C1(new_n325), .C2(new_n326), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G190gat), .B(G218gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT100), .ZN(new_n334));
  XOR2_X1   g133(.A(G134gat), .B(G162gat), .Z(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  XNOR2_X1  g135(.A(new_n332), .B(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n244), .A2(new_n291), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT89), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT17), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n320), .B2(new_n321), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n229), .B1(new_n342), .B2(new_n317), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n314), .A2(new_n229), .A3(new_n315), .ZN(new_n344));
  NAND2_X1  g143(.A1(G229gat), .A2(G233gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n340), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n230), .B1(new_n316), .B2(new_n318), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n322), .A2(new_n229), .B1(G229gat), .B2(G233gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT89), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n345), .B(KEYINPUT13), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n230), .B1(new_n320), .B2(new_n321), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(new_n344), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n343), .A2(new_n346), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n357), .B2(KEYINPUT18), .ZN(new_n358));
  XNOR2_X1  g157(.A(G113gat), .B(G141gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G197gat), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT11), .B(G169gat), .Z(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n352), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n352), .B2(new_n358), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n371));
  AND2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G141gat), .B(G148gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(G155gat), .B2(G162gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n374), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G141gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G148gat), .ZN(new_n380));
  INV_X1    g179(.A(G148gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G141gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G155gat), .B(G162gat), .ZN(new_n384));
  INV_X1    g183(.A(G155gat), .ZN(new_n385));
  INV_X1    g184(.A(G162gat), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT2), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G134gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G127gat), .ZN(new_n391));
  INV_X1    g190(.A(G127gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G134gat), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G113gat), .B(G120gat), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT1), .B1(new_n395), .B2(KEYINPUT66), .ZN(new_n396));
  INV_X1    g195(.A(G120gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G113gat), .ZN(new_n398));
  INV_X1    g197(.A(G113gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G120gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT66), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n394), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT67), .B1(new_n399), .B2(G120gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT67), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(new_n397), .A3(G113gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n407), .A3(new_n400), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT1), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n408), .A2(new_n409), .A3(new_n394), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n389), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n378), .A2(new_n388), .ZN(new_n412));
  INV_X1    g211(.A(new_n394), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT66), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n409), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n395), .A2(KEYINPUT66), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n394), .A3(new_n409), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n412), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n411), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n371), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT68), .B1(new_n404), .B2(new_n410), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT68), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n417), .A2(new_n425), .A3(new_n418), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n424), .A2(new_n426), .A3(KEYINPUT4), .A4(new_n412), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n419), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n378), .A2(new_n388), .A3(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n431), .B(new_n433), .C1(new_n404), .C2(new_n410), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(new_n434), .A3(new_n421), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n423), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  AND4_X1   g235(.A1(KEYINPUT4), .A2(new_n412), .A3(new_n417), .A4(new_n418), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n424), .A2(new_n412), .A3(new_n426), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(new_n429), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n434), .A2(new_n421), .A3(new_n371), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(G1gat), .B(G29gat), .Z(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G57gat), .B(G85gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n436), .B2(new_n441), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT79), .A3(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n441), .A3(new_n451), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n451), .B1(new_n442), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n427), .A2(new_n421), .A3(new_n434), .A4(new_n430), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n460), .A2(new_n423), .B1(new_n439), .B2(new_n440), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT80), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n457), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n454), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465));
  NAND2_X1  g264(.A1(G226gat), .A2(G233gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(G169gat), .A2(G176gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT26), .ZN(new_n469));
  NAND2_X1  g268(.A1(G169gat), .A2(G176gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n467), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT27), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(KEYINPUT65), .A3(G183gat), .ZN(new_n475));
  INV_X1    g274(.A(G190gat), .ZN(new_n476));
  AND2_X1   g275(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n475), .B(new_n476), .C1(new_n474), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT28), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G183gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(KEYINPUT28), .A3(new_n476), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n473), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G183gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G190gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(G183gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT24), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(G169gat), .B2(G176gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT24), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(G183gat), .A3(G190gat), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n470), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(KEYINPUT23), .B2(new_n467), .ZN(new_n495));
  NOR2_X1   g294(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n488), .A2(new_n493), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n496), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n467), .A2(KEYINPUT23), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n499), .A2(new_n490), .A3(new_n492), .A4(new_n470), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n491), .B1(new_n485), .B2(new_n486), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n483), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n466), .B1(new_n505), .B2(KEYINPUT29), .ZN(new_n506));
  XNOR2_X1  g305(.A(G197gat), .B(G204gat), .ZN(new_n507));
  INV_X1    g306(.A(G211gat), .ZN(new_n508));
  INV_X1    g307(.A(G218gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n507), .B1(KEYINPUT22), .B2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(G211gat), .B(G218gat), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n497), .A2(new_n502), .B1(KEYINPUT64), .B2(KEYINPUT25), .ZN(new_n514));
  OAI211_X1 g313(.A(G226gat), .B(G233gat), .C1(new_n514), .C2(new_n483), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n506), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n466), .B1(new_n505), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n515), .ZN(new_n521));
  INV_X1    g320(.A(new_n512), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n511), .B(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n516), .A2(new_n517), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n506), .A2(KEYINPUT72), .A3(new_n513), .A4(new_n515), .ZN(new_n525));
  XOR2_X1   g324(.A(G8gat), .B(G36gat), .Z(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT73), .ZN(new_n527));
  XNOR2_X1  g326(.A(G64gat), .B(G92gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n521), .A2(new_n513), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n523), .A3(new_n515), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n531), .A2(KEYINPUT81), .A3(new_n532), .A4(KEYINPUT37), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT38), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n529), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n524), .A2(new_n537), .A3(new_n525), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(KEYINPUT37), .A3(new_n532), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT81), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n535), .A2(new_n536), .A3(new_n538), .A4(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n464), .A2(new_n465), .A3(new_n530), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT6), .B1(new_n461), .B2(new_n451), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n447), .B1(new_n461), .B2(KEYINPUT80), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n436), .A2(new_n441), .A3(KEYINPUT80), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n547), .A2(new_n453), .A3(new_n450), .A4(new_n530), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n534), .A3(new_n533), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n538), .A2(new_n536), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT82), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n516), .A2(new_n517), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n521), .A2(new_n523), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n525), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(new_n537), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT38), .B1(new_n557), .B2(new_n550), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n513), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n412), .B1(new_n561), .B2(new_n432), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n433), .A2(new_n518), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(new_n513), .ZN(new_n564));
  OAI211_X1 g363(.A(G228gat), .B(G233gat), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G228gat), .A2(G233gat), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT3), .B1(new_n513), .B2(new_n518), .ZN(new_n567));
  OAI221_X1 g366(.A(new_n566), .B1(new_n513), .B2(new_n563), .C1(new_n567), .C2(new_n412), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT31), .B(G50gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n565), .B2(new_n568), .ZN(new_n572));
  XNOR2_X1  g371(.A(G78gat), .B(G106gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G22gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OR3_X1    g374(.A1(new_n571), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n571), .B2(new_n572), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n439), .A2(new_n434), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n422), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n580), .B(KEYINPUT39), .C1(new_n422), .C2(new_n420), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n582), .A3(new_n422), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n451), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT40), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n459), .A2(new_n462), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n581), .A2(KEYINPUT40), .A3(new_n451), .A4(new_n583), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT74), .B1(new_n555), .B2(new_n536), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n524), .A2(KEYINPUT30), .A3(new_n525), .A4(new_n529), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n556), .A2(KEYINPUT74), .A3(KEYINPUT30), .A4(new_n529), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n530), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n578), .B1(new_n589), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n559), .A2(KEYINPUT83), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT83), .B1(new_n559), .B2(new_n598), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n424), .A2(new_n426), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT69), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n424), .A2(KEYINPUT69), .A3(new_n426), .ZN(new_n605));
  INV_X1    g404(.A(new_n505), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n603), .A3(new_n505), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G227gat), .ZN(new_n610));
  INV_X1    g409(.A(G233gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n601), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  AOI211_X1 g413(.A(KEYINPUT34), .B(new_n612), .C1(new_n607), .C2(new_n608), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n607), .A2(new_n612), .A3(new_n608), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT32), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G15gat), .B(G43gat), .Z(new_n621));
  XNOR2_X1  g420(.A(G71gat), .B(G99gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n618), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n617), .B(KEYINPUT32), .C1(new_n619), .C2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n616), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n616), .A2(new_n624), .A3(new_n626), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(KEYINPUT36), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT70), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n624), .A3(KEYINPUT70), .A4(new_n626), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n630), .B1(new_n634), .B2(KEYINPUT36), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT75), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n592), .A2(new_n636), .A3(new_n593), .ZN(new_n637));
  NOR4_X1   g436(.A1(new_n461), .A2(new_n449), .A3(new_n456), .A4(new_n451), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT79), .B1(new_n452), .B2(KEYINPUT6), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT78), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n452), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT78), .B1(new_n461), .B2(new_n451), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n544), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n637), .A2(new_n645), .A3(new_n596), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n636), .B1(new_n592), .B2(new_n593), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n578), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n635), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n599), .A2(new_n600), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n627), .A2(new_n578), .A3(KEYINPUT35), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n633), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n594), .B(new_n596), .C1(new_n454), .C2(new_n463), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT84), .ZN(new_n655));
  INV_X1    g454(.A(new_n578), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n628), .A2(new_n656), .A3(new_n629), .ZN(new_n657));
  OR3_X1    g456(.A1(new_n657), .A2(new_n646), .A3(new_n647), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n653), .A2(new_n655), .B1(new_n658), .B2(KEYINPUT35), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n370), .B1(new_n650), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n559), .A2(new_n598), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT83), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n559), .A2(new_n598), .A3(KEYINPUT83), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n648), .A4(new_n635), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n655), .A2(new_n653), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n658), .A2(KEYINPUT35), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n668), .A3(KEYINPUT85), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n369), .B1(new_n660), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n645), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n597), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT103), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n676), .A3(new_n597), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(G8gat), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND4_X1  g478(.A1(new_n670), .A2(KEYINPUT42), .A3(new_n597), .A4(new_n679), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n675), .A2(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n679), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n682), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n679), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n675), .B2(new_n677), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(KEYINPUT104), .A3(new_n685), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n681), .B1(new_n687), .B2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n670), .ZN(new_n692));
  OAI21_X1  g491(.A(G15gat), .B1(new_n692), .B2(new_n635), .ZN(new_n693));
  INV_X1    g492(.A(new_n634), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n692), .B2(new_n695), .ZN(G1326gat));
  NAND2_X1  g495(.A1(new_n670), .A2(new_n578), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT43), .B(G22gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  NAND2_X1  g498(.A1(new_n660), .A2(new_n669), .ZN(new_n700));
  INV_X1    g499(.A(new_n336), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n332), .B(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n291), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n244), .A2(new_n367), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n293), .A3(new_n671), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT45), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n337), .B1(new_n665), .B2(new_n668), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n337), .B1(new_n660), .B2(new_n669), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n704), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n645), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n708), .A2(new_n715), .ZN(G1328gat));
  NOR2_X1   g515(.A1(new_n303), .A2(new_n304), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n706), .A2(new_n597), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT105), .B(KEYINPUT46), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n592), .A2(new_n593), .B1(new_n595), .B2(new_n530), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n717), .B2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(new_n635), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G43gat), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n705), .A2(new_n694), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n714), .A2(new_n725), .B1(new_n726), .B2(G43gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g527(.A(new_n710), .B1(new_n700), .B2(new_n702), .ZN(new_n729));
  INV_X1    g528(.A(new_n711), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n578), .B(new_n704), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n713), .A2(new_n733), .A3(new_n578), .A4(new_n704), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(G50gat), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n656), .A2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n705), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n705), .A2(new_n738), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n731), .A2(G50gat), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n739), .B1(new_n738), .B2(new_n705), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n736), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1331gat));
  NAND4_X1  g546(.A1(new_n244), .A2(new_n367), .A3(new_n337), .A4(new_n703), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n665), .B2(new_n668), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n671), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n205), .A2(new_n206), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1332gat));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n597), .B1(new_n753), .B2(new_n203), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT108), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n203), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  XOR2_X1   g557(.A(new_n634), .B(KEYINPUT109), .Z(new_n759));
  AOI21_X1  g558(.A(G71gat), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n724), .A2(G71gat), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n760), .B1(new_n749), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n578), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT112), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT111), .B(G78gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n244), .A2(new_n368), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n713), .A2(new_n703), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n645), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n709), .A2(new_n770), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n709), .A2(KEYINPUT51), .A3(new_n770), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n291), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n256), .A3(new_n671), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(G1336gat));
  NAND2_X1  g578(.A1(new_n770), .A2(new_n703), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n700), .A2(new_n702), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT44), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n782), .B2(new_n711), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n257), .B1(new_n783), .B2(new_n597), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n721), .A2(G92gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n777), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT52), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G92gat), .B1(new_n771), .B2(new_n721), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n790), .A3(new_n786), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n791), .ZN(G1337gat));
  OAI21_X1  g591(.A(G99gat), .B1(new_n771), .B2(new_n635), .ZN(new_n793));
  INV_X1    g592(.A(G99gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n794), .A3(new_n634), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(G1338gat));
  INV_X1    g595(.A(G106gat), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n783), .B2(new_n578), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n656), .A2(G106gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n777), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT53), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G106gat), .B1(new_n771), .B2(new_n656), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(new_n800), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(G1339gat));
  NOR2_X1   g605(.A1(new_n338), .A2(new_n368), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n352), .A2(new_n358), .A3(new_n364), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n345), .B1(new_n348), .B2(new_n344), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n355), .A2(new_n344), .A3(new_n354), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n362), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n271), .A2(new_n284), .A3(new_n273), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n276), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n281), .B1(new_n285), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n816), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n282), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n702), .A2(new_n812), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n289), .A2(new_n808), .A3(new_n290), .A4(new_n811), .ZN(new_n824));
  OAI211_X1 g623(.A(KEYINPUT114), .B(new_n824), .C1(new_n367), .C2(new_n821), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n337), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n820), .A2(new_n282), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(new_n819), .C1(new_n366), .C2(new_n365), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT114), .B1(new_n828), .B2(new_n824), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n823), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n807), .B1(new_n830), .B2(new_n243), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n831), .A2(new_n645), .A3(new_n657), .A4(new_n597), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n399), .A3(new_n368), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n243), .ZN(new_n834));
  INV_X1    g633(.A(new_n807), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(KEYINPUT115), .A3(new_n656), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n831), .B2(new_n578), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n597), .A2(new_n645), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n634), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n399), .B1(new_n842), .B2(new_n368), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n833), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n832), .B2(new_n703), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n291), .A2(new_n397), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n842), .B2(new_n849), .ZN(G1341gat));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n392), .A3(new_n244), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n842), .A2(new_n244), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n392), .ZN(G1342gat));
  NAND3_X1  g652(.A1(new_n832), .A2(new_n390), .A3(new_n702), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT56), .Z(new_n855));
  AND2_X1   g654(.A1(new_n842), .A2(new_n702), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n390), .B2(new_n856), .ZN(G1343gat));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n656), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n824), .B1(new_n367), .B2(new_n821), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n337), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n823), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n243), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n862), .B1(new_n835), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n337), .A3(new_n825), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n244), .B1(new_n870), .B2(new_n823), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n578), .B1(new_n871), .B2(new_n807), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n867), .B1(new_n872), .B2(new_n860), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n635), .A2(new_n841), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n859), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n874), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n836), .B2(new_n578), .ZN(new_n877));
  OAI211_X1 g676(.A(KEYINPUT117), .B(new_n876), .C1(new_n877), .C2(new_n867), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n878), .A3(new_n368), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G141gat), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n724), .A2(new_n656), .A3(new_n597), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n671), .B(new_n881), .C1(new_n871), .C2(new_n807), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n367), .A2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n858), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n368), .B(new_n876), .C1(new_n877), .C2(new_n867), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G141gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n858), .B1(new_n882), .B2(new_n884), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n888), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT118), .B(new_n891), .C1(new_n889), .C2(G141gat), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT119), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n885), .B1(new_n879), .B2(G141gat), .ZN(new_n898));
  OAI221_X1 g697(.A(new_n897), .B1(new_n893), .B2(new_n894), .C1(new_n898), .C2(new_n858), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(G1344gat));
  AOI21_X1  g699(.A(new_n244), .B1(new_n865), .B2(KEYINPUT120), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(KEYINPUT120), .B2(new_n865), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n835), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n903), .B2(new_n578), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n831), .A2(new_n862), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(new_n703), .A3(new_n876), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT59), .B1(new_n907), .B2(new_n381), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n381), .A2(KEYINPUT59), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n875), .A2(new_n878), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n291), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n882), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n381), .A3(new_n703), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n910), .B2(new_n243), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n385), .A3(new_n244), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1346gat));
  NOR3_X1   g717(.A1(new_n910), .A2(new_n386), .A3(new_n337), .ZN(new_n919));
  AOI21_X1  g718(.A(G162gat), .B1(new_n913), .B2(new_n702), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n657), .A2(new_n721), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT121), .Z(new_n923));
  NAND3_X1  g722(.A1(new_n836), .A2(new_n645), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n368), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n671), .A2(new_n721), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n759), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT122), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n840), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n368), .A2(G169gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(G1348gat));
  OAI21_X1  g732(.A(G176gat), .B1(new_n930), .B2(new_n291), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n924), .A2(G176gat), .A3(new_n291), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  NAND3_X1  g735(.A1(new_n925), .A2(new_n481), .A3(new_n244), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n930), .A2(new_n243), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(KEYINPUT123), .ZN(new_n939));
  OAI21_X1  g738(.A(G183gat), .B1(new_n938), .B2(KEYINPUT123), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT60), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n943), .B(new_n937), .C1(new_n939), .C2(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n930), .B2(new_n337), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT61), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n476), .A3(new_n702), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1351gat));
  NAND3_X1  g748(.A1(new_n635), .A2(new_n578), .A3(new_n597), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT124), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n951), .A2(new_n671), .A3(new_n831), .ZN(new_n952));
  XNOR2_X1  g751(.A(KEYINPUT125), .B(G197gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n368), .A3(new_n953), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT126), .Z(new_n955));
  AND2_X1   g754(.A1(new_n635), .A2(new_n927), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n906), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(new_n367), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n958), .B2(new_n953), .ZN(G1352gat));
  OAI21_X1  g758(.A(G204gat), .B1(new_n957), .B2(new_n291), .ZN(new_n960));
  INV_X1    g759(.A(G204gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n952), .A2(new_n961), .A3(new_n703), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(G1353gat));
  NAND3_X1  g763(.A1(new_n952), .A2(new_n508), .A3(new_n244), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n244), .B(new_n956), .C1(new_n904), .C2(new_n905), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G211gat), .ZN(new_n967));
  NOR2_X1   g766(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n967), .A2(new_n968), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(G218gat), .B1(new_n957), .B2(new_n337), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n952), .A2(new_n509), .A3(new_n702), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1355gat));
endmodule


