

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732;

  XNOR2_X1 U372 ( .A(n496), .B(n495), .ZN(n505) );
  OR2_X1 U373 ( .A1(n493), .A2(n492), .ZN(n496) );
  NAND2_X2 U374 ( .A1(n510), .A2(n408), .ZN(n409) );
  NAND2_X1 U375 ( .A1(n710), .A2(n725), .ZN(n652) );
  XNOR2_X2 U376 ( .A(n532), .B(n531), .ZN(n710) );
  XNOR2_X2 U377 ( .A(n395), .B(KEYINPUT80), .ZN(n510) );
  NOR2_X2 U378 ( .A1(n497), .A2(n675), .ZN(n395) );
  OR2_X2 U379 ( .A1(n622), .A2(G902), .ZN(n407) );
  XNOR2_X2 U380 ( .A(n394), .B(n393), .ZN(n513) );
  OR2_X2 U381 ( .A1(n629), .A2(G902), .ZN(n394) );
  AND2_X2 U382 ( .A1(n628), .A2(n486), .ZN(n488) );
  XNOR2_X1 U383 ( .A(n652), .B(KEYINPUT2), .ZN(n355) );
  AND2_X1 U384 ( .A1(n619), .A2(n353), .ZN(n525) );
  AND2_X1 U385 ( .A1(n357), .A2(n558), .ZN(n575) );
  XNOR2_X1 U386 ( .A(n437), .B(KEYINPUT19), .ZN(n545) );
  XNOR2_X1 U387 ( .A(n463), .B(n462), .ZN(n518) );
  OR2_X1 U388 ( .A1(n540), .A2(n668), .ZN(n675) );
  XNOR2_X1 U389 ( .A(n432), .B(n431), .ZN(n559) );
  XNOR2_X1 U390 ( .A(n513), .B(KEYINPUT1), .ZN(n497) );
  XNOR2_X1 U391 ( .A(n419), .B(n382), .ZN(n459) );
  BUF_X1 U392 ( .A(n697), .Z(n350) );
  AND2_X2 U393 ( .A1(n355), .A2(n354), .ZN(n697) );
  BUF_X1 U394 ( .A(n652), .Z(n351) );
  XNOR2_X2 U395 ( .A(n459), .B(n384), .ZN(n724) );
  XNOR2_X1 U396 ( .A(n672), .B(KEYINPUT107), .ZN(n555) );
  XNOR2_X1 U397 ( .A(G146), .B(G125), .ZN(n412) );
  XNOR2_X1 U398 ( .A(n654), .B(n653), .ZN(n689) );
  NAND2_X1 U399 ( .A1(n507), .A2(n669), .ZN(n640) );
  NOR2_X1 U400 ( .A1(n549), .A2(KEYINPUT71), .ZN(n551) );
  INV_X1 U401 ( .A(KEYINPUT106), .ZN(n520) );
  NAND2_X1 U402 ( .A1(n436), .A2(n435), .ZN(n437) );
  XNOR2_X1 U403 ( .A(n356), .B(n473), .ZN(n367) );
  XNOR2_X1 U404 ( .A(n366), .B(n363), .ZN(n356) );
  XNOR2_X1 U405 ( .A(KEYINPUT77), .B(KEYINPUT23), .ZN(n363) );
  INV_X1 U406 ( .A(G134), .ZN(n382) );
  XNOR2_X1 U407 ( .A(KEYINPUT85), .B(KEYINPUT2), .ZN(n653) );
  INV_X1 U408 ( .A(n656), .ZN(n358) );
  BUF_X1 U409 ( .A(n559), .Z(n596) );
  OR2_X1 U410 ( .A1(n675), .A2(n544), .ZN(n552) );
  AND2_X1 U411 ( .A1(n505), .A2(n565), .ZN(n523) );
  INV_X2 U412 ( .A(G953), .ZN(n726) );
  INV_X1 U413 ( .A(n600), .ZN(n354) );
  AND2_X1 U414 ( .A1(n607), .A2(G953), .ZN(n709) );
  NOR2_X1 U415 ( .A1(n695), .A2(G953), .ZN(n696) );
  INV_X1 U416 ( .A(n640), .ZN(n641) );
  XNOR2_X1 U417 ( .A(n412), .B(KEYINPUT10), .ZN(n473) );
  AND2_X1 U418 ( .A1(G217), .A2(n378), .ZN(n352) );
  AND2_X1 U419 ( .A1(n640), .A2(KEYINPUT70), .ZN(n353) );
  NOR2_X2 U420 ( .A1(n599), .A2(n598), .ZN(n725) );
  AND2_X1 U421 ( .A1(n557), .A2(n358), .ZN(n357) );
  AND2_X1 U422 ( .A1(n558), .A2(n557), .ZN(n360) );
  AND2_X1 U423 ( .A1(n360), .A2(n359), .ZN(n560) );
  INV_X1 U424 ( .A(n596), .ZN(n359) );
  XNOR2_X1 U425 ( .A(KEYINPUT18), .B(KEYINPUT82), .ZN(n410) );
  INV_X1 U426 ( .A(KEYINPUT47), .ZN(n550) );
  INV_X1 U427 ( .A(KEYINPUT24), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  BUF_X1 U429 ( .A(n513), .Z(n544) );
  BUF_X1 U430 ( .A(n493), .Z(n511) );
  XOR2_X1 U431 ( .A(KEYINPUT96), .B(G140), .Z(n362) );
  XNOR2_X1 U432 ( .A(G119), .B(G110), .ZN(n361) );
  XNOR2_X1 U433 ( .A(n362), .B(n361), .ZN(n368) );
  XNOR2_X1 U434 ( .A(G137), .B(G128), .ZN(n365) );
  XOR2_X1 U435 ( .A(n368), .B(n367), .Z(n372) );
  NAND2_X1 U436 ( .A1(n726), .A2(G234), .ZN(n370) );
  XNOR2_X1 U437 ( .A(KEYINPUT73), .B(KEYINPUT8), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n452) );
  NAND2_X1 U439 ( .A1(G221), .A2(n452), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n707) );
  NOR2_X1 U441 ( .A1(n707), .A2(G902), .ZN(n377) );
  XOR2_X1 U442 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n375) );
  XNOR2_X1 U443 ( .A(KEYINPUT91), .B(KEYINPUT15), .ZN(n373) );
  INV_X1 U444 ( .A(G902), .ZN(n430) );
  XNOR2_X1 U445 ( .A(n373), .B(n430), .ZN(n600) );
  NAND2_X1 U446 ( .A1(G234), .A2(n600), .ZN(n374) );
  XNOR2_X1 U447 ( .A(KEYINPUT20), .B(n374), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n375), .B(n352), .ZN(n376) );
  XNOR2_X1 U449 ( .A(n377), .B(n376), .ZN(n540) );
  AND2_X1 U450 ( .A1(n378), .A2(G221), .ZN(n380) );
  INV_X1 U451 ( .A(KEYINPUT21), .ZN(n379) );
  XNOR2_X1 U452 ( .A(n380), .B(n379), .ZN(n668) );
  XNOR2_X2 U453 ( .A(KEYINPUT66), .B(G143), .ZN(n381) );
  XNOR2_X2 U454 ( .A(n381), .B(G128), .ZN(n419) );
  XNOR2_X1 U455 ( .A(KEYINPUT65), .B(KEYINPUT72), .ZN(n383) );
  XNOR2_X1 U456 ( .A(n383), .B(KEYINPUT4), .ZN(n420) );
  XNOR2_X1 U457 ( .A(n420), .B(G137), .ZN(n384) );
  XNOR2_X1 U458 ( .A(KEYINPUT69), .B(G101), .ZN(n415) );
  XNOR2_X1 U459 ( .A(n415), .B(G146), .ZN(n385) );
  XNOR2_X2 U460 ( .A(n724), .B(n385), .ZN(n404) );
  XNOR2_X1 U461 ( .A(G110), .B(G107), .ZN(n387) );
  INV_X1 U462 ( .A(G104), .ZN(n386) );
  XNOR2_X1 U463 ( .A(n387), .B(n386), .ZN(n425) );
  INV_X1 U464 ( .A(n425), .ZN(n391) );
  XOR2_X1 U465 ( .A(G131), .B(G140), .Z(n474) );
  XNOR2_X1 U466 ( .A(KEYINPUT81), .B(n474), .ZN(n389) );
  NAND2_X1 U467 ( .A1(n726), .A2(G227), .ZN(n388) );
  XNOR2_X1 U468 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U469 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U470 ( .A(n404), .B(n392), .ZN(n629) );
  XNOR2_X1 U471 ( .A(KEYINPUT75), .B(G469), .ZN(n393) );
  XNOR2_X1 U472 ( .A(KEYINPUT76), .B(KEYINPUT3), .ZN(n396) );
  XNOR2_X1 U473 ( .A(n396), .B(G119), .ZN(n398) );
  XOR2_X1 U474 ( .A(G113), .B(G116), .Z(n397) );
  XNOR2_X1 U475 ( .A(n398), .B(n397), .ZN(n427) );
  NOR2_X1 U476 ( .A1(G953), .A2(G237), .ZN(n470) );
  NAND2_X1 U477 ( .A1(n470), .A2(G210), .ZN(n399) );
  XNOR2_X1 U478 ( .A(n399), .B(G131), .ZN(n401) );
  XNOR2_X1 U479 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n400) );
  XNOR2_X1 U480 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U481 ( .A(n427), .B(n402), .ZN(n403) );
  XNOR2_X1 U482 ( .A(n404), .B(n403), .ZN(n622) );
  INV_X1 U483 ( .A(KEYINPUT99), .ZN(n405) );
  XNOR2_X1 U484 ( .A(n405), .B(G472), .ZN(n406) );
  XNOR2_X2 U485 ( .A(n407), .B(n406), .ZN(n672) );
  XNOR2_X1 U486 ( .A(n672), .B(KEYINPUT6), .ZN(n565) );
  INV_X1 U487 ( .A(n565), .ZN(n408) );
  XNOR2_X2 U488 ( .A(n409), .B(KEYINPUT33), .ZN(n690) );
  XNOR2_X1 U489 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n411) );
  XNOR2_X1 U490 ( .A(n411), .B(n410), .ZN(n413) );
  XNOR2_X1 U491 ( .A(n413), .B(n412), .ZN(n418) );
  NAND2_X1 U492 ( .A1(G224), .A2(n726), .ZN(n414) );
  XNOR2_X1 U493 ( .A(n414), .B(KEYINPUT89), .ZN(n416) );
  XNOR2_X1 U494 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U495 ( .A(n418), .B(n417), .ZN(n422) );
  XNOR2_X1 U496 ( .A(n419), .B(n420), .ZN(n421) );
  XNOR2_X1 U497 ( .A(n422), .B(n421), .ZN(n428) );
  XNOR2_X1 U498 ( .A(KEYINPUT78), .B(KEYINPUT16), .ZN(n423) );
  XNOR2_X1 U499 ( .A(n423), .B(G122), .ZN(n424) );
  XNOR2_X1 U500 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U501 ( .A(n427), .B(n426), .ZN(n717) );
  XNOR2_X1 U502 ( .A(n428), .B(n717), .ZN(n601) );
  NAND2_X1 U503 ( .A1(n601), .A2(n600), .ZN(n432) );
  INV_X1 U504 ( .A(G237), .ZN(n429) );
  NAND2_X1 U505 ( .A1(n430), .A2(n429), .ZN(n433) );
  NAND2_X1 U506 ( .A1(n433), .A2(G210), .ZN(n431) );
  INV_X1 U507 ( .A(n559), .ZN(n436) );
  NAND2_X1 U508 ( .A1(n433), .A2(G214), .ZN(n434) );
  XNOR2_X1 U509 ( .A(n434), .B(KEYINPUT93), .ZN(n655) );
  INV_X1 U510 ( .A(n655), .ZN(n435) );
  NAND2_X1 U511 ( .A1(G234), .A2(G237), .ZN(n439) );
  INV_X1 U512 ( .A(KEYINPUT14), .ZN(n438) );
  XNOR2_X1 U513 ( .A(n439), .B(n438), .ZN(n687) );
  INV_X1 U514 ( .A(n687), .ZN(n538) );
  NAND2_X1 U515 ( .A1(G953), .A2(G902), .ZN(n533) );
  OR2_X1 U516 ( .A1(G898), .A2(n533), .ZN(n440) );
  NAND2_X1 U517 ( .A1(G952), .A2(n726), .ZN(n534) );
  NAND2_X1 U518 ( .A1(n440), .A2(n534), .ZN(n441) );
  NAND2_X1 U519 ( .A1(n538), .A2(n441), .ZN(n442) );
  NAND2_X1 U520 ( .A1(n442), .A2(KEYINPUT94), .ZN(n447) );
  NOR2_X1 U521 ( .A1(G898), .A2(KEYINPUT94), .ZN(n444) );
  INV_X1 U522 ( .A(n533), .ZN(n443) );
  NAND2_X1 U523 ( .A1(n444), .A2(n443), .ZN(n445) );
  OR2_X1 U524 ( .A1(n687), .A2(n445), .ZN(n446) );
  AND2_X1 U525 ( .A1(n447), .A2(n446), .ZN(n448) );
  NAND2_X1 U526 ( .A1(n545), .A2(n448), .ZN(n449) );
  XNOR2_X1 U527 ( .A(n449), .B(KEYINPUT0), .ZN(n493) );
  XNOR2_X1 U528 ( .A(n511), .B(KEYINPUT95), .ZN(n514) );
  NAND2_X1 U529 ( .A1(n690), .A2(n514), .ZN(n451) );
  INV_X1 U530 ( .A(KEYINPUT34), .ZN(n450) );
  XNOR2_X1 U531 ( .A(n451), .B(n450), .ZN(n481) );
  XOR2_X1 U532 ( .A(G122), .B(KEYINPUT103), .Z(n454) );
  NAND2_X1 U533 ( .A1(G217), .A2(n452), .ZN(n453) );
  XNOR2_X1 U534 ( .A(n454), .B(n453), .ZN(n458) );
  XOR2_X1 U535 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n456) );
  XNOR2_X1 U536 ( .A(G116), .B(G107), .ZN(n455) );
  XNOR2_X1 U537 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U538 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U539 ( .A(n459), .B(n460), .ZN(n703) );
  NOR2_X1 U540 ( .A1(G902), .A2(n703), .ZN(n461) );
  XOR2_X1 U541 ( .A(n461), .B(KEYINPUT104), .Z(n463) );
  INV_X1 U542 ( .A(G478), .ZN(n462) );
  INV_X1 U543 ( .A(n518), .ZN(n480) );
  XNOR2_X1 U544 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n477) );
  XOR2_X1 U545 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n465) );
  XNOR2_X1 U546 ( .A(G143), .B(G122), .ZN(n464) );
  XNOR2_X1 U547 ( .A(n465), .B(n464), .ZN(n469) );
  XOR2_X1 U548 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n467) );
  XNOR2_X1 U549 ( .A(G113), .B(G104), .ZN(n466) );
  XNOR2_X1 U550 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U551 ( .A(n469), .B(n468), .Z(n472) );
  NAND2_X1 U552 ( .A1(G214), .A2(n470), .ZN(n471) );
  XNOR2_X1 U553 ( .A(n472), .B(n471), .ZN(n475) );
  XNOR2_X1 U554 ( .A(n474), .B(n473), .ZN(n723) );
  XNOR2_X1 U555 ( .A(n475), .B(n723), .ZN(n698) );
  NOR2_X1 U556 ( .A1(G902), .A2(n698), .ZN(n476) );
  XNOR2_X1 U557 ( .A(n477), .B(n476), .ZN(n479) );
  INV_X1 U558 ( .A(G475), .ZN(n478) );
  XNOR2_X1 U559 ( .A(n479), .B(n478), .ZN(n489) );
  INV_X1 U560 ( .A(n489), .ZN(n517) );
  AND2_X1 U561 ( .A1(n480), .A2(n517), .ZN(n561) );
  NAND2_X1 U562 ( .A1(n481), .A2(n561), .ZN(n484) );
  INV_X1 U563 ( .A(KEYINPUT86), .ZN(n482) );
  XNOR2_X1 U564 ( .A(n482), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X2 U565 ( .A(n484), .B(n483), .ZN(n628) );
  INV_X1 U566 ( .A(KEYINPUT44), .ZN(n485) );
  AND2_X1 U567 ( .A1(n485), .A2(KEYINPUT70), .ZN(n486) );
  NOR2_X1 U568 ( .A1(n628), .A2(KEYINPUT70), .ZN(n487) );
  NOR2_X1 U569 ( .A1(n488), .A2(n487), .ZN(n509) );
  NAND2_X1 U570 ( .A1(n518), .A2(n489), .ZN(n658) );
  INV_X1 U571 ( .A(n658), .ZN(n491) );
  INV_X1 U572 ( .A(n668), .ZN(n490) );
  NAND2_X1 U573 ( .A1(n491), .A2(n490), .ZN(n492) );
  INV_X1 U574 ( .A(KEYINPUT68), .ZN(n494) );
  XNOR2_X1 U575 ( .A(n494), .B(KEYINPUT22), .ZN(n495) );
  BUF_X1 U576 ( .A(n540), .Z(n669) );
  INV_X1 U577 ( .A(n669), .ZN(n501) );
  BUF_X1 U578 ( .A(n497), .Z(n498) );
  INV_X1 U579 ( .A(KEYINPUT90), .ZN(n499) );
  XNOR2_X1 U580 ( .A(n498), .B(n499), .ZN(n568) );
  INV_X1 U581 ( .A(n568), .ZN(n500) );
  NOR2_X1 U582 ( .A1(n501), .A2(n500), .ZN(n502) );
  NAND2_X1 U583 ( .A1(n523), .A2(n502), .ZN(n503) );
  XNOR2_X2 U584 ( .A(n503), .B(KEYINPUT32), .ZN(n619) );
  AND2_X1 U585 ( .A1(n498), .A2(n555), .ZN(n504) );
  NAND2_X1 U586 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U587 ( .A(n506), .B(KEYINPUT67), .ZN(n507) );
  NAND2_X1 U588 ( .A1(n619), .A2(n640), .ZN(n508) );
  NOR2_X1 U589 ( .A1(n509), .A2(n508), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n510), .A2(n672), .ZN(n667) );
  NOR2_X1 U591 ( .A1(n667), .A2(n511), .ZN(n512) );
  XNOR2_X1 U592 ( .A(n512), .B(KEYINPUT31), .ZN(n644) );
  NOR2_X1 U593 ( .A1(n552), .A2(n672), .ZN(n515) );
  NAND2_X1 U594 ( .A1(n515), .A2(n514), .ZN(n636) );
  AND2_X1 U595 ( .A1(n644), .A2(n636), .ZN(n519) );
  NOR2_X1 U596 ( .A1(n518), .A2(n517), .ZN(n516) );
  XNOR2_X1 U597 ( .A(n516), .B(KEYINPUT105), .ZN(n648) );
  NAND2_X1 U598 ( .A1(n518), .A2(n517), .ZN(n645) );
  AND2_X1 U599 ( .A1(n648), .A2(n645), .ZN(n660) );
  NOR2_X1 U600 ( .A1(n519), .A2(n660), .ZN(n521) );
  XNOR2_X1 U601 ( .A(n521), .B(n520), .ZN(n524) );
  INV_X1 U602 ( .A(n498), .ZN(n593) );
  NOR2_X1 U603 ( .A1(n669), .A2(n593), .ZN(n522) );
  NAND2_X1 U604 ( .A1(n523), .A2(n522), .ZN(n634) );
  AND2_X1 U605 ( .A1(n524), .A2(n634), .ZN(n528) );
  NAND2_X1 U606 ( .A1(n628), .A2(n525), .ZN(n526) );
  NAND2_X1 U607 ( .A1(n526), .A2(KEYINPUT44), .ZN(n527) );
  NAND2_X1 U608 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X2 U609 ( .A1(n530), .A2(n529), .ZN(n532) );
  XOR2_X1 U610 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n531) );
  NOR2_X1 U611 ( .A1(G900), .A2(n533), .ZN(n536) );
  INV_X1 U612 ( .A(n534), .ZN(n535) );
  OR2_X1 U613 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U614 ( .A1(n538), .A2(n537), .ZN(n553) );
  NOR2_X1 U615 ( .A1(n668), .A2(n553), .ZN(n539) );
  AND2_X1 U616 ( .A1(n540), .A2(n539), .ZN(n564) );
  INV_X1 U617 ( .A(n564), .ZN(n541) );
  NOR2_X1 U618 ( .A1(n541), .A2(n555), .ZN(n543) );
  XNOR2_X1 U619 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n542) );
  XNOR2_X1 U620 ( .A(n543), .B(n542), .ZN(n582) );
  XNOR2_X1 U621 ( .A(n544), .B(KEYINPUT110), .ZN(n581) );
  INV_X1 U622 ( .A(n581), .ZN(n546) );
  NAND2_X1 U623 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X2 U624 ( .A1(n582), .A2(n547), .ZN(n548) );
  NOR2_X1 U625 ( .A1(n548), .A2(n648), .ZN(n613) );
  NOR2_X1 U626 ( .A1(n548), .A2(n645), .ZN(n617) );
  NOR2_X1 U627 ( .A1(n613), .A2(n617), .ZN(n549) );
  XNOR2_X1 U628 ( .A(n551), .B(n550), .ZN(n572) );
  XNOR2_X1 U629 ( .A(n552), .B(KEYINPUT108), .ZN(n554) );
  NOR2_X1 U630 ( .A1(n554), .A2(n553), .ZN(n558) );
  NOR2_X1 U631 ( .A1(n555), .A2(n655), .ZN(n556) );
  XNOR2_X1 U632 ( .A(n556), .B(KEYINPUT30), .ZN(n557) );
  XOR2_X1 U633 ( .A(n560), .B(KEYINPUT109), .Z(n562) );
  NAND2_X1 U634 ( .A1(n562), .A2(n561), .ZN(n643) );
  NOR2_X1 U635 ( .A1(n645), .A2(n655), .ZN(n563) );
  NAND2_X1 U636 ( .A1(n564), .A2(n563), .ZN(n566) );
  OR2_X1 U637 ( .A1(n566), .A2(n565), .ZN(n594) );
  NOR2_X1 U638 ( .A1(n594), .A2(n596), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT36), .ZN(n569) );
  AND2_X1 U640 ( .A1(n569), .A2(n568), .ZN(n650) );
  INV_X1 U641 ( .A(n650), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n643), .A2(n570), .ZN(n571) );
  NOR2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U644 ( .A(n573), .B(KEYINPUT74), .ZN(n588) );
  XNOR2_X1 U645 ( .A(KEYINPUT79), .B(KEYINPUT38), .ZN(n574) );
  XNOR2_X1 U646 ( .A(n596), .B(n574), .ZN(n656) );
  XNOR2_X1 U647 ( .A(n575), .B(KEYINPUT39), .ZN(n590) );
  NOR2_X1 U648 ( .A1(n590), .A2(n645), .ZN(n577) );
  XOR2_X1 U649 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n576) );
  XNOR2_X1 U650 ( .A(n577), .B(n576), .ZN(n616) );
  NOR2_X1 U651 ( .A1(n656), .A2(n655), .ZN(n578) );
  XNOR2_X1 U652 ( .A(n578), .B(KEYINPUT113), .ZN(n659) );
  NOR2_X1 U653 ( .A1(n659), .A2(n658), .ZN(n580) );
  XOR2_X1 U654 ( .A(KEYINPUT114), .B(KEYINPUT41), .Z(n579) );
  XNOR2_X1 U655 ( .A(n580), .B(n579), .ZN(n691) );
  NOR2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n691), .A2(n583), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n584), .B(KEYINPUT42), .ZN(n614) );
  NAND2_X1 U659 ( .A1(n616), .A2(n614), .ZN(n586) );
  XNOR2_X1 U660 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n585) );
  XNOR2_X1 U661 ( .A(n586), .B(n585), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U663 ( .A(n589), .B(KEYINPUT48), .ZN(n599) );
  INV_X1 U664 ( .A(n590), .ZN(n592) );
  INV_X1 U665 ( .A(n648), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n615) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U668 ( .A(n595), .B(KEYINPUT43), .Z(n597) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n611) );
  NAND2_X1 U670 ( .A1(n615), .A2(n611), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n697), .A2(G210), .ZN(n606) );
  XOR2_X1 U672 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n603) );
  XNOR2_X1 U673 ( .A(KEYINPUT88), .B(KEYINPUT83), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n601), .B(n604), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n606), .B(n605), .ZN(n608) );
  INV_X1 U677 ( .A(G952), .ZN(n607) );
  NOR2_X2 U678 ( .A1(n608), .A2(n709), .ZN(n610) );
  XNOR2_X1 U679 ( .A(KEYINPUT124), .B(KEYINPUT56), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n610), .B(n609), .ZN(G51) );
  XNOR2_X1 U681 ( .A(n611), .B(G140), .ZN(G42) );
  XNOR2_X1 U682 ( .A(G128), .B(KEYINPUT29), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n613), .B(n612), .ZN(G30) );
  XNOR2_X1 U684 ( .A(n614), .B(G137), .ZN(G39) );
  XNOR2_X1 U685 ( .A(n615), .B(G134), .ZN(G36) );
  XNOR2_X1 U686 ( .A(n616), .B(G131), .ZN(G33) );
  XOR2_X1 U687 ( .A(G146), .B(KEYINPUT118), .Z(n618) );
  XNOR2_X1 U688 ( .A(n617), .B(n618), .ZN(G48) );
  XNOR2_X1 U689 ( .A(G119), .B(KEYINPUT127), .ZN(n620) );
  XOR2_X1 U690 ( .A(n620), .B(n619), .Z(G21) );
  NAND2_X1 U691 ( .A1(n697), .A2(G472), .ZN(n624) );
  XOR2_X1 U692 ( .A(KEYINPUT115), .B(KEYINPUT62), .Z(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n624), .B(n623), .ZN(n625) );
  NOR2_X2 U695 ( .A1(n625), .A2(n709), .ZN(n627) );
  XOR2_X1 U696 ( .A(KEYINPUT116), .B(KEYINPUT63), .Z(n626) );
  XNOR2_X1 U697 ( .A(n627), .B(n626), .ZN(G57) );
  XNOR2_X1 U698 ( .A(n628), .B(G122), .ZN(G24) );
  NAND2_X1 U699 ( .A1(n350), .A2(G469), .ZN(n632) );
  XOR2_X1 U700 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n630) );
  XNOR2_X1 U701 ( .A(n629), .B(n630), .ZN(n631) );
  XNOR2_X1 U702 ( .A(n632), .B(n631), .ZN(n633) );
  NOR2_X1 U703 ( .A1(n633), .A2(n709), .ZN(G54) );
  XNOR2_X1 U704 ( .A(G101), .B(n634), .ZN(G3) );
  NOR2_X1 U705 ( .A1(n645), .A2(n636), .ZN(n635) );
  XOR2_X1 U706 ( .A(G104), .B(n635), .Z(G6) );
  NOR2_X1 U707 ( .A1(n648), .A2(n636), .ZN(n638) );
  XNOR2_X1 U708 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(G107), .B(n639), .ZN(G9) );
  XOR2_X1 U711 ( .A(G110), .B(n641), .Z(G12) );
  XOR2_X1 U712 ( .A(G143), .B(KEYINPUT117), .Z(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(G45) );
  NOR2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n647) );
  XNOR2_X1 U715 ( .A(G113), .B(KEYINPUT119), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(G15) );
  NOR2_X1 U717 ( .A1(n648), .A2(n644), .ZN(n649) );
  XOR2_X1 U718 ( .A(G116), .B(n649), .Z(G18) );
  XNOR2_X1 U719 ( .A(G125), .B(n650), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U721 ( .A1(n351), .A2(KEYINPUT84), .ZN(n654) );
  INV_X1 U722 ( .A(n690), .ZN(n665) );
  AND2_X1 U723 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n663) );
  NOR2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U726 ( .A(KEYINPUT121), .B(n661), .Z(n662) );
  NOR2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U728 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U729 ( .A(KEYINPUT122), .B(n666), .Z(n683) );
  NAND2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U731 ( .A(KEYINPUT120), .B(n670), .Z(n671) );
  XNOR2_X1 U732 ( .A(n671), .B(KEYINPUT49), .ZN(n674) );
  INV_X1 U733 ( .A(n672), .ZN(n673) );
  AND2_X1 U734 ( .A1(n674), .A2(n673), .ZN(n678) );
  NAND2_X1 U735 ( .A1(n675), .A2(n498), .ZN(n676) );
  XNOR2_X1 U736 ( .A(n676), .B(KEYINPUT50), .ZN(n677) );
  NAND2_X1 U737 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U738 ( .A1(n667), .A2(n679), .ZN(n680) );
  XOR2_X1 U739 ( .A(KEYINPUT51), .B(n680), .Z(n681) );
  NAND2_X1 U740 ( .A1(n681), .A2(n691), .ZN(n682) );
  NAND2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U742 ( .A(KEYINPUT52), .B(n684), .ZN(n685) );
  NAND2_X1 U743 ( .A1(n685), .A2(G952), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n689), .A2(n688), .ZN(n694) );
  NAND2_X1 U746 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U747 ( .A(KEYINPUT123), .B(n692), .Z(n693) );
  NAND2_X1 U748 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n696), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U750 ( .A1(n697), .A2(G475), .ZN(n700) );
  XOR2_X1 U751 ( .A(n698), .B(KEYINPUT59), .Z(n699) );
  XNOR2_X1 U752 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X2 U753 ( .A1(n701), .A2(n709), .ZN(n702) );
  XNOR2_X1 U754 ( .A(n702), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U755 ( .A1(n350), .A2(G478), .ZN(n704) );
  XNOR2_X1 U756 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U757 ( .A1(n709), .A2(n705), .ZN(G63) );
  NAND2_X1 U758 ( .A1(n350), .A2(G217), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(G66) );
  AND2_X1 U761 ( .A1(n710), .A2(n726), .ZN(n714) );
  INV_X1 U762 ( .A(G898), .ZN(n715) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n711) );
  XOR2_X1 U764 ( .A(KEYINPUT61), .B(n711), .Z(n712) );
  NOR2_X1 U765 ( .A1(n715), .A2(n712), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n722) );
  NAND2_X1 U767 ( .A1(n715), .A2(G953), .ZN(n719) );
  XOR2_X1 U768 ( .A(G101), .B(KEYINPUT126), .Z(n716) );
  XNOR2_X1 U769 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U770 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n720), .B(KEYINPUT125), .ZN(n721) );
  XOR2_X1 U772 ( .A(n722), .B(n721), .Z(G69) );
  XOR2_X1 U773 ( .A(n724), .B(n723), .Z(n728) );
  XNOR2_X1 U774 ( .A(n725), .B(n728), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(n726), .ZN(n732) );
  XOR2_X1 U776 ( .A(n728), .B(G227), .Z(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G900), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n730), .A2(G953), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n732), .A2(n731), .ZN(G72) );
endmodule

