//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G116), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT67), .A3(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n194), .A2(new_n195), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n194), .B2(new_n195), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n192), .A2(KEYINPUT67), .A3(G119), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT67), .B1(new_n192), .B2(G119), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n195), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n200), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n194), .A2(new_n195), .A3(new_n200), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT68), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT82), .B(G101), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G104), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n218), .A3(new_n215), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n219), .A2(KEYINPUT4), .B1(G101), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(KEYINPUT4), .A3(G101), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI22_X1  g037(.A1(new_n204), .A2(new_n211), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT87), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT83), .ZN(new_n226));
  XNOR2_X1  g040(.A(G104), .B(G107), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n217), .A2(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n215), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT83), .A3(G101), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n229), .A2(new_n219), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(new_n196), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT5), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n207), .B2(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n233), .A2(new_n210), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n203), .B1(new_n201), .B2(new_n202), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n209), .A2(KEYINPUT68), .A3(new_n210), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n219), .A2(KEYINPUT4), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n220), .A2(G101), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n222), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n243), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G110), .B(G122), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n225), .A2(new_n239), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT89), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n240), .A2(new_n241), .B1(new_n246), .B2(new_n222), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n238), .B1(new_n252), .B2(new_n243), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT89), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n225), .A3(new_n254), .A4(new_n249), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n249), .B(KEYINPUT8), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n233), .B1(new_n210), .B2(new_n237), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n238), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n260));
  INV_X1    g074(.A(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G143), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n266), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G125), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n260), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n261), .A2(G143), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n265), .A2(new_n275), .B1(KEYINPUT1), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n275), .A2(KEYINPUT1), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT66), .B1(new_n270), .B2(new_n278), .ZN(new_n279));
  AND4_X1   g093(.A1(KEYINPUT66), .A2(new_n278), .A3(new_n262), .A4(new_n264), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n273), .B(new_n277), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n269), .A2(KEYINPUT90), .A3(G125), .A4(new_n271), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n274), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G224), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n283), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT91), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT7), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n289), .B2(new_n286), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n274), .A2(new_n281), .A3(new_n282), .A4(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT92), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n259), .B(new_n288), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n256), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(KEYINPUT93), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT93), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n296), .B1(new_n251), .B2(new_n255), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n248), .A2(new_n239), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n252), .A2(new_n243), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n253), .A2(KEYINPUT88), .A3(new_n225), .ZN(new_n309));
  INV_X1    g123(.A(new_n249), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT6), .A4(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT6), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n251), .B2(new_n255), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n283), .B(new_n286), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n304), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G210), .B1(G237), .B2(G902), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n304), .A2(new_n318), .A3(new_n320), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n188), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G113), .B(G122), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(new_n213), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n273), .A2(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n273), .A2(KEYINPUT16), .A3(G140), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n330), .A2(G146), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT19), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT94), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n335), .A2(KEYINPUT94), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n339), .B(new_n261), .C1(new_n334), .C2(new_n337), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT69), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G953), .ZN(new_n343));
  INV_X1    g157(.A(G237), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n341), .A2(new_n343), .A3(G214), .A4(new_n344), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n345), .A2(new_n263), .ZN(new_n346));
  INV_X1    g160(.A(G131), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n263), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n333), .B(new_n340), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n346), .A2(new_n348), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT18), .A3(G131), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n334), .B(new_n261), .ZN(new_n355));
  NAND2_X1  g169(.A1(KEYINPUT18), .A2(G131), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n348), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n326), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(G146), .B1(new_n330), .B2(new_n331), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n360), .B(new_n332), .C1(new_n351), .C2(KEYINPUT17), .ZN(new_n361));
  INV_X1    g175(.A(new_n351), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT17), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n349), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n357), .A2(new_n355), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n361), .A2(new_n364), .B1(new_n354), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n359), .B1(new_n366), .B2(new_n326), .ZN(new_n367));
  NOR2_X1   g181(.A1(G475), .A2(G902), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n368), .B(KEYINPUT95), .Z(new_n369));
  OR2_X1    g183(.A1(new_n369), .A2(KEYINPUT96), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(KEYINPUT96), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT97), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT20), .B1(new_n367), .B2(new_n369), .ZN(new_n376));
  INV_X1    g190(.A(new_n359), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n332), .A2(new_n360), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n362), .B2(new_n363), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT17), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n326), .B(new_n358), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT97), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n373), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n375), .A2(new_n376), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n366), .A2(new_n326), .ZN(new_n386));
  INV_X1    g200(.A(new_n381), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n299), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G475), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n263), .A2(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n275), .A2(G143), .ZN(new_n393));
  INV_X1    g207(.A(G134), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G116), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n192), .A2(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n398), .A3(new_n217), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT13), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n392), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n393), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n392), .A2(new_n403), .ZN(new_n406));
  OAI21_X1  g220(.A(G134), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n192), .A2(KEYINPUT14), .A3(G122), .ZN(new_n409));
  OAI211_X1 g223(.A(G107), .B(new_n409), .C1(new_n399), .C2(KEYINPUT14), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n394), .B1(new_n392), .B2(new_n393), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n410), .B(new_n401), .C1(new_n395), .C2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT9), .B(G234), .ZN(new_n413));
  INV_X1    g227(.A(G217), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n413), .A2(new_n414), .A3(G953), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n408), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n408), .B2(new_n412), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT98), .A3(new_n299), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G478), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n420), .A2(KEYINPUT15), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(KEYINPUT15), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n341), .A2(new_n343), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n299), .B(new_n425), .C1(G234), .C2(G237), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(G898), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G952), .ZN(new_n429));
  AOI211_X1 g243(.A(G953), .B(new_n429), .C1(G234), .C2(G237), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n432), .B(KEYINPUT99), .Z(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n424), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G221), .B1(new_n413), .B2(G902), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT80), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n233), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n276), .A2(KEYINPUT1), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n270), .B2(G128), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n270), .A2(new_n278), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n270), .A2(KEYINPUT66), .A3(new_n278), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n229), .A2(new_n219), .A3(new_n232), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(KEYINPUT86), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n233), .A2(new_n439), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G137), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G134), .ZN(new_n453));
  AND2_X1   g267(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n454));
  NOR2_X1   g268(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT65), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n453), .B(KEYINPUT65), .C1(new_n454), .C2(new_n455), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n452), .A2(KEYINPUT11), .A3(G134), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n394), .A2(G137), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G131), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n458), .A2(new_n347), .A3(new_n459), .A4(new_n463), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT85), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n451), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT12), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n439), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n233), .A2(new_n439), .A3(KEYINPUT84), .A4(KEYINPUT10), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n466), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n462), .B1(new_n456), .B2(new_n457), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n347), .B1(new_n476), .B2(new_n459), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT10), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n272), .A2(new_n247), .B1(new_n450), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT12), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n451), .A2(new_n482), .A3(new_n467), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n469), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n425), .A2(G227), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT81), .ZN(new_n486));
  XNOR2_X1  g300(.A(G110), .B(G140), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n479), .B1(new_n447), .B2(new_n448), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n272), .B1(new_n221), .B2(new_n223), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n472), .B2(new_n473), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n488), .B1(new_n493), .B2(new_n478), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n474), .A2(new_n480), .ZN(new_n495));
  INV_X1    g309(.A(new_n478), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(new_n498), .A3(G469), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(new_n299), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n478), .B1(new_n474), .B2(new_n480), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n488), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n488), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n469), .A2(new_n481), .A3(new_n507), .A4(new_n483), .ZN(new_n508));
  AOI21_X1  g322(.A(G902), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n500), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n437), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n324), .A2(new_n391), .A3(new_n435), .A4(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n513));
  NOR2_X1   g327(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n514));
  OAI211_X1 g328(.A(G119), .B(new_n275), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G110), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n190), .A2(G128), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n190), .B2(G128), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n515), .A2(new_n516), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n275), .A2(G119), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n517), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT24), .B(G110), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT76), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT76), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n334), .A2(new_n261), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n332), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n514), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n521), .B1(new_n532), .B2(new_n518), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n519), .A2(new_n517), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT75), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT75), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n515), .A2(new_n536), .A3(new_n517), .A4(new_n519), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n535), .A2(G110), .A3(new_n537), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n332), .A2(new_n360), .B1(new_n522), .B2(new_n523), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n531), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n425), .A2(G221), .A3(G234), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT22), .B(G137), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n531), .B(new_n543), .C1(new_n538), .C2(new_n539), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G234), .ZN(new_n548));
  OAI21_X1  g362(.A(G217), .B1(new_n548), .B2(G902), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n299), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT78), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n299), .A3(new_n546), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT77), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT25), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n465), .A2(new_n466), .B1(new_n269), .B2(new_n271), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n453), .A2(new_n461), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G131), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n439), .A2(new_n466), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n242), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n204), .A2(new_n211), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n272), .B1(new_n475), .B2(new_n477), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n439), .A2(new_n466), .A3(new_n564), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT28), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT28), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n425), .A2(G210), .A3(new_n344), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT27), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT26), .B(G101), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n572), .A2(KEYINPUT71), .A3(new_n574), .A4(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT29), .ZN(new_n580));
  INV_X1    g394(.A(new_n578), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT30), .B1(new_n562), .B2(new_n565), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT30), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n568), .A2(new_n583), .A3(new_n569), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n567), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n562), .A2(new_n565), .A3(new_n242), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n579), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n574), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n573), .B1(new_n566), .B2(new_n570), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT71), .B1(new_n591), .B2(new_n578), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n561), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT71), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n572), .A2(new_n574), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n581), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n582), .A2(new_n584), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n242), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n570), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT29), .B1(new_n599), .B2(new_n581), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n596), .A2(new_n600), .A3(KEYINPUT72), .A4(new_n579), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n590), .A2(KEYINPUT73), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n595), .B2(KEYINPUT73), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n581), .A2(new_n580), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n593), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n606), .A2(G472), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n595), .A2(new_n581), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT70), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n598), .A2(new_n609), .A3(new_n570), .A4(new_n578), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT31), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n585), .A2(new_n581), .A3(new_n586), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT31), .B1(new_n613), .B2(new_n609), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n608), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(G472), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(KEYINPUT32), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT32), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n610), .A2(new_n611), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n585), .A2(new_n586), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n620), .A2(new_n609), .A3(KEYINPUT31), .A4(new_n578), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n619), .A2(new_n621), .B1(new_n595), .B2(new_n581), .ZN(new_n622));
  INV_X1    g436(.A(new_n616), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n560), .B1(new_n607), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT79), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n606), .A2(G472), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n624), .A3(new_n617), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT79), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n560), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n512), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n212), .ZN(G3));
  OAI21_X1  g447(.A(KEYINPUT101), .B1(new_n416), .B2(new_n417), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n421), .A2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n418), .A2(new_n299), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n636), .A2(new_n637), .B1(new_n638), .B2(new_n421), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n391), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n324), .A2(new_n433), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n622), .B2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n615), .A2(new_n616), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n437), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n499), .A2(new_n502), .ZN(new_n647));
  AOI211_X1 g461(.A(G469), .B(G902), .C1(new_n506), .C2(new_n508), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n560), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n642), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n649), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n651), .A2(KEYINPUT100), .A3(new_n644), .A4(new_n643), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n641), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT34), .B(G104), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  INV_X1    g470(.A(new_n424), .ZN(new_n657));
  INV_X1    g471(.A(new_n376), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n367), .A2(KEYINPUT20), .A3(new_n369), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n389), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n324), .A2(new_n433), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n653), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT35), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  INV_X1    g479(.A(new_n645), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n558), .A2(new_n559), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT36), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n543), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n540), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n540), .A2(new_n669), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n671), .A3(new_n552), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n391), .A2(new_n673), .A3(new_n435), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n324), .A2(new_n511), .A3(new_n666), .A4(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  NAND2_X1  g491(.A1(new_n511), .A2(new_n673), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n617), .A2(new_n624), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n679), .B2(new_n628), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n426), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n431), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n657), .A2(new_n660), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT102), .B1(new_n324), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n304), .A2(new_n320), .A3(new_n318), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n320), .B1(new_n304), .B2(new_n318), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n187), .B(new_n685), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n680), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XOR2_X1   g507(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n683), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n511), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n698));
  NOR4_X1   g512(.A1(new_n697), .A2(new_n698), .A3(new_n188), .A4(new_n673), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n581), .A2(new_n571), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n299), .B1(new_n702), .B2(new_n613), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G472), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n617), .A2(new_n624), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n391), .A2(new_n657), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n322), .A2(new_n323), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT38), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n699), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT105), .B(G143), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G45));
  NAND2_X1  g526(.A1(new_n636), .A2(new_n637), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n638), .A2(new_n421), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n390), .A2(new_n715), .A3(new_n683), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n188), .B(new_n716), .C1(new_n322), .C2(new_n323), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n680), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  INV_X1    g533(.A(new_n436), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n509), .B2(new_n500), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n497), .A2(new_n481), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n451), .A2(new_n482), .A3(new_n467), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n482), .B1(new_n451), .B2(new_n467), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n723), .A2(new_n488), .B1(new_n494), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(G469), .B1(new_n727), .B2(G902), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n722), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n721), .B(G469), .C1(new_n727), .C2(G902), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n720), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n629), .A2(new_n560), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n641), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT41), .B(G113), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NOR2_X1   g549(.A1(new_n662), .A2(new_n732), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n192), .ZN(G18));
  NAND4_X1  g551(.A1(new_n324), .A2(new_n629), .A3(new_n674), .A4(new_n731), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  OAI22_X1  g553(.A1(new_n612), .A2(new_n614), .B1(new_n603), .B2(new_n578), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n616), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n643), .A2(new_n741), .A3(new_n560), .ZN(new_n742));
  AOI211_X1 g556(.A(new_n434), .B(new_n720), .C1(new_n729), .C2(new_n730), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n324), .A2(new_n742), .A3(new_n706), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  OAI211_X1 g559(.A(new_n731), .B(new_n187), .C1(new_n687), .C2(new_n688), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n639), .B(new_n684), .C1(new_n385), .C2(new_n389), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n643), .A3(new_n673), .A4(new_n741), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT107), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n748), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n324), .A3(new_n751), .A4(new_n731), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  OR2_X1    g568(.A1(new_n624), .A2(KEYINPUT108), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n624), .A2(KEYINPUT108), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n628), .A3(new_n756), .A4(new_n617), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n720), .B1(new_n503), .B2(new_n510), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n322), .A2(new_n187), .A3(new_n758), .A4(new_n323), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n757), .A2(new_n760), .A3(new_n560), .A4(new_n747), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n626), .A2(new_n759), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n761), .A2(KEYINPUT42), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n760), .A2(new_n629), .A3(new_n560), .A4(new_n685), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  AOI21_X1  g581(.A(KEYINPUT43), .B1(new_n715), .B2(KEYINPUT109), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(KEYINPUT109), .B2(new_n715), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n390), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n639), .B1(new_n390), .B2(KEYINPUT110), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(KEYINPUT110), .B2(new_n390), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n770), .B1(new_n772), .B2(KEYINPUT43), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n645), .A3(new_n673), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT44), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n687), .A2(new_n688), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n187), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n489), .A2(new_n498), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT45), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n780), .B2(KEYINPUT45), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n502), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n648), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n436), .A3(new_n695), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n779), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n775), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n436), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT47), .ZN(new_n792));
  OR4_X1    g606(.A1(new_n629), .A2(new_n777), .A3(new_n560), .A4(new_n716), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT112), .B(G140), .Z(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G42));
  NAND2_X1  g610(.A1(new_n729), .A2(new_n730), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT49), .Z(new_n798));
  NAND3_X1  g612(.A1(new_n560), .A2(new_n187), .A3(new_n646), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n798), .A2(new_n772), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n705), .ZN(new_n801));
  INV_X1    g615(.A(new_n709), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n773), .A2(new_n430), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n742), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n746), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n731), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n777), .A2(new_n809), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n560), .A2(new_n810), .A3(new_n430), .A4(new_n801), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n429), .B(G953), .C1(new_n811), .C2(new_n640), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n808), .A2(KEYINPUT119), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT119), .B1(new_n808), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n731), .A2(new_n188), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT117), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n816), .A2(KEYINPUT117), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n802), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT50), .B1(new_n819), .B2(new_n805), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n804), .A2(new_n810), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n643), .A2(new_n741), .A3(new_n673), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n811), .A2(new_n391), .A3(new_n639), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n797), .A2(new_n437), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n792), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n779), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n819), .A2(KEYINPUT50), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(KEYINPUT51), .B(new_n826), .C1(new_n832), .C2(new_n805), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n805), .B1(new_n830), .B2(new_n831), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(new_n825), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n757), .A2(new_n560), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n821), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT48), .B1(new_n838), .B2(KEYINPUT120), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(KEYINPUT120), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n815), .A2(new_n833), .A3(new_n836), .A4(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n187), .B1(new_n687), .B2(new_n688), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n672), .B(new_n684), .C1(new_n558), .C2(new_n559), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n844), .B(new_n436), .C1(new_n647), .C2(new_n648), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT114), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n510), .A2(new_n502), .A3(new_n499), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n436), .A4(new_n844), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n851), .A2(new_n707), .B1(new_n717), .B2(new_n680), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n692), .A2(new_n852), .A3(new_n753), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n689), .A2(new_n690), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n708), .A2(KEYINPUT102), .A3(new_n187), .A4(new_n685), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n857), .A2(new_n680), .B1(new_n749), .B2(new_n752), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n852), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n675), .A2(new_n738), .A3(new_n744), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n632), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n660), .A2(new_n424), .A3(new_n684), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n776), .A2(new_n864), .A3(new_n187), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n322), .A2(new_n187), .A3(new_n323), .A4(new_n865), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT113), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n868), .A3(new_n680), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n760), .A2(new_n750), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n869), .A2(new_n766), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n732), .B1(new_n641), .B2(new_n662), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n390), .A2(new_n715), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n390), .B2(new_n657), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n324), .A2(new_n433), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n653), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n863), .A2(new_n871), .A3(new_n877), .A4(new_n764), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n861), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n859), .B1(new_n858), .B2(new_n852), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n859), .A2(new_n692), .A3(new_n753), .A4(new_n852), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT115), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n854), .A2(new_n860), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n878), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n880), .B1(new_n887), .B2(new_n879), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n879), .B1(new_n861), .B2(new_n878), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n887), .B2(new_n879), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT116), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n895), .A3(KEYINPUT54), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n842), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n803), .B1(new_n897), .B2(new_n898), .ZN(G75));
  NAND2_X1  g713(.A1(new_n887), .A2(new_n879), .ZN(new_n900));
  INV_X1    g714(.A(new_n880), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(G210), .A3(G902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n315), .B(new_n316), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n425), .A2(G952), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(G51));
  XNOR2_X1  g724(.A(new_n501), .B(KEYINPUT57), .ZN(new_n911));
  AOI211_X1 g725(.A(KEYINPUT54), .B(new_n880), .C1(new_n879), .C2(new_n887), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n889), .B1(new_n900), .B2(new_n901), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n727), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR4_X1    g730(.A1(new_n299), .A2(new_n888), .A3(new_n781), .A4(new_n782), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n909), .B1(new_n916), .B2(new_n917), .ZN(G54));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT121), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n902), .A2(G902), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n921), .A2(new_n367), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n367), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n909), .ZN(G60));
  INV_X1    g738(.A(new_n636), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n912), .B2(new_n913), .ZN(new_n929));
  INV_X1    g743(.A(new_n909), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n927), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n894), .A2(new_n896), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n925), .B2(new_n933), .ZN(G63));
  NOR2_X1   g748(.A1(new_n670), .A2(new_n671), .ZN(new_n935));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT122), .Z(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n902), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n938), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n547), .B1(new_n888), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n930), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n939), .A2(new_n941), .A3(KEYINPUT61), .A4(new_n930), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(G66));
  NAND2_X1  g760(.A1(new_n863), .A2(new_n877), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n425), .ZN(new_n948));
  INV_X1    g762(.A(G224), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n427), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n315), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(G898), .B2(new_n425), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(G69));
  XNOR2_X1  g768(.A(new_n874), .B(KEYINPUT123), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n955), .A2(new_n777), .A3(new_n696), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n627), .A2(new_n631), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT124), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n959), .A2(new_n794), .A3(new_n789), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n858), .A2(new_n718), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n710), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n339), .B1(new_n334), .B2(new_n337), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n597), .B(new_n966), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n425), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n425), .A2(G900), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT125), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n324), .A2(new_n706), .ZN(new_n972));
  OR3_X1    g786(.A1(new_n787), .A2(new_n972), .A3(new_n837), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n973), .A2(new_n764), .A3(new_n766), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n794), .A2(new_n974), .A3(new_n789), .A4(new_n961), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n971), .B1(new_n975), .B2(new_n425), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n969), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n425), .B1(G227), .B2(G900), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n981), .B(new_n969), .C1(new_n978), .C2(new_n979), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(G72));
  XOR2_X1   g799(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n986));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n965), .B2(new_n947), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n989), .A2(new_n578), .A3(new_n599), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n620), .A2(new_n578), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n892), .B(new_n988), .C1(new_n991), .C2(new_n613), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n988), .B1(new_n975), .B2(new_n947), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n599), .A2(new_n578), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n909), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n990), .A2(new_n992), .A3(new_n995), .ZN(G57));
endmodule


