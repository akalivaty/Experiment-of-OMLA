//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G20), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n211), .B1(KEYINPUT1), .B2(new_n223), .C1(new_n225), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(KEYINPUT64), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND2_X1  g0048(.A1(new_n227), .A2(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n206), .A2(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NOR3_X1   g0052(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n249), .B1(new_n202), .B2(new_n250), .C1(new_n254), .C2(new_n218), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G1), .A2(G13), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n255), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G68), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT12), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n261), .B(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n256), .A2(new_n257), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G1), .B2(new_n206), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n259), .B(new_n263), .C1(new_n227), .C2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT11), .B1(new_n255), .B2(new_n258), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT14), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT13), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n220), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G226), .A2(G1698), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n235), .B2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n273), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n274), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n272), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n219), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n235), .A2(G1698), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n286), .B(new_n287), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n274), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n257), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(KEYINPUT69), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n283), .A2(G238), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT65), .ZN(new_n299));
  OAI21_X1  g0099(.A(G274), .B1(new_n293), .B2(new_n257), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n297), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n224), .B2(new_n282), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  AOI21_X1  g0105(.A(G1), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(KEYINPUT65), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n298), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n271), .B1(new_n296), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT69), .B1(new_n292), .B2(new_n294), .ZN(new_n310));
  AOI211_X1 g0110(.A(new_n272), .B(new_n283), .C1(new_n290), .C2(new_n291), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n271), .B(new_n308), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n270), .B(G169), .C1(new_n309), .C2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(G179), .A3(new_n312), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n312), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n270), .B1(new_n319), .B2(G169), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n269), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(G200), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(new_n268), .C1(new_n323), .C2(new_n319), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n285), .A2(G222), .ZN(new_n326));
  AND2_X1   g0126(.A1(G223), .A2(G1698), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n280), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n202), .B2(new_n280), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT66), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n283), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n330), .B2(new_n329), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n301), .A2(new_n307), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n294), .A2(new_n306), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(G226), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G200), .ZN(new_n338));
  MUX2_X1   g0138(.A(new_n260), .B(new_n265), .S(G50), .Z(new_n339));
  INV_X1    g0139(.A(G150), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n254), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n342), .A2(new_n250), .B1(new_n206), .B2(new_n201), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n258), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT9), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n332), .A2(G190), .A3(new_n336), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n338), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n348), .B(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n345), .B1(new_n337), .B2(G179), .ZN(new_n351));
  INV_X1    g0151(.A(G169), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n337), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n260), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n342), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n265), .B2(new_n342), .ZN(new_n357));
  XOR2_X1   g0157(.A(new_n357), .B(KEYINPUT73), .Z(new_n358));
  NOR2_X1   g0158(.A1(new_n288), .A2(new_n289), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n359), .B2(new_n206), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n279), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT70), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n278), .A2(new_n206), .A3(new_n279), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n361), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT70), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(G68), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G58), .A2(G68), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(G58), .A2(G68), .ZN(new_n375));
  OAI21_X1  g0175(.A(G20), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n372), .B(new_n376), .C1(new_n254), .C2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT67), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(new_n206), .A3(new_n273), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n380), .B2(new_n251), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n206), .B1(new_n228), .B2(new_n373), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT71), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n264), .B1(new_n371), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT72), .B1(new_n360), .B2(new_n362), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT72), .B1(new_n365), .B2(new_n366), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n227), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n378), .A2(new_n383), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n358), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n219), .A2(G1698), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(G223), .B2(G1698), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n396), .A2(new_n359), .B1(new_n273), .B2(new_n214), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n294), .B1(G232), .B2(new_n335), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n333), .ZN(new_n399));
  INV_X1    g0199(.A(G179), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n352), .B1(new_n398), .B2(new_n333), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT18), .B1(new_n394), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n357), .B(KEYINPUT73), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n369), .B1(new_n368), .B2(G68), .ZN(new_n406));
  AOI211_X1 g0206(.A(KEYINPUT70), .B(new_n227), .C1(new_n367), .C2(new_n361), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n258), .B1(new_n408), .B2(new_n384), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT72), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n367), .B2(new_n361), .ZN(new_n411));
  OAI21_X1  g0211(.A(G68), .B1(new_n411), .B2(new_n389), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n378), .A2(new_n383), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT16), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n405), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n403), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n413), .B(KEYINPUT16), .C1(new_n407), .C2(new_n406), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n393), .A2(new_n419), .A3(new_n258), .ZN(new_n420));
  INV_X1    g0220(.A(G200), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n399), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT74), .B(G190), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n399), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(new_n405), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(KEYINPUT17), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n394), .B2(new_n424), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n404), .B(new_n418), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n334), .B1(G244), .B2(new_n335), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n280), .A2(KEYINPUT68), .A3(G232), .A4(new_n285), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n359), .A2(new_n235), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n432), .B1(new_n433), .B2(new_n280), .C1(new_n434), .C2(KEYINPUT68), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n280), .A2(G238), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n285), .B1(new_n436), .B2(KEYINPUT68), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n294), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n352), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G20), .A2(G77), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT15), .B(G87), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n441), .B1(new_n250), .B2(new_n442), .C1(new_n254), .C2(new_n342), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n443), .A2(new_n258), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n355), .A2(new_n202), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n265), .B2(new_n202), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n440), .B(new_n448), .C1(G179), .C2(new_n439), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n431), .A2(new_n438), .A3(G190), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n447), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n421), .B1(new_n431), .B2(new_n438), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  AND4_X1   g0255(.A1(new_n325), .A2(new_n354), .A3(new_n430), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(KEYINPUT76), .B2(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n305), .A2(G1), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT76), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(new_n304), .A3(KEYINPUT5), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n303), .A2(new_n458), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n458), .A3(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n283), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(new_n221), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n215), .B1(new_n278), .B2(new_n279), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT75), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(KEYINPUT4), .ZN(new_n468));
  OAI21_X1  g0268(.A(G1698), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(G244), .B1(new_n288), .B2(new_n289), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(new_n468), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n213), .B1(new_n278), .B2(new_n279), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n467), .B1(new_n474), .B2(new_n285), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n469), .B(new_n473), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n465), .B1(new_n477), .B2(new_n294), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT77), .B1(new_n478), .B2(new_n421), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT77), .ZN(new_n480));
  INV_X1    g0280(.A(new_n468), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n470), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(G250), .B1(new_n288), .B2(new_n289), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n285), .B1(new_n483), .B2(new_n481), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(G244), .B(new_n285), .C1(new_n288), .C2(new_n289), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n476), .B1(new_n486), .B2(KEYINPUT75), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n283), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n480), .B(G200), .C1(new_n489), .C2(new_n465), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n479), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n433), .B1(new_n388), .B2(new_n390), .ZN(new_n492));
  XNOR2_X1  g0292(.A(G97), .B(G107), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n433), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n497), .A2(new_n206), .B1(new_n202), .B2(new_n254), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n258), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n260), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n205), .A2(G33), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n264), .A2(new_n260), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n500), .B1(new_n503), .B2(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n469), .A2(new_n473), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n294), .B1(new_n505), .B2(new_n487), .ZN(new_n506));
  INV_X1    g0306(.A(new_n465), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(G190), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n499), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n506), .A2(new_n400), .A3(new_n507), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(G169), .B2(new_n478), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n499), .A2(new_n504), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n491), .A2(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n214), .A2(new_n220), .A3(new_n433), .ZN(new_n516));
  OAI211_X1 g0316(.A(KEYINPUT19), .B(new_n516), .C1(new_n274), .C2(G20), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n206), .B(G68), .C1(new_n288), .C2(new_n289), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT19), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n250), .B2(new_n220), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT79), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n517), .A2(KEYINPUT79), .A3(new_n518), .A4(new_n520), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n258), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n442), .A2(new_n355), .ZN(new_n526));
  INV_X1    g0326(.A(new_n442), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n503), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n215), .B1(new_n305), .B2(G1), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n205), .A2(new_n302), .A3(G45), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n283), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(G238), .B(new_n285), .C1(new_n288), .C2(new_n289), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G116), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n535), .C1(new_n472), .C2(new_n285), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n536), .B2(new_n294), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n400), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT78), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n537), .A2(G169), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT78), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n537), .A2(new_n541), .A3(new_n400), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n529), .A2(new_n539), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n264), .B1(new_n521), .B2(new_n522), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n524), .B1(new_n355), .B2(new_n442), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n503), .A2(G87), .ZN(new_n546));
  AOI211_X1 g0346(.A(G190), .B(new_n533), .C1(new_n536), .C2(new_n294), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n536), .A2(new_n294), .ZN(new_n548));
  AOI21_X1  g0348(.A(G200), .B1(new_n548), .B2(new_n532), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n221), .A2(new_n285), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n288), .B2(new_n289), .ZN(new_n553));
  OAI211_X1 g0353(.A(G250), .B(new_n285), .C1(new_n288), .C2(new_n289), .ZN(new_n554));
  INV_X1    g0354(.A(G294), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n273), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n294), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n463), .A2(G264), .A3(new_n283), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n559), .A2(G179), .A3(new_n462), .A4(new_n560), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n559), .A2(new_n462), .A3(new_n560), .ZN(new_n563));
  AOI22_X1  g0363(.A1(KEYINPUT83), .A2(new_n561), .B1(new_n563), .B2(G169), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n206), .B(G87), .C1(new_n288), .C2(new_n289), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n280), .A2(new_n206), .A3(G87), .A4(new_n567), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n535), .B2(G20), .ZN(new_n575));
  OR3_X1    g0375(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n206), .A2(KEYINPUT82), .A3(G33), .A4(G116), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n578));
  AND4_X1   g0378(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n572), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n573), .B1(new_n572), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n258), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT25), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n260), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n433), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n503), .A2(G107), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n562), .A2(new_n564), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n559), .A2(new_n323), .A3(new_n462), .A4(new_n560), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n556), .B1(new_n280), .B2(new_n552), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n283), .B1(new_n589), .B2(new_n554), .ZN(new_n590));
  INV_X1    g0390(.A(new_n462), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n463), .A2(G264), .A3(new_n283), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n588), .B1(new_n593), .B2(G200), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n582), .A2(new_n594), .A3(new_n586), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n260), .A2(G116), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G116), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n502), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(G20), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n258), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(G20), .B1(G33), .B2(G283), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n273), .A2(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT80), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT80), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT20), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n470), .B(new_n206), .C1(G33), .C2(new_n220), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT80), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n256), .A2(new_n257), .B1(G20), .B2(new_n598), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n611), .A2(KEYINPUT20), .A3(new_n607), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n600), .B1(new_n608), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G303), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n278), .A2(new_n616), .A3(new_n279), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n285), .A2(G257), .ZN(new_n618));
  NAND2_X1  g0418(.A1(G264), .A2(G1698), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n617), .B(new_n294), .C1(new_n359), .C2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n463), .A2(G270), .A3(new_n283), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n622), .A3(new_n462), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(G169), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n615), .A2(new_n624), .A3(KEYINPUT21), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n611), .A2(new_n607), .A3(new_n612), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n599), .B1(new_n629), .B2(new_n613), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n623), .A2(G169), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n623), .A2(new_n400), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n621), .A2(new_n622), .A3(new_n462), .A4(new_n423), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n623), .A2(G200), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n630), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n625), .A2(new_n632), .A3(new_n634), .A4(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n587), .A2(new_n595), .A3(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n456), .A2(new_n515), .A3(new_n551), .A4(new_n639), .ZN(G372));
  NAND3_X1  g0440(.A1(new_n529), .A2(new_n538), .A3(new_n540), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n352), .B1(new_n489), .B2(new_n465), .ZN(new_n643));
  OAI21_X1  g0443(.A(G107), .B1(new_n411), .B2(new_n389), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n495), .A2(new_n496), .ZN(new_n645));
  INV_X1    g0445(.A(new_n254), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n645), .A2(G20), .B1(new_n646), .B2(G77), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n264), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n504), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n643), .B(new_n511), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n582), .A2(new_n594), .A3(new_n586), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n479), .A2(new_n490), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n509), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n625), .A2(new_n632), .A3(new_n634), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n582), .A2(new_n586), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n564), .A2(new_n562), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n538), .B1(G169), .B2(new_n537), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n549), .A2(new_n547), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n525), .A2(new_n546), .A3(new_n526), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n659), .A2(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT84), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n550), .A2(new_n641), .A3(KEYINPUT84), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n642), .B1(new_n658), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n650), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n551), .A2(KEYINPUT26), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT85), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n644), .A2(new_n647), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n649), .B1(new_n672), .B2(new_n258), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n671), .B1(new_n512), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n514), .A2(KEYINPUT85), .A3(new_n643), .A4(new_n511), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n665), .A2(new_n666), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n670), .B1(new_n676), .B2(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n456), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n404), .A2(new_n418), .ZN(new_n680));
  INV_X1    g0480(.A(new_n321), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n324), .B2(new_n450), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n425), .A2(KEYINPUT17), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n394), .A2(new_n427), .A3(new_n424), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n680), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n350), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n353), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n679), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT86), .Z(G369));
  NAND2_X1  g0491(.A1(new_n656), .A2(new_n655), .ZN(new_n692));
  INV_X1    g0492(.A(G13), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n693), .A2(G1), .A3(G20), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(G213), .B1(new_n695), .B2(KEYINPUT27), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT27), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n694), .A2(KEYINPUT87), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT87), .B1(new_n694), .B2(new_n697), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G343), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n582), .B2(new_n586), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n692), .B(new_n651), .C1(KEYINPUT88), .C2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(KEYINPUT88), .B2(new_n703), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n692), .A2(new_n702), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n630), .A2(new_n702), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n654), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n638), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT89), .Z(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n654), .A2(new_n702), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n705), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n587), .A2(new_n702), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n209), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G1), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n516), .A2(G116), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n725), .A2(new_n726), .B1(new_n229), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n658), .A2(new_n667), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n641), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT26), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n551), .A2(new_n731), .A3(new_n669), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n676), .B2(new_n731), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n702), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .ZN(new_n735));
  INV_X1    g0535(.A(new_n702), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n668), .B2(new_n677), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n735), .B1(KEYINPUT29), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n639), .A2(new_n515), .A3(new_n551), .A4(new_n702), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n537), .A2(new_n560), .A3(new_n559), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n478), .A3(new_n633), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n623), .A2(new_n400), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n593), .A2(new_n745), .A3(new_n537), .ZN(new_n746));
  INV_X1    g0546(.A(new_n478), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n743), .A2(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n742), .A2(new_n478), .A3(KEYINPUT30), .A4(new_n633), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n702), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT31), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n741), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n743), .A2(new_n744), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n746), .A2(new_n747), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n736), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT31), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G330), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n740), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n728), .B1(new_n764), .B2(G1), .ZN(G364));
  AOI21_X1  g0565(.A(new_n257), .B1(G20), .B2(new_n352), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n206), .A2(new_n400), .A3(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n323), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n323), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n206), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G311), .A2(new_n770), .B1(new_n773), .B2(G294), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n423), .A2(new_n768), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n280), .B1(new_n776), .B2(G322), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n206), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n774), .B(new_n777), .C1(new_n616), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n206), .A2(new_n400), .A3(new_n421), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT92), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(KEYINPUT92), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n782), .A2(new_n423), .A3(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT95), .Z(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT96), .B(G326), .Z(new_n787));
  AOI21_X1  g0587(.A(new_n780), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n778), .A2(new_n323), .A3(new_n421), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT93), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT93), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n778), .A2(new_n323), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(G329), .B1(G283), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT97), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n782), .A2(new_n323), .A3(new_n783), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT94), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  OAI211_X1 g0603(.A(new_n788), .B(new_n797), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n779), .A2(new_n214), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n776), .B2(G58), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n806), .B1(new_n202), .B2(new_n769), .C1(new_n433), .C2(new_n794), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n359), .B(new_n807), .C1(G97), .C2(new_n773), .ZN(new_n808));
  INV_X1    g0608(.A(new_n802), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G68), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n793), .A2(G159), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n811), .A2(KEYINPUT32), .ZN(new_n812));
  INV_X1    g0612(.A(new_n784), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n811), .A2(KEYINPUT32), .B1(new_n813), .B2(G50), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n808), .A2(new_n810), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n767), .B1(new_n804), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n693), .A2(G20), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n725), .B1(G45), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n206), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT91), .Z(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n767), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n244), .A2(G45), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n722), .A2(new_n280), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n824), .B(new_n825), .C1(G45), .C2(new_n229), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n722), .A2(new_n359), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(G355), .B1(new_n598), .B2(new_n722), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n823), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n816), .A2(new_n819), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT98), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n710), .A2(new_n822), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n710), .A2(G330), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT90), .Z(new_n835));
  NOR2_X1   g0635(.A1(new_n712), .A2(new_n818), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n359), .B1(new_n220), .B2(new_n772), .C1(new_n792), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n794), .A2(new_n214), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n776), .B2(G294), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n842), .B1(new_n433), .B2(new_n779), .C1(new_n598), .C2(new_n769), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n840), .B(new_n843), .C1(G303), .C2(new_n813), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n802), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT100), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n776), .A2(G143), .B1(new_n770), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n849), .B2(new_n784), .C1(new_n802), .C2(new_n340), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n280), .B1(new_n779), .B2(new_n218), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n772), .A2(new_n226), .B1(new_n794), .B2(new_n227), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(new_n793), .C2(G132), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n766), .B1(new_n847), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n766), .A2(new_n820), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT99), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n818), .C1(G77), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n862));
  INV_X1    g0662(.A(new_n820), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n452), .A2(new_n453), .B1(new_n447), .B2(new_n702), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n449), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n448), .B1(new_n439), .B2(G179), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(new_n440), .A3(new_n702), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n862), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n738), .A2(new_n869), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n737), .A2(new_n870), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n761), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n818), .B1(new_n762), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n873), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G384));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n227), .B2(G50), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n218), .A2(KEYINPUT102), .A3(G68), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n373), .A2(G77), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n882), .B(new_n883), .C1(new_n229), .C2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(G1), .A3(new_n693), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT103), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n598), .B(new_n225), .C1(new_n645), .C2(KEYINPUT35), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(KEYINPUT35), .B2(new_n645), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT36), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n890), .B2(new_n889), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n875), .A2(new_n868), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(new_n425), .ZN(new_n895));
  INV_X1    g0695(.A(new_n701), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n420), .A2(new_n405), .B1(new_n403), .B2(new_n896), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n895), .A2(new_n897), .A3(KEYINPUT37), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n387), .B1(new_n408), .B2(new_n392), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n386), .ZN(new_n900));
  INV_X1    g0700(.A(new_n357), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n701), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n416), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n425), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n898), .B1(KEYINPUT37), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n680), .B2(new_n685), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n894), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n903), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n429), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n357), .B1(new_n899), .B2(new_n386), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n425), .B1(new_n911), .B2(new_n896), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n403), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT37), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n415), .B1(new_n416), .B2(new_n701), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(new_n425), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n918), .A3(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n908), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n268), .A2(new_n702), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n321), .A2(new_n324), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n318), .B2(new_n320), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n893), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n680), .A2(new_n701), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n681), .A2(new_n702), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n919), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n394), .A2(new_n896), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n915), .A2(new_n425), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT37), .B1(new_n897), .B2(KEYINPUT104), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n429), .A2(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n935), .A2(new_n934), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT105), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n429), .A2(new_n933), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n934), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n894), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT105), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n943), .A2(new_n944), .A3(new_n931), .A4(new_n919), .ZN(new_n945));
  INV_X1    g0745(.A(new_n919), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT38), .B1(new_n910), .B2(new_n918), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT39), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n939), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n928), .B1(new_n930), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n739), .A2(new_n456), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n689), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n950), .B(new_n952), .Z(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT106), .B1(new_n750), .B2(KEYINPUT31), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT106), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n756), .A2(new_n955), .A3(new_n757), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n741), .A2(new_n954), .A3(new_n956), .A4(new_n751), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n869), .B1(new_n923), .B2(new_n924), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n920), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT40), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n943), .A2(new_n919), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT40), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n961), .A2(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n456), .A2(new_n957), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n760), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n965), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n953), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n205), .B2(new_n817), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n953), .A2(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n892), .B1(new_n970), .B2(new_n971), .ZN(G367));
  OAI21_X1  g0772(.A(new_n515), .B1(new_n673), .B2(new_n702), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n669), .A2(new_n736), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n714), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n662), .A2(new_n736), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n667), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n641), .B2(new_n978), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT107), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n714), .A2(new_n982), .A3(new_n975), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n977), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n981), .B1(new_n977), .B2(new_n983), .ZN(new_n985));
  INV_X1    g0785(.A(new_n975), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n717), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n973), .A2(new_n692), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n736), .B1(new_n990), .B2(new_n650), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n988), .B2(KEYINPUT42), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n989), .A2(new_n992), .B1(KEYINPUT43), .B2(new_n980), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OR3_X1    g0794(.A1(new_n984), .A2(new_n985), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n984), .B2(new_n985), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n723), .B(KEYINPUT41), .Z(new_n997));
  INV_X1    g0797(.A(KEYINPUT108), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n720), .A2(new_n998), .A3(new_n975), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT108), .B1(new_n719), .B2(new_n986), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n719), .A2(new_n986), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT44), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n715), .B1(new_n1009), .B2(KEYINPUT109), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT109), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1011), .A3(new_n714), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n707), .A2(new_n716), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n705), .B2(new_n716), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(KEYINPUT110), .B2(new_n712), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n711), .B(KEYINPUT110), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n763), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1010), .A2(new_n1012), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n997), .B1(new_n1019), .B2(new_n764), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n205), .B1(new_n817), .B2(G45), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n995), .B(new_n996), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n823), .B1(new_n722), .B2(new_n527), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n825), .A2(new_n239), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n819), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n809), .A2(G159), .B1(G50), .B2(new_n770), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT112), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT112), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n794), .A2(new_n202), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G68), .B2(new_n773), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n226), .B2(new_n779), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n359), .B1(new_n776), .B2(G150), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n792), .B2(new_n849), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(new_n786), .C2(G143), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1028), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G294), .A2(new_n809), .B1(new_n786), .B2(G311), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n779), .A2(new_n598), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT46), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT111), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n359), .B1(new_n769), .B2(new_n845), .C1(new_n1038), .C2(KEYINPUT46), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n773), .A2(G107), .B1(new_n795), .B2(G97), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n616), .B2(new_n775), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(G317), .C2(new_n793), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1037), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1036), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT47), .Z(new_n1047));
  OAI221_X1 g0847(.A(new_n1026), .B1(new_n980), .B2(new_n822), .C1(new_n1047), .C2(new_n767), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1023), .A2(new_n1048), .ZN(G387));
  INV_X1    g0849(.A(new_n1018), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1017), .A2(new_n763), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n723), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n707), .A2(new_n822), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n825), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n342), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n726), .C1(G68), .C2(G77), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n236), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n305), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n827), .A2(new_n726), .B1(new_n433), .B2(new_n722), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT113), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(KEYINPUT113), .A3(new_n1061), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n823), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(G317), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n775), .A2(new_n1066), .B1(new_n769), .B2(new_n616), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT116), .Z(new_n1068));
  INV_X1    g0868(.A(G322), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1068), .B1(new_n785), .B2(new_n1069), .C1(new_n839), .C2(new_n802), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n779), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n773), .A2(G283), .B1(new_n1074), .B2(G294), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT49), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n359), .B1(new_n794), .B2(new_n598), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n793), .B2(new_n787), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1074), .A2(G77), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n792), .B2(new_n340), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT114), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n280), .B1(new_n220), .B2(new_n794), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT115), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n776), .A2(G50), .B1(new_n773), .B2(new_n527), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n227), .B2(new_n769), .C1(new_n377), .C2(new_n784), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n342), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n809), .B2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1077), .A2(new_n1079), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n818), .B1(new_n1062), .B2(new_n1065), .C1(new_n1090), .C2(new_n767), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1053), .B1(new_n1091), .B2(KEYINPUT117), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(KEYINPUT117), .B2(new_n1091), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1052), .B(new_n1093), .C1(new_n1021), .C2(new_n1017), .ZN(G393));
  NOR2_X1   g0894(.A1(new_n1054), .A2(new_n247), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1064), .B1(new_n220), .B2(new_n209), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n818), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n784), .A2(new_n340), .B1(new_n775), .B2(new_n377), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT118), .Z(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n359), .B(new_n841), .C1(new_n793), .C2(G143), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n772), .A2(new_n202), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G68), .B2(new_n1074), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n342), .C2(new_n769), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G50), .B2(new_n809), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n784), .A2(new_n1066), .B1(new_n775), .B2(new_n839), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT52), .Z(new_n1108));
  OAI22_X1  g0908(.A1(new_n769), .A2(new_n555), .B1(new_n772), .B2(new_n598), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n359), .B1(new_n433), .B2(new_n794), .C1(new_n792), .C2(new_n1069), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G283), .C2(new_n1074), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n616), .B2(new_n802), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1106), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1097), .B1(new_n1113), .B2(new_n766), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n975), .B2(new_n822), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1009), .A2(new_n714), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1008), .A2(new_n715), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1115), .B1(new_n1119), .B2(new_n1021), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n724), .B1(new_n1119), .B2(new_n1050), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1019), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(G390));
  INV_X1    g0923(.A(new_n868), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n737), .B2(new_n870), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n925), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n929), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1127), .A2(new_n945), .A3(new_n948), .A4(new_n939), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n865), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n868), .B1(new_n734), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n925), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n930), .B1(new_n943), .B2(new_n919), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n760), .B(new_n869), .C1(new_n752), .C2(new_n758), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n925), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1128), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n869), .A2(new_n760), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n957), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n925), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1136), .B1(new_n1140), .B2(KEYINPUT119), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT119), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1142), .B(new_n1139), .C1(new_n1128), .C2(new_n1133), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n949), .A2(new_n863), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n818), .B1(new_n860), .B2(new_n1088), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n280), .B(new_n805), .C1(new_n793), .C2(G294), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n775), .A2(new_n598), .B1(new_n769), .B2(new_n220), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1102), .B(new_n1148), .C1(G68), .C2(new_n795), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n433), .B2(new_n802), .C1(new_n845), .C2(new_n784), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n802), .A2(new_n849), .ZN(new_n1152));
  XOR2_X1   g0952(.A(KEYINPUT54), .B(G143), .Z(new_n1153));
  AOI22_X1  g0953(.A1(new_n776), .A2(G132), .B1(new_n770), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n218), .B2(new_n794), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G128), .B2(new_n813), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n779), .A2(new_n340), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT53), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n359), .B(new_n1159), .C1(G159), .C2(new_n773), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n793), .A2(G125), .B1(new_n1158), .B2(new_n1157), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1156), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1151), .B1(new_n1152), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1146), .B1(new_n1163), .B2(new_n766), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1144), .A2(new_n1022), .B1(new_n1145), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n456), .A2(G330), .A3(new_n957), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT120), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT120), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n456), .A2(new_n1170), .A3(G330), .A4(new_n957), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(new_n951), .A3(new_n689), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1138), .A2(new_n925), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n925), .B2(new_n1134), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1130), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1139), .B1(new_n1134), .B2(new_n925), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1175), .A2(new_n1176), .B1(new_n893), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1173), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1167), .B1(new_n1144), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(KEYINPUT121), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n724), .B1(new_n1144), .B2(new_n1179), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1166), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G378));
  OAI21_X1  g0986(.A(new_n818), .B1(new_n860), .B2(G50), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n354), .B(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n345), .A2(new_n701), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(new_n863), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n795), .A2(G58), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1080), .A2(new_n1194), .A3(new_n304), .A4(new_n359), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G283), .B2(new_n793), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT122), .Z(new_n1197));
  AOI22_X1  g0997(.A1(new_n776), .A2(G107), .B1(new_n773), .B2(G68), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n442), .B2(new_n769), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G116), .B2(new_n813), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1197), .B(new_n1200), .C1(new_n220), .C2(new_n802), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT123), .Z(new_n1202));
  OR2_X1    g1002(.A1(new_n1202), .A2(KEYINPUT58), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(KEYINPUT58), .ZN(new_n1204));
  AOI21_X1  g1004(.A(G50), .B1(new_n279), .B2(new_n304), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n793), .A2(G124), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n273), .B(new_n304), .C1(new_n794), .C2(new_n377), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n770), .A2(G137), .B1(new_n1074), .B2(new_n1153), .ZN(new_n1208));
  INV_X1    g1008(.A(G128), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n775), .C1(new_n340), .C2(new_n772), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G125), .B2(new_n813), .ZN(new_n1211));
  INV_X1    g1011(.A(G132), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n802), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1206), .B(new_n1207), .C1(new_n1213), .C2(KEYINPUT59), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1205), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1203), .A2(new_n1204), .A3(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1187), .B(new_n1193), .C1(new_n766), .C2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n964), .B1(new_n938), .B2(new_n946), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n959), .B1(new_n919), .B2(new_n908), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(G330), .C1(KEYINPUT40), .C2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT124), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n961), .A2(new_n962), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1224), .A2(KEYINPUT124), .A3(G330), .A4(new_n1219), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1225), .A3(new_n1192), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n965), .A2(new_n1191), .A3(KEYINPUT124), .A4(G330), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1226), .A2(new_n950), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n950), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1218), .B1(new_n1230), .B2(new_n1022), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1173), .B1(new_n1144), .B2(new_n1179), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1229), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1226), .A2(new_n950), .A3(new_n1227), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(KEYINPUT57), .A3(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n723), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n930), .B1(new_n893), .B2(new_n925), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1133), .B1(new_n949), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1139), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1142), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1140), .A2(KEYINPUT119), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(new_n1136), .A4(new_n1179), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1173), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1245), .B2(new_n1230), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1231), .B1(new_n1236), .B2(new_n1246), .ZN(G375));
  INV_X1    g1047(.A(new_n997), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1173), .A2(new_n1178), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1181), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n809), .A2(new_n1153), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n280), .B(new_n1194), .C1(new_n792), .C2(new_n1209), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n770), .A2(G150), .B1(new_n1074), .B2(G159), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n218), .B2(new_n772), .C1(new_n849), .C2(new_n775), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1252), .B(new_n1254), .C1(G132), .C2(new_n813), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1030), .A2(new_n280), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n784), .A2(new_n555), .B1(new_n1256), .B2(KEYINPUT125), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n776), .A2(G283), .B1(new_n770), .B2(G107), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n773), .A2(new_n527), .B1(new_n1074), .B2(G97), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(new_n616), .C2(new_n792), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1257), .B(new_n1260), .C1(KEYINPUT125), .C2(new_n1256), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n809), .A2(G116), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1251), .A2(new_n1255), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n818), .B1(G68), .B2(new_n860), .C1(new_n1263), .C2(new_n767), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1126), .B2(new_n820), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1178), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(new_n1022), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1250), .A2(new_n1267), .ZN(G381));
  NAND3_X1  g1068(.A1(new_n1122), .A2(new_n1023), .A3(new_n1048), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(G375), .ZN(new_n1271));
  NOR4_X1   g1071(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1185), .A4(new_n1272), .ZN(G407));
  INV_X1    g1073(.A(G343), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1271), .A2(G213), .A3(new_n1274), .A4(new_n1185), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(G407), .A2(new_n1275), .A3(G213), .ZN(G409));
  NAND3_X1  g1076(.A1(new_n1245), .A2(new_n1248), .A3(new_n1230), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1231), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1182), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1241), .A2(new_n1242), .A3(new_n1136), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT121), .B1(new_n1280), .B2(new_n1181), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1184), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1278), .A2(new_n1282), .A3(new_n1165), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(G375), .B2(new_n1185), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1274), .A2(G213), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1181), .B(new_n723), .C1(new_n1286), .C2(new_n1249), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT60), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1267), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n879), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G384), .B(new_n1267), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1284), .A2(new_n1285), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1274), .A2(G213), .A3(G2897), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1290), .A2(new_n1296), .A3(new_n1291), .A4(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1290), .A2(new_n1296), .A3(new_n1291), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1297), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1296), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1299), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1295), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT62), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1284), .A2(new_n1306), .A3(new_n1285), .A4(new_n1292), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1294), .A2(new_n1304), .A3(new_n1305), .A4(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1122), .B1(new_n1023), .B2(new_n1048), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(G393), .B(new_n837), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1310), .A2(new_n1269), .A3(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1311), .B1(new_n1270), .B2(new_n1309), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1308), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1315), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1303), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1293), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1285), .A4(new_n1292), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1317), .A2(new_n1318), .A3(new_n1320), .A4(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1316), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT127), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT127), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1316), .A2(new_n1325), .A3(new_n1322), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1326), .ZN(G405));
  XNOR2_X1  g1127(.A(G375), .B(new_n1185), .ZN(new_n1328));
  XOR2_X1   g1128(.A(new_n1328), .B(new_n1292), .Z(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(new_n1317), .ZN(G402));
endmodule


