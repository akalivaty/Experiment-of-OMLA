

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U323 ( .A(n347), .B(n346), .Z(n559) );
  XOR2_X1 U324 ( .A(n311), .B(n300), .Z(n291) );
  XOR2_X1 U325 ( .A(n302), .B(G71GAT), .Z(n292) );
  AND2_X1 U326 ( .A1(n534), .A2(n524), .ZN(n468) );
  XNOR2_X1 U327 ( .A(G50GAT), .B(KEYINPUT80), .ZN(n326) );
  XNOR2_X1 U328 ( .A(KEYINPUT117), .B(KEYINPUT54), .ZN(n418) );
  NOR2_X1 U329 ( .A1(n482), .A2(n481), .ZN(n495) );
  XNOR2_X1 U330 ( .A(n419), .B(n418), .ZN(n439) );
  NOR2_X1 U331 ( .A1(n439), .A2(n522), .ZN(n565) );
  XNOR2_X1 U332 ( .A(n484), .B(KEYINPUT37), .ZN(n521) );
  XOR2_X1 U333 ( .A(n307), .B(n306), .Z(n308) );
  NOR2_X1 U334 ( .A1(n459), .A2(n458), .ZN(n562) );
  XOR2_X1 U335 ( .A(KEYINPUT84), .B(n559), .Z(n543) );
  XNOR2_X1 U336 ( .A(n490), .B(G190GAT), .ZN(n491) );
  XNOR2_X1 U337 ( .A(n487), .B(G43GAT), .ZN(n488) );
  XNOR2_X1 U338 ( .A(n492), .B(n491), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n489), .B(n488), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT19), .B(KEYINPUT91), .Z(n294) );
  XNOR2_X1 U341 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U343 ( .A(G169GAT), .B(n295), .ZN(n415) );
  XOR2_X1 U344 ( .A(KEYINPUT20), .B(KEYINPUT90), .Z(n297) );
  XNOR2_X1 U345 ( .A(G183GAT), .B(G176GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n307) );
  XOR2_X1 U347 ( .A(G15GAT), .B(G127GAT), .Z(n311) );
  XOR2_X1 U348 ( .A(KEYINPUT89), .B(G99GAT), .Z(n299) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n300) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n291), .B(n301), .ZN(n302) );
  XOR2_X1 U353 ( .A(G120GAT), .B(KEYINPUT0), .Z(n304) );
  XNOR2_X1 U354 ( .A(G113GAT), .B(G134GAT), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n428) );
  XNOR2_X1 U356 ( .A(n428), .B(KEYINPUT92), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n292), .B(n305), .ZN(n306) );
  XOR2_X2 U358 ( .A(n415), .B(n308), .Z(n534) );
  INV_X1 U359 ( .A(n534), .ZN(n459) );
  XOR2_X1 U360 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n349) );
  XOR2_X1 U361 ( .A(G64GAT), .B(KEYINPUT15), .Z(n310) );
  XNOR2_X1 U362 ( .A(KEYINPUT12), .B(KEYINPUT86), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n315) );
  XOR2_X1 U364 ( .A(G22GAT), .B(G155GAT), .Z(n441) );
  XOR2_X1 U365 ( .A(n441), .B(G78GAT), .Z(n313) );
  XNOR2_X1 U366 ( .A(n311), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U368 ( .A(n315), .B(n314), .Z(n317) );
  NAND2_X1 U369 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U371 ( .A(KEYINPUT14), .B(KEYINPUT88), .Z(n319) );
  XNOR2_X1 U372 ( .A(G1GAT), .B(KEYINPUT87), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n325) );
  XNOR2_X1 U375 ( .A(G8GAT), .B(G183GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n322), .B(KEYINPUT85), .ZN(n412) );
  XNOR2_X1 U377 ( .A(G71GAT), .B(G57GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n323), .B(KEYINPUT13), .ZN(n358) );
  XNOR2_X1 U379 ( .A(n412), .B(n358), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n576) );
  INV_X1 U381 ( .A(n576), .ZN(n540) );
  XNOR2_X1 U382 ( .A(n326), .B(G162GAT), .ZN(n445) );
  INV_X1 U383 ( .A(KEYINPUT66), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n445), .B(n327), .ZN(n329) );
  NAND2_X1 U385 ( .A1(G232GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U387 ( .A(KEYINPUT75), .B(G85GAT), .Z(n331) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(G99GAT), .B(n332), .Z(n371) );
  XNOR2_X1 U391 ( .A(n333), .B(n371), .ZN(n347) );
  XOR2_X1 U392 ( .A(KEYINPUT83), .B(KEYINPUT9), .Z(n335) );
  XNOR2_X1 U393 ( .A(KEYINPUT67), .B(KEYINPUT81), .ZN(n334) );
  XNOR2_X1 U394 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U395 ( .A(KEYINPUT11), .B(KEYINPUT82), .Z(n337) );
  XNOR2_X1 U396 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U398 ( .A(n339), .B(n338), .Z(n345) );
  XOR2_X1 U399 ( .A(G29GAT), .B(G43GAT), .Z(n341) );
  XNOR2_X1 U400 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n380) );
  XOR2_X1 U402 ( .A(G92GAT), .B(G218GAT), .Z(n343) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(G190GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n406) );
  XNOR2_X1 U405 ( .A(n380), .B(n406), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U407 ( .A(KEYINPUT36), .B(n543), .ZN(n579) );
  NAND2_X1 U408 ( .A1(n540), .A2(n579), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n350), .B(KEYINPUT68), .ZN(n374) );
  XNOR2_X1 U411 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n352) );
  XNOR2_X1 U412 ( .A(KEYINPUT33), .B(KEYINPUT79), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U414 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n354) );
  XNOR2_X1 U415 ( .A(KEYINPUT77), .B(KEYINPUT72), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n360) );
  XNOR2_X1 U418 ( .A(G78GAT), .B(KEYINPUT74), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n357), .B(G148GAT), .ZN(n452) );
  XNOR2_X1 U420 ( .A(n452), .B(n358), .ZN(n359) );
  XNOR2_X1 U421 ( .A(n360), .B(n359), .ZN(n370) );
  INV_X1 U422 ( .A(G64GAT), .ZN(n361) );
  NAND2_X1 U423 ( .A1(KEYINPUT78), .A2(n361), .ZN(n364) );
  INV_X1 U424 ( .A(KEYINPUT78), .ZN(n362) );
  NAND2_X1 U425 ( .A1(n362), .A2(G64GAT), .ZN(n363) );
  NAND2_X1 U426 ( .A1(n364), .A2(n363), .ZN(n366) );
  XNOR2_X1 U427 ( .A(G176GAT), .B(G204GAT), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n409) );
  XOR2_X1 U429 ( .A(n409), .B(G92GAT), .Z(n368) );
  NAND2_X1 U430 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U432 ( .A(n370), .B(n369), .Z(n373) );
  XNOR2_X1 U433 ( .A(G120GAT), .B(n371), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n572) );
  NAND2_X1 U435 ( .A1(n374), .A2(n572), .ZN(n375) );
  XNOR2_X1 U436 ( .A(KEYINPUT113), .B(n375), .ZN(n392) );
  XOR2_X1 U437 ( .A(G141GAT), .B(G22GAT), .Z(n377) );
  XNOR2_X1 U438 ( .A(G169GAT), .B(G197GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n391) );
  XOR2_X1 U440 ( .A(G50GAT), .B(G36GAT), .Z(n379) );
  NAND2_X1 U441 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U443 ( .A(n381), .B(n380), .Z(n389) );
  XOR2_X1 U444 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n383) );
  XNOR2_X1 U445 ( .A(G15GAT), .B(G113GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U447 ( .A(G1GAT), .B(G8GAT), .Z(n385) );
  XNOR2_X1 U448 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n561) );
  INV_X1 U453 ( .A(n561), .ZN(n566) );
  NAND2_X1 U454 ( .A1(n392), .A2(n566), .ZN(n403) );
  XOR2_X1 U455 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n400) );
  XNOR2_X1 U456 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n572), .B(KEYINPUT65), .ZN(n393) );
  XNOR2_X1 U458 ( .A(KEYINPUT41), .B(n393), .ZN(n553) );
  INV_X1 U459 ( .A(n553), .ZN(n394) );
  NAND2_X1 U460 ( .A1(n394), .A2(n561), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n397) );
  NOR2_X1 U462 ( .A1(n540), .A2(n397), .ZN(n398) );
  NAND2_X1 U463 ( .A1(n398), .A2(n559), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U465 ( .A(KEYINPUT47), .B(n401), .Z(n402) );
  NAND2_X1 U466 ( .A1(n403), .A2(n402), .ZN(n405) );
  XOR2_X1 U467 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n404) );
  XNOR2_X1 U468 ( .A(n405), .B(n404), .ZN(n548) );
  XOR2_X1 U469 ( .A(KEYINPUT96), .B(n406), .Z(n408) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U472 ( .A(n410), .B(n409), .Z(n414) );
  XNOR2_X1 U473 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n411), .B(G211GAT), .ZN(n453) );
  XNOR2_X1 U475 ( .A(n453), .B(n412), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U477 ( .A(n416), .B(n415), .Z(n524) );
  XOR2_X1 U478 ( .A(n524), .B(KEYINPUT116), .Z(n417) );
  NOR2_X1 U479 ( .A1(n548), .A2(n417), .ZN(n419) );
  XOR2_X1 U480 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n421) );
  XNOR2_X1 U481 ( .A(G1GAT), .B(G57GAT), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n438) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G155GAT), .Z(n423) );
  XNOR2_X1 U484 ( .A(G127GAT), .B(G148GAT), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U486 ( .A(G29GAT), .B(G162GAT), .Z(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n434) );
  XOR2_X1 U488 ( .A(KEYINPUT2), .B(KEYINPUT93), .Z(n427) );
  XNOR2_X1 U489 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n428), .B(n440), .ZN(n432) );
  XOR2_X1 U492 ( .A(KEYINPUT94), .B(KEYINPUT6), .Z(n430) );
  XNOR2_X1 U493 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n436) );
  NAND2_X1 U497 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U499 ( .A(n438), .B(n437), .Z(n474) );
  INV_X1 U500 ( .A(n474), .ZN(n522) );
  XOR2_X1 U501 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U502 ( .A1(G228GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U504 ( .A(n444), .B(KEYINPUT23), .Z(n447) );
  XNOR2_X1 U505 ( .A(n445), .B(KEYINPUT22), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U507 ( .A(G204GAT), .B(KEYINPUT24), .Z(n449) );
  XNOR2_X1 U508 ( .A(G218GAT), .B(G106GAT), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U510 ( .A(n451), .B(n450), .Z(n455) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(n477) );
  NAND2_X1 U513 ( .A1(n565), .A2(n477), .ZN(n457) );
  XOR2_X1 U514 ( .A(KEYINPUT118), .B(KEYINPUT55), .Z(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U516 ( .A1(n562), .A2(n540), .ZN(n461) );
  XNOR2_X1 U517 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n461), .B(n460), .ZN(G1350GAT) );
  NAND2_X1 U519 ( .A1(n562), .A2(n394), .ZN(n467) );
  XOR2_X1 U520 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U523 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n467), .B(n466), .ZN(G1349GAT) );
  XNOR2_X1 U526 ( .A(KEYINPUT99), .B(n468), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n477), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(n470), .Z(n473) );
  XNOR2_X1 U529 ( .A(n524), .B(KEYINPUT27), .ZN(n478) );
  NOR2_X1 U530 ( .A1(n534), .A2(n477), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT26), .ZN(n564) );
  NAND2_X1 U532 ( .A1(n478), .A2(n564), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT100), .B(n476), .Z(n482) );
  XOR2_X1 U536 ( .A(n477), .B(KEYINPUT28), .Z(n530) );
  NAND2_X1 U537 ( .A1(n478), .A2(n522), .ZN(n547) );
  NOR2_X1 U538 ( .A1(n530), .A2(n547), .ZN(n535) );
  XNOR2_X1 U539 ( .A(KEYINPUT97), .B(n535), .ZN(n479) );
  NOR2_X1 U540 ( .A1(n534), .A2(n479), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(KEYINPUT98), .ZN(n481) );
  NAND2_X1 U542 ( .A1(n579), .A2(n576), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n495), .A2(n483), .ZN(n484) );
  NAND2_X1 U544 ( .A1(n572), .A2(n561), .ZN(n497) );
  NOR2_X1 U545 ( .A1(n521), .A2(n497), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n508) );
  NAND2_X1 U548 ( .A1(n508), .A2(n534), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n487) );
  NAND2_X1 U550 ( .A1(n562), .A2(n543), .ZN(n492) );
  XOR2_X1 U551 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n490) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n499) );
  NOR2_X1 U553 ( .A1(n543), .A2(n576), .ZN(n493) );
  XOR2_X1 U554 ( .A(KEYINPUT16), .B(n493), .Z(n494) );
  NOR2_X1 U555 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT101), .B(n496), .ZN(n510) );
  NOR2_X1 U557 ( .A1(n497), .A2(n510), .ZN(n503) );
  NAND2_X1 U558 ( .A1(n503), .A2(n522), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1324GAT) );
  NAND2_X1 U560 ( .A1(n524), .A2(n503), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U562 ( .A(G15GAT), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U563 ( .A1(n503), .A2(n534), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n530), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .Z(n506) );
  NAND2_X1 U568 ( .A1(n508), .A2(n522), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NAND2_X1 U570 ( .A1(n524), .A2(n508), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n507), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n508), .A2(n530), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n512) );
  NAND2_X1 U575 ( .A1(n566), .A2(n394), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n510), .A2(n520), .ZN(n516) );
  NAND2_X1 U577 ( .A1(n516), .A2(n522), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n524), .A2(n516), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n513), .B(KEYINPUT104), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n534), .A2(n516), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U585 ( .A1(n516), .A2(n530), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U587 ( .A(G78GAT), .B(n519), .Z(G1335GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n531), .A2(n522), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n531), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(KEYINPUT106), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n528) );
  NAND2_X1 U595 ( .A1(n531), .A2(n534), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n548), .A2(n536), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n561), .A2(n544), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U606 ( .A1(n544), .A2(n394), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n544), .A2(n540), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n549), .A2(n564), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n566), .A2(n558), .ZN(n550) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n550), .Z(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n553), .A2(n558), .ZN(n554) );
  XOR2_X1 U622 ( .A(n555), .B(n554), .Z(G1345GAT) );
  NOR2_X1 U623 ( .A1(n576), .A2(n558), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT115), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n578) );
  NOR2_X1 U631 ( .A1(n566), .A2(n578), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT59), .B(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n578), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n578), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n582) );
  INV_X1 U644 ( .A(n578), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

