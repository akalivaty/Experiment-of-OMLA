

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765;

  XOR2_X1 U366 ( .A(G122), .B(G104), .Z(n502) );
  XNOR2_X1 U367 ( .A(n516), .B(n461), .ZN(n538) );
  INV_X1 U368 ( .A(G953), .ZN(n757) );
  NAND2_X2 U369 ( .A1(n521), .A2(n520), .ZN(n418) );
  XNOR2_X2 U370 ( .A(n434), .B(n433), .ZN(n362) );
  NAND2_X2 U371 ( .A1(n435), .A2(n620), .ZN(n434) );
  XNOR2_X1 U372 ( .A(G143), .B(G113), .ZN(n501) );
  NOR2_X1 U373 ( .A1(n582), .A2(n697), .ZN(n694) );
  NOR2_X2 U374 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X2 U375 ( .A(n686), .B(KEYINPUT6), .ZN(n621) );
  NOR2_X1 U376 ( .A1(n764), .A2(n765), .ZN(n587) );
  XNOR2_X1 U377 ( .A(n581), .B(KEYINPUT42), .ZN(n765) );
  NOR2_X1 U378 ( .A1(n711), .A2(n580), .ZN(n581) );
  INV_X2 U379 ( .A(n623), .ZN(n444) );
  INV_X1 U380 ( .A(KEYINPUT16), .ZN(n387) );
  XNOR2_X1 U381 ( .A(n373), .B(n449), .ZN(n764) );
  XNOR2_X1 U382 ( .A(n619), .B(n618), .ZN(n710) );
  INV_X1 U383 ( .A(n607), .ZN(n344) );
  XNOR2_X1 U384 ( .A(n382), .B(G469), .ZN(n605) );
  XNOR2_X1 U385 ( .A(n532), .B(n387), .ZN(n386) );
  XNOR2_X1 U386 ( .A(n536), .B(n470), .ZN(n500) );
  XOR2_X1 U387 ( .A(G146), .B(G125), .Z(n536) );
  XNOR2_X1 U388 ( .A(n570), .B(n569), .ZN(n580) );
  NOR2_X2 U389 ( .A1(n644), .A2(G902), .ZN(n554) );
  XNOR2_X1 U390 ( .A(n554), .B(n553), .ZN(n607) );
  BUF_X1 U391 ( .A(n723), .Z(n345) );
  BUF_X1 U392 ( .A(n395), .Z(n346) );
  XNOR2_X1 U393 ( .A(n372), .B(n542), .ZN(n723) );
  NOR2_X1 U394 ( .A1(n683), .A2(n551), .ZN(n496) );
  XNOR2_X1 U395 ( .A(n538), .B(n462), .ZN(n751) );
  XNOR2_X1 U396 ( .A(n751), .B(G146), .ZN(n529) );
  AND2_X1 U397 ( .A1(n369), .A2(n368), .ZN(n706) );
  INV_X1 U398 ( .A(KEYINPUT45), .ZN(n441) );
  XNOR2_X1 U399 ( .A(n517), .B(G478), .ZN(n576) );
  XNOR2_X1 U400 ( .A(n487), .B(n486), .ZN(n683) );
  XNOR2_X1 U401 ( .A(n388), .B(G122), .ZN(n532) );
  INV_X1 U402 ( .A(G116), .ZN(n388) );
  XNOR2_X1 U403 ( .A(n605), .B(n381), .ZN(n623) );
  INV_X1 U404 ( .A(KEYINPUT1), .ZN(n381) );
  AND2_X1 U405 ( .A1(n560), .A2(n605), .ZN(n561) );
  INV_X1 U406 ( .A(n411), .ZN(n410) );
  XNOR2_X1 U407 ( .A(n573), .B(n371), .ZN(n370) );
  INV_X1 U408 ( .A(KEYINPUT77), .ZN(n371) );
  INV_X1 U409 ( .A(G101), .ZN(n519) );
  XNOR2_X1 U410 ( .A(n506), .B(n504), .ZN(n424) );
  XOR2_X1 U411 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n504) );
  XOR2_X1 U412 ( .A(G101), .B(G140), .Z(n464) );
  INV_X1 U413 ( .A(KEYINPUT81), .ZN(n547) );
  NOR2_X1 U414 ( .A1(n344), .A2(n564), .ZN(n567) );
  XNOR2_X1 U415 ( .A(n565), .B(KEYINPUT28), .ZN(n566) );
  XNOR2_X1 U416 ( .A(n529), .B(n458), .ZN(n644) );
  XNOR2_X1 U417 ( .A(n528), .B(n530), .ZN(n458) );
  XNOR2_X1 U418 ( .A(n500), .B(n430), .ZN(n429) );
  XNOR2_X1 U419 ( .A(n476), .B(KEYINPUT23), .ZN(n430) );
  NOR2_X1 U420 ( .A1(n753), .A2(KEYINPUT65), .ZN(n406) );
  XNOR2_X1 U421 ( .A(n538), .B(n374), .ZN(n542) );
  XNOR2_X1 U422 ( .A(n537), .B(n541), .ZN(n374) );
  INV_X1 U423 ( .A(KEYINPUT36), .ZN(n378) );
  AND2_X1 U424 ( .A1(n625), .A2(n615), .ZN(n416) );
  INV_X1 U425 ( .A(KEYINPUT97), .ZN(n384) );
  AND2_X1 U426 ( .A1(n687), .A2(n394), .ZN(n393) );
  OR2_X1 U427 ( .A1(n726), .A2(G902), .ZN(n382) );
  XNOR2_X1 U428 ( .A(n511), .B(n375), .ZN(n514) );
  XNOR2_X1 U429 ( .A(KEYINPUT85), .B(n640), .ZN(n725) );
  NOR2_X1 U430 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U431 ( .A1(n437), .A2(KEYINPUT44), .ZN(n398) );
  NAND2_X1 U432 ( .A1(n665), .A2(n695), .ZN(n588) );
  XOR2_X1 U433 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n482) );
  NOR2_X1 U434 ( .A1(G237), .A2(G953), .ZN(n497) );
  NAND2_X1 U435 ( .A1(n638), .A2(KEYINPUT65), .ZN(n411) );
  XNOR2_X1 U436 ( .A(n365), .B(KEYINPUT117), .ZN(n691) );
  OR2_X1 U437 ( .A1(n689), .A2(n690), .ZN(n365) );
  AND2_X1 U438 ( .A1(G953), .A2(G902), .ZN(n489) );
  XOR2_X1 U439 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n484) );
  XNOR2_X1 U440 ( .A(G137), .B(KEYINPUT5), .ZN(n524) );
  XOR2_X1 U441 ( .A(G116), .B(KEYINPUT96), .Z(n525) );
  NAND2_X1 U442 ( .A1(n408), .A2(n447), .ZN(n407) );
  INV_X1 U443 ( .A(KEYINPUT18), .ZN(n539) );
  INV_X1 U444 ( .A(KEYINPUT4), .ZN(n461) );
  INV_X1 U445 ( .A(KEYINPUT48), .ZN(n452) );
  OR2_X1 U446 ( .A1(G237), .A2(G902), .ZN(n546) );
  AND2_X1 U447 ( .A1(n687), .A2(n428), .ZN(n427) );
  NOR2_X1 U448 ( .A1(n582), .A2(n551), .ZN(n428) );
  XNOR2_X1 U449 ( .A(n614), .B(KEYINPUT22), .ZN(n624) );
  XNOR2_X1 U450 ( .A(n532), .B(n348), .ZN(n375) );
  XNOR2_X1 U451 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n509) );
  XOR2_X1 U452 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n510) );
  XNOR2_X1 U453 ( .A(n423), .B(n422), .ZN(n639) );
  XNOR2_X1 U454 ( .A(n503), .B(n500), .ZN(n422) );
  XNOR2_X1 U455 ( .A(n505), .B(n424), .ZN(n423) );
  XNOR2_X1 U456 ( .A(n529), .B(n469), .ZN(n726) );
  XNOR2_X1 U457 ( .A(n468), .B(n467), .ZN(n469) );
  AND2_X1 U458 ( .A1(n687), .A2(n621), .ZN(n442) );
  XNOR2_X1 U459 ( .A(n707), .B(n366), .ZN(n708) );
  XNOR2_X1 U460 ( .A(n367), .B(KEYINPUT119), .ZN(n366) );
  INV_X1 U461 ( .A(KEYINPUT52), .ZN(n367) );
  NAND2_X1 U462 ( .A1(n744), .A2(n631), .ZN(n632) );
  NAND2_X1 U463 ( .A1(G214), .A2(n546), .ZN(n699) );
  INV_X1 U464 ( .A(KEYINPUT35), .ZN(n433) );
  AND2_X1 U465 ( .A1(n568), .A2(n605), .ZN(n570) );
  NOR2_X1 U466 ( .A1(n624), .A2(n444), .ZN(n627) );
  XOR2_X1 U467 ( .A(G128), .B(G119), .Z(n459) );
  INV_X1 U468 ( .A(KEYINPUT40), .ZN(n449) );
  XNOR2_X1 U469 ( .A(n548), .B(n377), .ZN(n549) );
  XNOR2_X1 U470 ( .A(n378), .B(KEYINPUT110), .ZN(n377) );
  INV_X1 U471 ( .A(KEYINPUT32), .ZN(n359) );
  XNOR2_X1 U472 ( .A(n383), .B(n609), .ZN(n670) );
  NOR2_X1 U473 ( .A1(n577), .A2(n572), .ZN(n664) );
  XNOR2_X1 U474 ( .A(n392), .B(n391), .ZN(n563) );
  INV_X1 U475 ( .A(KEYINPUT106), .ZN(n391) );
  NAND2_X1 U476 ( .A1(n561), .A2(n393), .ZN(n392) );
  AND2_X2 U477 ( .A1(n627), .A2(n421), .ZN(n657) );
  AND2_X1 U478 ( .A1(n686), .A2(n615), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n732), .B(n413), .ZN(n735) );
  XNOR2_X1 U480 ( .A(n734), .B(n733), .ZN(n413) );
  INV_X1 U481 ( .A(KEYINPUT56), .ZN(n414) );
  NOR2_X1 U482 ( .A1(n718), .A2(G953), .ZN(n719) );
  INV_X1 U483 ( .A(KEYINPUT44), .ZN(n628) );
  NOR2_X1 U484 ( .A1(n657), .A2(n628), .ZN(n347) );
  XOR2_X1 U485 ( .A(G134), .B(G107), .Z(n348) );
  OR2_X1 U486 ( .A1(KEYINPUT47), .A2(n588), .ZN(n349) );
  AND2_X1 U487 ( .A1(n617), .A2(n650), .ZN(n350) );
  XNOR2_X1 U488 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n351) );
  XOR2_X1 U489 ( .A(KEYINPUT34), .B(KEYINPUT74), .Z(n352) );
  XOR2_X1 U490 ( .A(n639), .B(n351), .Z(n353) );
  XNOR2_X1 U491 ( .A(G902), .B(KEYINPUT15), .ZN(n636) );
  INV_X1 U492 ( .A(KEYINPUT65), .ZN(n447) );
  NAND2_X1 U493 ( .A1(n737), .A2(G475), .ZN(n420) );
  NOR2_X1 U494 ( .A1(n633), .A2(n632), .ZN(n354) );
  NOR2_X1 U495 ( .A1(n633), .A2(n632), .ZN(n680) );
  AND2_X1 U496 ( .A1(n446), .A2(n445), .ZN(n355) );
  AND2_X2 U497 ( .A1(n446), .A2(n445), .ZN(n737) );
  XNOR2_X1 U498 ( .A(n397), .B(n545), .ZN(n550) );
  BUF_X1 U499 ( .A(n390), .Z(n356) );
  NAND2_X1 U500 ( .A1(n629), .A2(n664), .ZN(n373) );
  AND2_X1 U501 ( .A1(n763), .A2(n437), .ZN(n357) );
  NAND2_X1 U502 ( .A1(n626), .A2(KEYINPUT32), .ZN(n360) );
  NAND2_X1 U503 ( .A1(n358), .A2(n359), .ZN(n361) );
  NAND2_X1 U504 ( .A1(n360), .A2(n361), .ZN(n763) );
  INV_X1 U505 ( .A(n626), .ZN(n358) );
  NAND2_X1 U506 ( .A1(n417), .A2(n416), .ZN(n626) );
  BUF_X1 U507 ( .A(n599), .Z(n363) );
  XNOR2_X1 U508 ( .A(n434), .B(n433), .ZN(n762) );
  NAND2_X1 U509 ( .A1(n737), .A2(G210), .ZN(n440) );
  XNOR2_X1 U510 ( .A(n436), .B(n352), .ZN(n435) );
  NAND2_X1 U511 ( .A1(n412), .A2(n406), .ZN(n405) );
  AND2_X1 U512 ( .A1(n762), .A2(n763), .ZN(n400) );
  OR2_X2 U513 ( .A1(n364), .A2(n432), .ZN(n431) );
  NAND2_X1 U514 ( .A1(n364), .A2(n432), .ZN(n535) );
  NAND2_X1 U515 ( .A1(n364), .A2(n747), .ZN(n748) );
  XNOR2_X2 U516 ( .A(n389), .B(n386), .ZN(n364) );
  INV_X1 U517 ( .A(n711), .ZN(n368) );
  XNOR2_X1 U518 ( .A(n693), .B(KEYINPUT51), .ZN(n369) );
  XNOR2_X1 U519 ( .A(n440), .B(n724), .ZN(n419) );
  NOR2_X1 U520 ( .A1(n456), .A2(n370), .ZN(n455) );
  NAND2_X1 U521 ( .A1(n431), .A2(n535), .ZN(n372) );
  NAND2_X1 U522 ( .A1(n550), .A2(n699), .ZN(n396) );
  XNOR2_X1 U523 ( .A(n390), .B(KEYINPUT19), .ZN(n599) );
  XNOR2_X1 U524 ( .A(n420), .B(n353), .ZN(n641) );
  INV_X1 U525 ( .A(n585), .ZN(n584) );
  NAND2_X1 U526 ( .A1(n427), .A2(n561), .ZN(n585) );
  XNOR2_X1 U527 ( .A(n592), .B(n575), .ZN(n696) );
  NAND2_X1 U528 ( .A1(n419), .A2(n725), .ZN(n415) );
  NOR2_X1 U529 ( .A1(n412), .A2(n411), .ZN(n404) );
  NAND2_X1 U530 ( .A1(n376), .A2(n663), .ZN(n573) );
  NAND2_X1 U531 ( .A1(n588), .A2(KEYINPUT47), .ZN(n376) );
  NAND2_X1 U532 ( .A1(n401), .A2(n379), .ZN(n439) );
  NAND2_X1 U533 ( .A1(n400), .A2(n347), .ZN(n379) );
  XNOR2_X1 U534 ( .A(n474), .B(n429), .ZN(n480) );
  XNOR2_X1 U535 ( .A(n380), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U536 ( .A1(n649), .A2(n725), .ZN(n380) );
  NAND2_X1 U537 ( .A1(n670), .A2(n653), .ZN(n610) );
  NAND2_X1 U538 ( .A1(n692), .A2(n385), .ZN(n383) );
  XNOR2_X1 U539 ( .A(n608), .B(n384), .ZN(n692) );
  NAND2_X1 U540 ( .A1(n385), .A2(n613), .ZN(n614) );
  XNOR2_X1 U541 ( .A(n385), .B(KEYINPUT90), .ZN(n395) );
  XNOR2_X2 U542 ( .A(n602), .B(n601), .ZN(n385) );
  XNOR2_X2 U543 ( .A(n534), .B(n533), .ZN(n389) );
  XNOR2_X2 U544 ( .A(n466), .B(G107), .ZN(n533) );
  XNOR2_X2 U545 ( .A(n418), .B(n522), .ZN(n534) );
  NOR2_X1 U546 ( .A1(n589), .A2(n356), .ZN(n548) );
  XNOR2_X2 U547 ( .A(n396), .B(n547), .ZN(n390) );
  NOR2_X1 U548 ( .A1(n592), .A2(n551), .ZN(n394) );
  NAND2_X1 U549 ( .A1(n395), .A2(n710), .ZN(n436) );
  NAND2_X1 U550 ( .A1(n346), .A2(n686), .ZN(n603) );
  NOR2_X2 U551 ( .A1(n723), .A2(n635), .ZN(n397) );
  NAND2_X1 U552 ( .A1(n399), .A2(n398), .ZN(n401) );
  NAND2_X1 U553 ( .A1(n357), .A2(n362), .ZN(n399) );
  NAND2_X1 U554 ( .A1(n402), .A2(n405), .ZN(n446) );
  NOR2_X1 U555 ( .A1(n404), .A2(n403), .ZN(n402) );
  NAND2_X1 U556 ( .A1(n409), .A2(n407), .ZN(n403) );
  NAND2_X1 U557 ( .A1(n753), .A2(n410), .ZN(n409) );
  INV_X1 U558 ( .A(n638), .ZN(n408) );
  NOR2_X2 U559 ( .A1(n634), .A2(n636), .ZN(n412) );
  XNOR2_X1 U560 ( .A(n415), .B(n414), .ZN(G51) );
  INV_X1 U561 ( .A(n624), .ZN(n417) );
  NAND2_X1 U562 ( .A1(n599), .A2(n600), .ZN(n602) );
  NAND2_X1 U563 ( .A1(n451), .A2(n450), .ZN(n629) );
  XNOR2_X2 U564 ( .A(n453), .B(n452), .ZN(n426) );
  NAND2_X1 U565 ( .A1(n426), .A2(n677), .ZN(n633) );
  NAND2_X1 U566 ( .A1(n426), .A2(n425), .ZN(n448) );
  AND2_X1 U567 ( .A1(n677), .A2(n676), .ZN(n425) );
  INV_X1 U568 ( .A(n687), .ZN(n606) );
  INV_X1 U569 ( .A(KEYINPUT83), .ZN(n432) );
  NAND2_X1 U570 ( .A1(n657), .A2(n628), .ZN(n437) );
  XNOR2_X2 U571 ( .A(n438), .B(n441), .ZN(n634) );
  NAND2_X1 U572 ( .A1(n439), .A2(n350), .ZN(n438) );
  XNOR2_X2 U573 ( .A(G119), .B(KEYINPUT3), .ZN(n522) );
  XNOR2_X1 U574 ( .A(n587), .B(KEYINPUT46), .ZN(n454) );
  XNOR2_X2 U575 ( .A(n554), .B(n552), .ZN(n686) );
  NAND2_X1 U576 ( .A1(n457), .A2(n349), .ZN(n456) );
  XNOR2_X1 U577 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U578 ( .A1(n444), .A2(n442), .ZN(n618) );
  NAND2_X1 U579 ( .A1(n444), .A2(n687), .ZN(n443) );
  NOR2_X1 U580 ( .A1(n443), .A2(n344), .ZN(n608) );
  INV_X1 U581 ( .A(n354), .ZN(n445) );
  NOR2_X1 U582 ( .A1(n753), .A2(n634), .ZN(n678) );
  XNOR2_X2 U583 ( .A(n448), .B(KEYINPUT80), .ZN(n753) );
  NAND2_X1 U584 ( .A1(n584), .A2(n583), .ZN(n450) );
  NAND2_X1 U585 ( .A1(n585), .A2(n586), .ZN(n451) );
  NAND2_X1 U586 ( .A1(n455), .A2(n454), .ZN(n453) );
  INV_X1 U587 ( .A(n675), .ZN(n457) );
  XNOR2_X1 U588 ( .A(G140), .B(KEYINPUT10), .ZN(n470) );
  INV_X1 U589 ( .A(KEYINPUT38), .ZN(n574) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n574), .B(KEYINPUT71), .ZN(n575) );
  INV_X1 U592 ( .A(KEYINPUT107), .ZN(n565) );
  XNOR2_X1 U593 ( .A(n498), .B(G134), .ZN(n462) );
  XNOR2_X1 U594 ( .A(n540), .B(n539), .ZN(n541) );
  INV_X1 U595 ( .A(KEYINPUT0), .ZN(n601) );
  XNOR2_X1 U596 ( .A(n579), .B(n578), .ZN(n711) );
  XNOR2_X2 U597 ( .A(G128), .B(KEYINPUT64), .ZN(n460) );
  XNOR2_X2 U598 ( .A(n460), .B(G143), .ZN(n516) );
  XNOR2_X1 U599 ( .A(KEYINPUT66), .B(G131), .ZN(n498) );
  NAND2_X1 U600 ( .A1(G227), .A2(n757), .ZN(n463) );
  XNOR2_X1 U601 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U602 ( .A(G137), .B(KEYINPUT67), .ZN(n475) );
  XNOR2_X1 U603 ( .A(KEYINPUT91), .B(n475), .ZN(n750) );
  XOR2_X1 U604 ( .A(n465), .B(n750), .Z(n468) );
  XNOR2_X2 U605 ( .A(G110), .B(G104), .ZN(n466) );
  BUF_X1 U606 ( .A(n533), .Z(n467) );
  XOR2_X1 U607 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n472) );
  XNOR2_X1 U608 ( .A(KEYINPUT68), .B(KEYINPUT24), .ZN(n471) );
  XNOR2_X1 U609 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U610 ( .A(G110), .B(n473), .ZN(n474) );
  INV_X1 U611 ( .A(n475), .ZN(n476) );
  NAND2_X1 U612 ( .A1(G234), .A2(n757), .ZN(n477) );
  XOR2_X1 U613 ( .A(KEYINPUT8), .B(n477), .Z(n512) );
  NAND2_X1 U614 ( .A1(n512), .A2(G221), .ZN(n478) );
  XNOR2_X1 U615 ( .A(n478), .B(n459), .ZN(n479) );
  XNOR2_X1 U616 ( .A(n480), .B(n479), .ZN(n736) );
  NOR2_X1 U617 ( .A1(G902), .A2(n736), .ZN(n487) );
  NAND2_X1 U618 ( .A1(G234), .A2(n636), .ZN(n481) );
  XNOR2_X1 U619 ( .A(n482), .B(n481), .ZN(n494) );
  NAND2_X1 U620 ( .A1(G217), .A2(n494), .ZN(n483) );
  XNOR2_X1 U621 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U622 ( .A(KEYINPUT94), .B(n485), .ZN(n486) );
  NAND2_X1 U623 ( .A1(G234), .A2(G237), .ZN(n488) );
  XNOR2_X1 U624 ( .A(KEYINPUT14), .B(n488), .ZN(n491) );
  NAND2_X1 U625 ( .A1(n491), .A2(n489), .ZN(n594) );
  XOR2_X1 U626 ( .A(n594), .B(KEYINPUT105), .Z(n490) );
  NOR2_X1 U627 ( .A1(G900), .A2(n490), .ZN(n493) );
  NAND2_X1 U628 ( .A1(G952), .A2(n491), .ZN(n709) );
  NOR2_X1 U629 ( .A1(n709), .A2(G953), .ZN(n492) );
  XNOR2_X1 U630 ( .A(n492), .B(KEYINPUT88), .ZN(n596) );
  NOR2_X1 U631 ( .A1(n493), .A2(n596), .ZN(n551) );
  NAND2_X1 U632 ( .A1(n494), .A2(G221), .ZN(n495) );
  XOR2_X1 U633 ( .A(KEYINPUT21), .B(n495), .Z(n682) );
  NAND2_X1 U634 ( .A1(n496), .A2(n682), .ZN(n564) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(G475), .ZN(n508) );
  XNOR2_X1 U636 ( .A(n497), .B(KEYINPUT72), .ZN(n523) );
  NAND2_X1 U637 ( .A1(n523), .A2(G214), .ZN(n506) );
  INV_X1 U638 ( .A(n498), .ZN(n499) );
  XNOR2_X1 U639 ( .A(n499), .B(KEYINPUT12), .ZN(n505) );
  XNOR2_X1 U640 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U641 ( .A1(G902), .A2(n639), .ZN(n507) );
  XOR2_X1 U642 ( .A(n508), .B(n507), .Z(n577) );
  XNOR2_X1 U643 ( .A(n510), .B(n509), .ZN(n511) );
  NAND2_X1 U644 ( .A1(G217), .A2(n512), .ZN(n513) );
  XNOR2_X1 U645 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U646 ( .A(n516), .B(n515), .ZN(n734) );
  NOR2_X1 U647 ( .A1(n734), .A2(G902), .ZN(n517) );
  INV_X1 U648 ( .A(n576), .ZN(n572) );
  INV_X1 U649 ( .A(n664), .ZN(n667) );
  NOR2_X1 U650 ( .A1(n564), .A2(n667), .ZN(n531) );
  INV_X1 U651 ( .A(G113), .ZN(n518) );
  NAND2_X1 U652 ( .A1(n518), .A2(G101), .ZN(n521) );
  NAND2_X1 U653 ( .A1(n519), .A2(G113), .ZN(n520) );
  BUF_X1 U654 ( .A(n534), .Z(n530) );
  AND2_X1 U655 ( .A1(G210), .A2(n523), .ZN(n527) );
  XNOR2_X1 U656 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U657 ( .A(G472), .B(KEYINPUT70), .ZN(n552) );
  NAND2_X1 U658 ( .A1(n531), .A2(n621), .ZN(n589) );
  XNOR2_X1 U659 ( .A(n536), .B(KEYINPUT17), .ZN(n537) );
  NAND2_X1 U660 ( .A1(G224), .A2(n757), .ZN(n540) );
  INV_X1 U661 ( .A(n636), .ZN(n635) );
  XOR2_X1 U662 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n544) );
  NAND2_X1 U663 ( .A1(G210), .A2(n546), .ZN(n543) );
  XNOR2_X1 U664 ( .A(n544), .B(n543), .ZN(n545) );
  NOR2_X1 U665 ( .A1(n623), .A2(n549), .ZN(n675) );
  INV_X1 U666 ( .A(n550), .ZN(n592) );
  INV_X1 U667 ( .A(n682), .ZN(n611) );
  INV_X1 U668 ( .A(n683), .ZN(n615) );
  NOR2_X2 U669 ( .A1(n611), .A2(n615), .ZN(n687) );
  INV_X1 U670 ( .A(KEYINPUT30), .ZN(n555) );
  INV_X1 U671 ( .A(n552), .ZN(n553) );
  NAND2_X1 U672 ( .A1(n607), .A2(n699), .ZN(n556) );
  NAND2_X1 U673 ( .A1(n555), .A2(n556), .ZN(n559) );
  INV_X1 U674 ( .A(n556), .ZN(n557) );
  NAND2_X1 U675 ( .A1(KEYINPUT30), .A2(n557), .ZN(n558) );
  NAND2_X1 U676 ( .A1(n559), .A2(n558), .ZN(n560) );
  OR2_X1 U677 ( .A1(n576), .A2(n577), .ZN(n562) );
  XOR2_X1 U678 ( .A(KEYINPUT104), .B(n562), .Z(n620) );
  NAND2_X1 U679 ( .A1(n563), .A2(n620), .ZN(n663) );
  INV_X1 U680 ( .A(KEYINPUT108), .ZN(n569) );
  INV_X1 U681 ( .A(n363), .ZN(n571) );
  NOR2_X2 U682 ( .A1(n580), .A2(n571), .ZN(n665) );
  NAND2_X1 U683 ( .A1(n572), .A2(n577), .ZN(n669) );
  NAND2_X1 U684 ( .A1(n667), .A2(n669), .ZN(n695) );
  INV_X1 U685 ( .A(n696), .ZN(n582) );
  NAND2_X1 U686 ( .A1(n577), .A2(n576), .ZN(n697) );
  NAND2_X1 U687 ( .A1(n699), .A2(n694), .ZN(n579) );
  XNOR2_X1 U688 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n578) );
  XNOR2_X1 U689 ( .A(KEYINPUT69), .B(KEYINPUT39), .ZN(n583) );
  INV_X1 U690 ( .A(n583), .ZN(n586) );
  NOR2_X1 U691 ( .A1(n444), .A2(n589), .ZN(n590) );
  NAND2_X1 U692 ( .A1(n590), .A2(n699), .ZN(n591) );
  XNOR2_X1 U693 ( .A(KEYINPUT43), .B(n591), .ZN(n593) );
  NAND2_X1 U694 ( .A1(n593), .A2(n592), .ZN(n677) );
  NOR2_X1 U695 ( .A1(G898), .A2(n594), .ZN(n595) );
  XNOR2_X1 U696 ( .A(KEYINPUT89), .B(n595), .ZN(n598) );
  INV_X1 U697 ( .A(n596), .ZN(n597) );
  NAND2_X1 U698 ( .A1(n598), .A2(n597), .ZN(n600) );
  NOR2_X1 U699 ( .A1(n606), .A2(n603), .ZN(n604) );
  NAND2_X1 U700 ( .A1(n605), .A2(n604), .ZN(n653) );
  XOR2_X1 U701 ( .A(KEYINPUT98), .B(KEYINPUT31), .Z(n609) );
  NAND2_X1 U702 ( .A1(n610), .A2(n695), .ZN(n617) );
  NOR2_X1 U703 ( .A1(n611), .A2(n697), .ZN(n612) );
  XNOR2_X1 U704 ( .A(KEYINPUT102), .B(n612), .ZN(n613) );
  NOR2_X1 U705 ( .A1(n621), .A2(n615), .ZN(n616) );
  NAND2_X1 U706 ( .A1(n627), .A2(n616), .ZN(n650) );
  XOR2_X1 U707 ( .A(KEYINPUT103), .B(KEYINPUT33), .Z(n619) );
  XOR2_X1 U708 ( .A(KEYINPUT75), .B(n621), .Z(n622) );
  NOR2_X1 U709 ( .A1(n623), .A2(n622), .ZN(n625) );
  INV_X1 U710 ( .A(n634), .ZN(n744) );
  INV_X1 U711 ( .A(n669), .ZN(n659) );
  NAND2_X1 U712 ( .A1(n659), .A2(n629), .ZN(n676) );
  NAND2_X1 U713 ( .A1(KEYINPUT2), .A2(n676), .ZN(n630) );
  XOR2_X1 U714 ( .A(KEYINPUT76), .B(n630), .Z(n631) );
  XNOR2_X1 U715 ( .A(n636), .B(KEYINPUT79), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n637), .A2(KEYINPUT2), .ZN(n638) );
  NOR2_X1 U717 ( .A1(G952), .A2(n757), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n725), .ZN(n643) );
  INV_X1 U719 ( .A(KEYINPUT60), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n643), .B(n642), .ZN(G60) );
  NAND2_X1 U721 ( .A1(n737), .A2(G472), .ZN(n648) );
  XOR2_X1 U722 ( .A(KEYINPUT84), .B(KEYINPUT62), .Z(n646) );
  XOR2_X1 U723 ( .A(n644), .B(KEYINPUT111), .Z(n645) );
  XNOR2_X1 U724 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U726 ( .A(G101), .B(n650), .ZN(G3) );
  NOR2_X1 U727 ( .A1(n667), .A2(n653), .ZN(n651) );
  XOR2_X1 U728 ( .A(KEYINPUT112), .B(n651), .Z(n652) );
  XNOR2_X1 U729 ( .A(G104), .B(n652), .ZN(G6) );
  NOR2_X1 U730 ( .A1(n669), .A2(n653), .ZN(n655) );
  XNOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U733 ( .A(G107), .B(n656), .ZN(G9) );
  XNOR2_X1 U734 ( .A(G110), .B(n657), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(KEYINPUT113), .ZN(G12) );
  XOR2_X1 U736 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n661) );
  NAND2_X1 U737 ( .A1(n665), .A2(n659), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U739 ( .A(G128), .B(n662), .ZN(G30) );
  XNOR2_X1 U740 ( .A(G143), .B(n663), .ZN(G45) );
  NAND2_X1 U741 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n666), .B(G146), .ZN(G48) );
  NOR2_X1 U743 ( .A1(n670), .A2(n667), .ZN(n668) );
  XOR2_X1 U744 ( .A(G113), .B(n668), .Z(G15) );
  NOR2_X1 U745 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U746 ( .A(G116), .B(n671), .Z(G18) );
  XOR2_X1 U747 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n673) );
  XNOR2_X1 U748 ( .A(G125), .B(KEYINPUT37), .ZN(n672) );
  XNOR2_X1 U749 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U750 ( .A(n675), .B(n674), .ZN(G27) );
  XNOR2_X1 U751 ( .A(G134), .B(n676), .ZN(G36) );
  XNOR2_X1 U752 ( .A(G140), .B(n677), .ZN(G42) );
  NOR2_X1 U753 ( .A1(KEYINPUT2), .A2(n678), .ZN(n679) );
  XOR2_X1 U754 ( .A(KEYINPUT78), .B(n681), .Z(n717) );
  NOR2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n684), .B(KEYINPUT49), .ZN(n685) );
  NAND2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n687), .A2(n444), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT50), .ZN(n689) );
  NOR2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  INV_X1 U761 ( .A(n694), .ZN(n702) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U766 ( .A1(n710), .A2(n703), .ZN(n704) );
  XOR2_X1 U767 ( .A(KEYINPUT118), .B(n704), .Z(n705) );
  NOR2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U769 ( .A1(n709), .A2(n708), .ZN(n714) );
  INV_X1 U770 ( .A(n710), .ZN(n712) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U772 ( .A(KEYINPUT120), .B(n715), .ZN(n716) );
  NAND2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n719), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U775 ( .A(KEYINPUT55), .B(KEYINPUT82), .Z(n721) );
  XNOR2_X1 U776 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n720) );
  XNOR2_X1 U777 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n345), .B(n722), .ZN(n724) );
  INV_X1 U779 ( .A(n725), .ZN(n741) );
  XOR2_X1 U780 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n728) );
  XNOR2_X1 U781 ( .A(n726), .B(KEYINPUT122), .ZN(n727) );
  XNOR2_X1 U782 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n355), .A2(G469), .ZN(n729) );
  XNOR2_X1 U784 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U785 ( .A1(n741), .A2(n731), .ZN(G54) );
  XOR2_X1 U786 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n733) );
  NAND2_X1 U787 ( .A1(n355), .A2(G478), .ZN(n732) );
  NOR2_X1 U788 ( .A1(n741), .A2(n735), .ZN(G63) );
  XNOR2_X1 U789 ( .A(n736), .B(KEYINPUT126), .ZN(n739) );
  NAND2_X1 U790 ( .A1(G217), .A2(n355), .ZN(n738) );
  XNOR2_X1 U791 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U792 ( .A1(n741), .A2(n740), .ZN(G66) );
  NAND2_X1 U793 ( .A1(G953), .A2(G224), .ZN(n742) );
  XNOR2_X1 U794 ( .A(KEYINPUT61), .B(n742), .ZN(n743) );
  NAND2_X1 U795 ( .A1(n743), .A2(G898), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n744), .A2(n757), .ZN(n745) );
  NAND2_X1 U797 ( .A1(n746), .A2(n745), .ZN(n749) );
  OR2_X1 U798 ( .A1(n757), .A2(G898), .ZN(n747) );
  XOR2_X1 U799 ( .A(n749), .B(n748), .Z(G69) );
  XNOR2_X1 U800 ( .A(n750), .B(n500), .ZN(n752) );
  XOR2_X1 U801 ( .A(n751), .B(n752), .Z(n755) );
  XOR2_X1 U802 ( .A(n755), .B(n753), .Z(n754) );
  NAND2_X1 U803 ( .A1(n754), .A2(n757), .ZN(n760) );
  XOR2_X1 U804 ( .A(G227), .B(n755), .Z(n756) );
  NOR2_X1 U805 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U806 ( .A1(G900), .A2(n758), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U808 ( .A(KEYINPUT127), .B(n761), .ZN(G72) );
  XNOR2_X1 U809 ( .A(n362), .B(G122), .ZN(G24) );
  XNOR2_X1 U810 ( .A(n763), .B(G119), .ZN(G21) );
  XOR2_X1 U811 ( .A(n764), .B(G131), .Z(G33) );
  XOR2_X1 U812 ( .A(G137), .B(n765), .Z(G39) );
endmodule

