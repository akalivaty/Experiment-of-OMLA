//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT31), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G50gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT77), .B(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT78), .ZN(new_n213));
  XOR2_X1   g012(.A(G211gat), .B(G218gat), .Z(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n214), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(KEYINPUT78), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT29), .ZN(new_n218));
  XNOR2_X1  g017(.A(G141gat), .B(G148gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n222), .B(new_n221), .C1(new_n219), .C2(KEYINPUT2), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n215), .A2(new_n217), .B1(new_n218), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(G228gat), .B2(G233gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n225), .A2(new_n226), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n212), .A2(new_n216), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT29), .B1(new_n212), .B2(new_n216), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n230), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G22gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n218), .A3(new_n217), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n232), .B1(new_n238), .B2(new_n227), .ZN(new_n239));
  OAI211_X1 g038(.A(G228gat), .B(G233gat), .C1(new_n239), .C2(new_n229), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n237), .B1(new_n236), .B2(new_n240), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n206), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n241), .A3(new_n205), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G169gat), .ZN(new_n249));
  INV_X1    g048(.A(G176gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT23), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(G169gat), .B2(G176gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT24), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n261), .A2(new_n262), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT25), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT25), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n255), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n256), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n257), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n260), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT68), .B(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n269), .A2(KEYINPUT67), .A3(new_n257), .A4(new_n270), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n267), .B1(new_n279), .B2(KEYINPUT69), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n273), .A2(new_n277), .A3(new_n281), .A4(new_n278), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n265), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n254), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n249), .A2(new_n250), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n284), .B1(KEYINPUT26), .B2(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(KEYINPUT26), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n286), .A2(new_n287), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n275), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT28), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n218), .B1(new_n283), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G226gat), .A2(G233gat), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT79), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n215), .A2(new_n217), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n302));
  INV_X1    g101(.A(new_n267), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n282), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n265), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n295), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n297), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(new_n297), .B2(new_n296), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n299), .B(new_n301), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n297), .B1(new_n312), .B2(KEYINPUT29), .ZN(new_n313));
  OAI211_X1 g112(.A(G226gat), .B(G233gat), .C1(new_n283), .C2(new_n295), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n301), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G64gat), .B(G92gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT80), .ZN(new_n318));
  XOR2_X1   g117(.A(G8gat), .B(G36gat), .Z(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n311), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G57gat), .B(G85gat), .Z(new_n322));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G120gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G113gat), .ZN(new_n329));
  INV_X1    g128(.A(G113gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT71), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G134gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT72), .B1(new_n336), .B2(G127gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n335), .A3(G134gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n334), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n332), .A2(new_n346), .A3(new_n333), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n348), .A2(new_n228), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n231), .A2(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n348), .A2(new_n231), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n348), .A2(new_n231), .A3(KEYINPUT4), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n351), .B(new_n352), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n352), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n348), .A2(new_n231), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n353), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT5), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT5), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n361), .B1(new_n357), .B2(new_n363), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n327), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n363), .ZN(new_n368));
  INV_X1    g167(.A(new_n361), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n326), .B(KEYINPUT85), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n372), .A3(new_n364), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n367), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n365), .A2(new_n366), .A3(new_n327), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT6), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n321), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n299), .B(new_n300), .C1(new_n309), .C2(new_n310), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT37), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n313), .A2(new_n314), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n381), .B2(new_n301), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT38), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n320), .B1(new_n311), .B2(new_n316), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n320), .A2(new_n380), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT38), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n298), .B1(new_n381), .B2(KEYINPUT79), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n315), .B1(new_n389), .B2(new_n301), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n320), .B1(new_n390), .B2(new_n380), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n311), .A2(new_n316), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT37), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n248), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n345), .A2(new_n347), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n232), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n398));
  INV_X1    g197(.A(new_n356), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n398), .A2(new_n399), .B1(new_n349), .B2(new_n350), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT86), .B1(new_n400), .B2(new_n352), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT86), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n358), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n348), .A2(new_n231), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n397), .A2(new_n352), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT39), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT88), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(new_n404), .A3(new_n401), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n412), .A3(new_n371), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT40), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n407), .A2(new_n412), .A3(KEYINPUT40), .A4(new_n371), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n373), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n311), .A2(KEYINPUT30), .A3(new_n316), .A4(new_n320), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT81), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n390), .A2(new_n420), .A3(KEYINPUT30), .A4(new_n320), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n384), .B1(new_n423), .B2(new_n321), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n417), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n395), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n367), .A2(new_n374), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n377), .B1(new_n427), .B2(new_n376), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n428), .A3(new_n424), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n247), .ZN(new_n430));
  XOR2_X1   g229(.A(G15gat), .B(G43gat), .Z(new_n431));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G227gat), .ZN(new_n434));
  INV_X1    g233(.A(G233gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n436), .B(KEYINPUT64), .Z(new_n437));
  NAND3_X1  g236(.A1(new_n306), .A2(new_n396), .A3(new_n307), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n348), .B1(new_n283), .B2(new_n295), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(KEYINPUT32), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n433), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT74), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n433), .A2(KEYINPUT73), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT33), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n433), .A2(KEYINPUT73), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT32), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n444), .B1(new_n440), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n437), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n396), .B1(new_n306), .B2(new_n307), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n348), .B(new_n295), .C1(new_n304), .C2(new_n305), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n448), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(KEYINPUT74), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n443), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT75), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT75), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n443), .A2(new_n449), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n438), .A2(new_n439), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n461), .A2(KEYINPUT34), .A3(new_n450), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT34), .B1(new_n461), .B2(new_n436), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n464), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n457), .A2(new_n466), .A3(new_n459), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(KEYINPUT36), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT36), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n457), .A2(new_n466), .A3(new_n459), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n457), .B2(new_n459), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n430), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n426), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n430), .A2(KEYINPUT84), .A3(new_n468), .A4(new_n472), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n248), .B1(new_n470), .B2(new_n471), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n478));
  INV_X1    g277(.A(new_n429), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(new_n248), .C1(new_n470), .C2(new_n471), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n248), .A2(new_n422), .A3(new_n424), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n470), .B2(new_n471), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n465), .A2(KEYINPUT89), .A3(new_n467), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT35), .B1(new_n375), .B2(new_n377), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n475), .A2(new_n476), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(G113gat), .B(G141gat), .Z(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT91), .B(G197gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT11), .B(G169gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(KEYINPUT12), .Z(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g304(.A1(G43gat), .A2(G50gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT92), .B(G50gat), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n505), .B(new_n506), .C1(new_n507), .C2(G43gat), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n508), .B2(KEYINPUT93), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(KEYINPUT93), .B2(new_n508), .ZN(new_n510));
  NOR2_X1   g309(.A1(G43gat), .A2(G50gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n505), .B1(new_n512), .B2(new_n506), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n514), .A2(new_n504), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G15gat), .B(G22gat), .Z(new_n519));
  INV_X1    g318(.A(G1gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(G8gat), .B1(new_n521), .B2(KEYINPUT94), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(KEYINPUT16), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n523), .B2(new_n519), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n524), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT95), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n518), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n530), .A3(new_n516), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n528), .B1(new_n532), .B2(KEYINPUT95), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n499), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT18), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n517), .B(new_n527), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(new_n499), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(KEYINPUT18), .B(new_n499), .C1(new_n531), .C2(new_n533), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n498), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n536), .A2(new_n498), .A3(new_n542), .A4(new_n540), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n536), .A2(new_n540), .ZN(new_n548));
  INV_X1    g347(.A(new_n542), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n497), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(new_n545), .A3(new_n544), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n202), .B1(new_n491), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n429), .A2(new_n247), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n472), .A2(new_n468), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n474), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n426), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n557), .A2(new_n558), .A3(new_n476), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n482), .A2(KEYINPUT35), .B1(new_n488), .B2(new_n489), .ZN(new_n560));
  OAI211_X1 g359(.A(KEYINPUT98), .B(new_n554), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G230gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(new_n435), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT102), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT101), .Z(new_n571));
  OAI21_X1  g370(.A(KEYINPUT7), .B1(new_n566), .B2(new_n567), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT100), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n568), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G99gat), .B(G106gat), .Z(new_n575));
  AOI21_X1  g374(.A(new_n564), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n575), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n574), .B(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n579), .B2(KEYINPUT102), .ZN(new_n580));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G71gat), .B(G78gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT104), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n574), .B(new_n575), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(new_n585), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n580), .A2(KEYINPUT104), .A3(new_n585), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n588), .A2(new_n589), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n580), .A2(new_n589), .A3(new_n585), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n563), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n563), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n592), .A2(new_n591), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n597), .B2(new_n588), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n602), .B1(new_n595), .B2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n576), .B1(new_n590), .B2(new_n564), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n517), .B1(new_n608), .B2(KEYINPUT17), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n580), .A2(new_n530), .A3(new_n518), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n613));
  XOR2_X1   g412(.A(G190gat), .B(G218gat), .Z(new_n614));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n618), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n615), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  OR2_X1    g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT21), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n585), .B1(new_n527), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT99), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G183gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G211gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n631), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n527), .A2(new_n628), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n636), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n607), .A2(new_n627), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n553), .A2(new_n561), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n428), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g445(.A1(new_n422), .A2(new_n424), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n553), .A2(new_n647), .A3(new_n561), .A4(new_n642), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n648), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT105), .B1(new_n648), .B2(G8gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT16), .B(G8gat), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n643), .A2(KEYINPUT42), .A3(new_n647), .A4(new_n654), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n651), .A2(new_n652), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n648), .A2(G8gat), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n648), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n661), .A2(new_n657), .A3(new_n656), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT106), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(G1325gat));
  NAND2_X1  g464(.A1(new_n486), .A2(new_n487), .ZN(new_n666));
  AOI21_X1  g465(.A(G15gat), .B1(new_n643), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n556), .B(KEYINPUT107), .Z(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G15gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n643), .B2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n643), .A2(new_n247), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NOR3_X1   g472(.A1(new_n627), .A2(new_n640), .A3(new_n606), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n428), .A2(G29gat), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n553), .A2(new_n561), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n627), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n473), .A2(new_n426), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n560), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n684), .C1(new_n559), .C2(new_n560), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n543), .A2(new_n546), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n545), .B(new_n498), .C1(new_n541), .C2(new_n542), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n547), .A2(KEYINPUT110), .A3(new_n551), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(new_n640), .A3(new_n606), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n428), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n699), .A3(new_n700), .ZN(G1328gat));
  AND2_X1   g500(.A1(new_n553), .A2(new_n561), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n674), .ZN(new_n703));
  INV_X1    g502(.A(G36gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n647), .A2(new_n704), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n703), .A2(KEYINPUT46), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n647), .ZN(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n698), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT46), .B1(new_n703), .B2(new_n705), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(G1329gat));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711));
  INV_X1    g510(.A(G43gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n698), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(new_n668), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n702), .A2(new_n712), .A3(new_n666), .A4(new_n674), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n711), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n556), .ZN(new_n718));
  OAI21_X1  g517(.A(G43gat), .B1(new_n698), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(KEYINPUT47), .A3(new_n715), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(G1330gat));
  OAI21_X1  g520(.A(new_n507), .B1(new_n698), .B2(new_n248), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n248), .A2(new_n507), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n703), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n722), .B(KEYINPUT48), .C1(new_n703), .C2(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1331gat));
  OR2_X1    g527(.A1(new_n560), .A2(new_n685), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n694), .A2(new_n695), .ZN(new_n730));
  INV_X1    g529(.A(new_n640), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n730), .A2(new_n684), .A3(new_n607), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(new_n644), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT111), .B(G57gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1332gat));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n732), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n707), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  INV_X1    g542(.A(new_n668), .ZN(new_n744));
  OAI21_X1  g543(.A(G71gat), .B1(new_n738), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n666), .A3(new_n732), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT113), .ZN(new_n747));
  INV_X1    g546(.A(G71gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n745), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n745), .B2(new_n749), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n248), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g554(.A1(new_n730), .A2(new_n640), .A3(new_n607), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n690), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n428), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n730), .A2(new_n640), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n759), .B(new_n684), .C1(new_n560), .C2(new_n685), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n606), .A2(new_n566), .A3(new_n644), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n758), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n757), .B2(new_n707), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n729), .A2(KEYINPUT51), .A3(new_n684), .A4(new_n759), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n760), .A2(new_n761), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(KEYINPUT114), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n762), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n607), .A2(G92gat), .A3(new_n707), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT52), .ZN(new_n776));
  INV_X1    g575(.A(new_n764), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(new_n777), .B2(new_n773), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n767), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n757), .B2(new_n744), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n607), .B1(new_n487), .B2(new_n486), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n783), .A2(G99gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n764), .B2(new_n784), .ZN(G1338gat));
  NOR3_X1   g584(.A1(new_n607), .A2(G106gat), .A3(new_n248), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n772), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n688), .A2(new_n689), .A3(new_n247), .A4(new_n756), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n762), .B2(new_n763), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(KEYINPUT115), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n787), .B2(new_n789), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n789), .A2(new_n792), .A3(new_n793), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1339gat));
  NAND4_X1  g599(.A1(new_n696), .A2(new_n640), .A3(new_n627), .A4(new_n607), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n593), .A2(new_n594), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n596), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n593), .A2(new_n563), .A3(new_n594), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n806));
  AOI21_X1  g605(.A(new_n603), .B1(new_n595), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n604), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n531), .A2(new_n533), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n813), .A2(new_n499), .B1(new_n537), .B2(new_n539), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n496), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n544), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n625), .A2(new_n626), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n606), .A2(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n696), .B2(new_n812), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n627), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n801), .B1(new_n821), .B2(new_n640), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n644), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n554), .A3(new_n488), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G113gat), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n478), .A2(new_n481), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n707), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n823), .A2(new_n330), .A3(new_n730), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n825), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1340gat));
  AND2_X1   g632(.A1(new_n823), .A2(new_n488), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n606), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n823), .A2(new_n827), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n606), .A2(new_n328), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n835), .A2(new_n328), .B1(new_n836), .B2(new_n837), .ZN(G1341gat));
  INV_X1    g637(.A(new_n836), .ZN(new_n839));
  AOI21_X1  g638(.A(G127gat), .B1(new_n839), .B2(new_n640), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n731), .A2(new_n335), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n834), .B2(new_n841), .ZN(G1342gat));
  AOI21_X1  g641(.A(new_n627), .B1(new_n337), .B2(new_n339), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n823), .A2(new_n488), .A3(new_n684), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n844), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n844), .B2(KEYINPUT56), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n839), .A2(KEYINPUT118), .A3(new_n849), .A4(new_n843), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(G141gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n811), .A2(new_n604), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n805), .B2(new_n807), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n552), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n819), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n627), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n818), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n640), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n801), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n247), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT57), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n822), .A2(new_n863), .A3(new_n247), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n556), .A2(new_n428), .A3(new_n647), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n852), .B1(new_n866), .B2(new_n730), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n668), .A2(new_n428), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n822), .A2(new_n247), .A3(new_n868), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n869), .A2(G141gat), .A3(new_n552), .A4(new_n647), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT58), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n552), .A2(G141gat), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n822), .A2(new_n874), .A3(new_n247), .A4(new_n868), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n872), .A2(new_n707), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT120), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n864), .A3(new_n554), .A4(new_n865), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT58), .B1(new_n878), .B2(G141gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n647), .B1(new_n869), .B2(KEYINPUT119), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n873), .A4(new_n875), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n877), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n871), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n822), .A2(new_n247), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT57), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n641), .A2(new_n554), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT121), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n863), .B(new_n247), .C1(new_n889), .C2(new_n859), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n887), .A2(new_n890), .A3(new_n606), .A4(new_n865), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n885), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n885), .A2(G148gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n866), .B2(new_n606), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n880), .A2(new_n875), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n607), .A2(G148gat), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n892), .A2(new_n894), .B1(new_n895), .B2(new_n896), .ZN(G1345gat));
  NAND3_X1  g696(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n898));
  OAI21_X1  g697(.A(G155gat), .B1(new_n898), .B2(new_n731), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n731), .A2(G155gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n880), .A2(new_n875), .A3(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n899), .B2(new_n901), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(G1346gat));
  INV_X1    g704(.A(G162gat), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n898), .A2(new_n906), .A3(new_n627), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n880), .A2(new_n684), .A3(new_n875), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n707), .A2(new_n644), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n247), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n822), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n554), .A3(new_n666), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(G169gat), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n826), .A2(new_n910), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n822), .A2(new_n249), .A3(new_n730), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT123), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n915), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1348gat));
  NOR2_X1   g721(.A1(new_n783), .A2(new_n250), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n822), .A2(new_n606), .A3(new_n916), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n913), .A2(new_n923), .B1(new_n924), .B2(new_n250), .ZN(G1349gat));
  NAND3_X1  g724(.A1(new_n913), .A2(new_n666), .A3(new_n640), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G183gat), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n822), .A2(new_n289), .A3(new_n640), .A4(new_n916), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1350gat));
  NAND4_X1  g733(.A1(new_n822), .A2(new_n666), .A3(new_n684), .A4(new_n912), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n936), .A3(G190gat), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(KEYINPUT126), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(KEYINPUT126), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n935), .A2(G190gat), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n938), .B(new_n939), .C1(new_n936), .C2(new_n940), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n822), .A2(new_n275), .A3(new_n684), .A4(new_n916), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT125), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1351gat));
  AND2_X1   g743(.A1(new_n887), .A2(new_n890), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n668), .A2(new_n911), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n552), .ZN(new_n948));
  INV_X1    g747(.A(new_n946), .ZN(new_n949));
  NOR4_X1   g748(.A1(new_n886), .A2(G197gat), .A3(new_n696), .A4(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT127), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n948), .A2(new_n951), .ZN(G1352gat));
  NAND3_X1  g751(.A1(new_n945), .A2(new_n606), .A3(new_n946), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NOR4_X1   g753(.A1(new_n886), .A2(G204gat), .A3(new_n607), .A4(new_n949), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1353gat));
  NOR2_X1   g756(.A1(new_n886), .A2(new_n949), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n208), .A3(new_n640), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n887), .A2(new_n890), .A3(new_n640), .A4(new_n946), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  AOI21_X1  g762(.A(G218gat), .B1(new_n958), .B2(new_n684), .ZN(new_n964));
  INV_X1    g763(.A(new_n947), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n627), .A2(new_n209), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(G1355gat));
endmodule


