//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1308, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n215), .B1(new_n202), .B2(new_n216), .C1(new_n203), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n208), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n208), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n225), .B(new_n231), .C1(KEYINPUT1), .C2(new_n219), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n221), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n216), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n213), .ZN(new_n240));
  INV_X1    g0040(.A(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n237), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G169), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n216), .A2(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n252), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G97), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  AND2_X1   g0069(.A1(G1), .A2(G13), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(new_n263), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n268), .A2(G238), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n261), .A2(new_n262), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n264), .B1(new_n257), .B2(new_n258), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(new_n264), .A3(G274), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(new_n217), .B2(new_n267), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT13), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n251), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT14), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n276), .A2(new_n280), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT75), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n281), .A2(new_n286), .A3(new_n282), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n262), .B1(new_n261), .B2(new_n275), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT13), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n282), .B(G169), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT75), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n285), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT74), .B1(new_n294), .B2(new_n203), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT12), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n228), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n265), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n229), .A2(G33), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G77), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n303), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT11), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n292), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n283), .A2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n314), .B(new_n311), .C1(new_n315), .C2(new_n283), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n299), .A2(G50), .A3(new_n300), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(G50), .B2(new_n293), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT8), .B(G58), .Z(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(new_n305), .B1(G150), .B2(new_n307), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n204), .A2(G20), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n303), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT9), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n254), .A2(G222), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G223), .A2(G1698), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n252), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n328), .B(new_n260), .C1(G77), .C2(new_n252), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(new_n278), .C1(new_n253), .C2(new_n267), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT71), .B(G200), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n315), .B2(new_n330), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(KEYINPUT73), .C1(new_n315), .C2(new_n330), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT10), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n336), .B(new_n335), .C1(new_n325), .C2(new_n333), .ZN(new_n339));
  INV_X1    g0139(.A(new_n324), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n330), .A2(new_n251), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n340), .B(new_n341), .C1(G179), .C2(new_n330), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT15), .B(G87), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT70), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n305), .ZN(new_n348));
  INV_X1    g0148(.A(new_n307), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT69), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT69), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n307), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n320), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G20), .A2(G77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n303), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n300), .A2(G77), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n299), .A2(new_n359), .B1(new_n210), .B2(new_n294), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G33), .ZN(new_n364));
  INV_X1    g0164(.A(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G238), .A2(G1698), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n216), .B2(G1698), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n260), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT68), .B(G107), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n370), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n278), .B1(new_n211), .B2(new_n267), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n251), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n344), .B1(new_n362), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n373), .A2(new_n374), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n284), .ZN(new_n379));
  OAI211_X1 g0179(.A(KEYINPUT72), .B(new_n375), .C1(new_n357), .C2(new_n361), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(G190), .ZN(new_n382));
  INV_X1    g0182(.A(new_n331), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n362), .B(new_n382), .C1(new_n383), .C2(new_n378), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n343), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT76), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n365), .B2(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n363), .A2(KEYINPUT76), .A3(G33), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n366), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n253), .A2(G1698), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(G223), .B2(G1698), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n390), .A2(new_n392), .B1(new_n365), .B2(new_n212), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n260), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n278), .B1(new_n216), .B2(new_n267), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n315), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n260), .B2(new_n393), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(G200), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n320), .A2(new_n300), .ZN(new_n400));
  INV_X1    g0200(.A(new_n320), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n400), .A2(new_n299), .B1(new_n294), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n202), .A2(new_n203), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G58), .A2(G68), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n307), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n390), .A2(new_n229), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n203), .B1(new_n409), .B2(KEYINPUT7), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n390), .A2(new_n411), .A3(new_n229), .ZN(new_n412));
  AOI211_X1 g0212(.A(new_n403), .B(new_n408), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n252), .B2(G20), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n367), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n408), .B1(new_n416), .B2(G68), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n298), .B1(new_n417), .B2(KEYINPUT16), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n399), .B(new_n402), .C1(new_n413), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n420));
  INV_X1    g0220(.A(new_n402), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n252), .A2(new_n411), .A3(G20), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT7), .B1(new_n367), .B2(new_n229), .ZN(new_n423));
  OAI21_X1  g0223(.A(G68), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n408), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n303), .B1(new_n426), .B2(new_n403), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n409), .A2(KEYINPUT7), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(G68), .A3(new_n412), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n421), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n399), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n420), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n398), .A2(G179), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n251), .B2(new_n398), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT18), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n402), .B1(new_n413), .B2(new_n418), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n436), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n317), .A2(new_n386), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n388), .A2(new_n389), .A3(new_n229), .A4(new_n366), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT22), .B1(new_n446), .B2(new_n212), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT87), .B(KEYINPUT22), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n252), .A2(new_n448), .A3(new_n229), .A4(G87), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n229), .A2(KEYINPUT23), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G116), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n451), .A2(G107), .B1(G20), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n372), .A2(G20), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(KEYINPUT23), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT24), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n450), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n303), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT88), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT25), .ZN(new_n462));
  AOI211_X1 g0262(.A(G107), .B(new_n293), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n461), .A2(new_n462), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n265), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n293), .A2(new_n467), .A3(new_n228), .A4(new_n297), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n465), .A2(new_n466), .B1(G107), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G41), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n265), .A2(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n476), .B2(KEYINPUT80), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n265), .B(G45), .C1(new_n272), .C2(KEYINPUT5), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n477), .A2(KEYINPUT81), .A3(new_n271), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n472), .A2(G41), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n482), .A2(KEYINPUT80), .A3(new_n265), .A4(G45), .ZN(new_n483));
  INV_X1    g0283(.A(new_n473), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n480), .A2(new_n483), .A3(new_n271), .A4(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  MUX2_X1   g0288(.A(new_n213), .B(new_n241), .S(G1698), .Z(new_n489));
  INV_X1    g0289(.A(G294), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n390), .A2(new_n489), .B1(new_n365), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n260), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n483), .A2(new_n484), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n478), .A2(new_n479), .ZN(new_n494));
  OAI211_X1 g0294(.A(G264), .B(new_n264), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n488), .A2(new_n496), .A3(new_n284), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n492), .A2(new_n495), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n481), .A2(new_n487), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n251), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n460), .A2(new_n471), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n450), .A2(new_n458), .A3(new_n455), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n458), .B1(new_n450), .B2(new_n455), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n298), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n488), .A2(new_n496), .A3(G190), .ZN(new_n505));
  AOI21_X1  g0305(.A(G200), .B1(new_n498), .B2(new_n499), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n504), .B(new_n470), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G264), .A2(G1698), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n241), .B2(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n511), .A2(new_n388), .A3(new_n366), .A4(new_n389), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n367), .A2(G303), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT85), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n260), .A3(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G270), .B(new_n264), .C1(new_n493), .C2(new_n494), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n499), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n229), .C1(G33), .C2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n298), .C1(new_n229), .C2(G116), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n294), .A2(KEYINPUT86), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT86), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n293), .B2(G116), .ZN(new_n530));
  AOI22_X1  g0330(.A1(G116), .A2(new_n469), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n520), .A2(G169), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n260), .B1(new_n477), .B2(new_n480), .ZN(new_n536));
  AOI22_X1  g0336(.A1(G270), .A2(new_n536), .B1(new_n481), .B2(new_n487), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n537), .A2(new_n532), .A3(G179), .A4(new_n518), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n520), .A2(KEYINPUT21), .A3(G169), .A4(new_n532), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n532), .B1(new_n520), .B2(G200), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n315), .B2(new_n520), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT19), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n258), .B2(new_n229), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n212), .A2(new_n522), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n371), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n544), .B1(new_n304), .B2(new_n522), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n446), .A2(new_n203), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n298), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n345), .B(KEYINPUT70), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n294), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n347), .A2(new_n469), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n213), .B1(new_n273), .B2(G1), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n265), .A2(new_n269), .A3(G45), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n264), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT83), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n264), .A2(new_n556), .A3(new_n557), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G244), .A2(G1698), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n217), .B2(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(new_n388), .A3(new_n366), .A4(new_n389), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n264), .B1(new_n565), .B2(new_n452), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n284), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n251), .B1(new_n562), .B2(new_n566), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n555), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n547), .B(new_n548), .C1(new_n203), .C2(new_n446), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n298), .B1(new_n294), .B2(new_n552), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n559), .A2(new_n561), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n565), .A2(new_n452), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n260), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(G190), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n469), .A2(G87), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n331), .B1(new_n562), .B2(new_n566), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n572), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n570), .A2(new_n579), .A3(KEYINPUT84), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT84), .B1(new_n570), .B2(new_n579), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n372), .B1(new_n414), .B2(new_n415), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g0384(.A(G97), .B(G107), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n586), .A2(new_n522), .A3(G107), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G20), .B1(G77), .B2(new_n307), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n468), .A2(G97), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G97), .B2(new_n294), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT77), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n593), .B(KEYINPUT77), .C1(G97), .C2(new_n294), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n592), .A2(new_n298), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G257), .B(new_n264), .C1(new_n493), .C2(new_n494), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n499), .A2(new_n284), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n521), .B1(new_n367), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(G250), .A2(G1698), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n364), .A2(new_n366), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT78), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT78), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n252), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n603), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT4), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n254), .A2(G244), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n390), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT79), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n606), .A2(new_n608), .ZN(new_n614));
  INV_X1    g0414(.A(new_n602), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n252), .A2(new_n615), .B1(G33), .B2(G283), .ZN(new_n616));
  AND4_X1   g0416(.A1(KEYINPUT79), .A2(new_n614), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n260), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n598), .B1(new_n601), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n614), .A2(new_n612), .A3(new_n616), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT79), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n614), .A2(new_n612), .A3(KEYINPUT79), .A4(new_n616), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n264), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n499), .A2(new_n599), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n251), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(G200), .B1(new_n624), .B2(new_n625), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n624), .A2(new_n315), .A3(new_n625), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n598), .B(new_n628), .C1(new_n629), .C2(KEYINPUT82), .ZN(new_n630));
  INV_X1    g0430(.A(new_n625), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n618), .A2(new_n631), .A3(KEYINPUT82), .A4(G190), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n582), .B(new_n627), .C1(new_n630), .C2(new_n633), .ZN(new_n634));
  NOR4_X1   g0434(.A1(new_n445), .A2(new_n509), .A3(new_n543), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n342), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT92), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n380), .A2(new_n379), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n552), .A2(new_n304), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n298), .B1(new_n639), .B2(new_n355), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n360), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT72), .B1(new_n641), .B2(new_n375), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n637), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n377), .A2(KEYINPUT92), .A3(new_n379), .A4(new_n380), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n643), .A2(new_n644), .A3(new_n316), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n434), .B1(new_n645), .B2(new_n312), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n439), .A2(new_n440), .A3(new_n436), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n440), .B1(new_n439), .B2(new_n436), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n338), .A2(new_n339), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n636), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n566), .A2(KEYINPUT89), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n566), .A2(KEYINPUT89), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n573), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n331), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(new_n572), .A3(new_n577), .A4(new_n576), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n251), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n555), .A3(new_n568), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT82), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n618), .A2(new_n631), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n315), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(new_n598), .A3(new_n632), .A4(new_n628), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n501), .A2(new_n535), .A3(new_n538), .A4(new_n539), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n507), .A4(new_n627), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT91), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n619), .A2(new_n667), .A3(new_n626), .ZN(new_n668));
  AOI21_X1  g0468(.A(G169), .B1(new_n618), .B2(new_n631), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n596), .A2(new_n597), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n588), .B1(new_n586), .B2(new_n585), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n671), .A2(new_n229), .B1(new_n210), .B2(new_n349), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n298), .B1(new_n672), .B2(new_n583), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n624), .B2(new_n600), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT91), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n660), .B1(new_n666), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n659), .B(KEYINPUT90), .Z(new_n681));
  NAND2_X1  g0481(.A1(new_n570), .A2(new_n579), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT84), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n570), .A2(new_n579), .A3(KEYINPUT84), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n626), .A4(new_n619), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n652), .B1(new_n690), .B2(new_n445), .ZN(G369));
  INV_X1    g0491(.A(new_n540), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n265), .A2(new_n229), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n526), .B2(new_n531), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n692), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n543), .B2(new_n700), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n501), .A2(new_n699), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT93), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n698), .B1(new_n460), .B2(new_n471), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n508), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT94), .Z(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n540), .A2(new_n698), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n501), .A2(new_n698), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(G399));
  NOR3_X1   g0517(.A1(new_n371), .A2(G116), .A3(new_n546), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n222), .A2(new_n272), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n226), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n723), .B(new_n699), .C1(new_n680), .C2(new_n688), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n659), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n677), .A2(new_n727), .B1(new_n686), .B2(new_n678), .ZN(new_n728));
  INV_X1    g0528(.A(new_n681), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT96), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n669), .A2(new_n675), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n624), .A2(new_n625), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT82), .B1(new_n732), .B2(G190), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n628), .A2(new_n598), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n731), .B1(new_n735), .B2(new_n632), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n660), .B1(new_n540), .B2(new_n501), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT97), .A4(new_n507), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT97), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n664), .A2(new_n507), .A3(new_n627), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n665), .A2(new_n659), .A3(new_n657), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT96), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n726), .B1(new_n676), .B2(new_n668), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT26), .B1(new_n582), .B2(new_n731), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n743), .B(new_n681), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n730), .A2(new_n738), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n699), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n725), .B1(new_n748), .B2(KEYINPUT29), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n567), .A2(new_n495), .A3(new_n492), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n618), .A2(new_n631), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n518), .A2(new_n499), .A3(G179), .A4(new_n519), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT95), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n537), .A2(KEYINPUT95), .A3(G179), .A4(new_n518), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(G179), .B1(new_n498), .B2(new_n499), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n520), .A3(new_n655), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT30), .B1(new_n760), .B2(new_n732), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n698), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n756), .A2(new_n757), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT30), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n763), .A2(new_n764), .A3(new_n732), .A4(new_n752), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n750), .B1(new_n762), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n624), .A2(new_n625), .A3(new_n751), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n662), .A2(new_n520), .A3(new_n655), .A4(new_n759), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(KEYINPUT30), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n771), .A2(KEYINPUT31), .A3(new_n698), .A4(new_n765), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n508), .A2(new_n540), .A3(new_n542), .A4(new_n699), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n767), .B(new_n772), .C1(new_n634), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G330), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n749), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n722), .B1(new_n776), .B2(G1), .ZN(G364));
  AND2_X1   g0577(.A1(new_n229), .A2(G13), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n265), .B1(new_n778), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n719), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n703), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G330), .B2(new_n702), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n252), .A2(new_n222), .ZN(new_n785));
  INV_X1    g0585(.A(G355), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n786), .B1(G116), .B2(new_n222), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n246), .A2(G45), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n390), .A2(new_n222), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n273), .B2(new_n227), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n228), .B1(G20), .B2(new_n251), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n782), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(G20), .A2(G179), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT98), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n315), .ZN(new_n801));
  INV_X1    g0601(.A(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n801), .A2(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n203), .A2(new_n804), .B1(new_n806), .B2(new_n210), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n800), .A2(G190), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G200), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(G58), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n229), .A2(G179), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n331), .A2(new_n315), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(G107), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n331), .A2(G190), .A3(new_n811), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G87), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n815), .A2(new_n252), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G179), .A2(G200), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(G20), .A3(new_n315), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G159), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT32), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT99), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n808), .A2(new_n802), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n229), .B1(new_n820), .B2(G190), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT100), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n826), .A2(G50), .B1(new_n828), .B2(G97), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n810), .A2(new_n819), .A3(new_n825), .A4(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G311), .A2(new_n805), .B1(new_n809), .B2(G322), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT33), .B(G317), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n803), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n252), .B1(new_n822), .B2(G329), .ZN(new_n834));
  INV_X1    g0634(.A(G283), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n812), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G303), .B2(new_n817), .ZN(new_n837));
  XOR2_X1   g0637(.A(KEYINPUT101), .B(G326), .Z(new_n838));
  AOI22_X1  g0638(.A1(new_n826), .A2(new_n838), .B1(new_n828), .B2(G294), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n831), .A2(new_n833), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n830), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n798), .B1(new_n841), .B2(new_n795), .ZN(new_n842));
  INV_X1    g0642(.A(new_n794), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n702), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n784), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G396));
  NAND2_X1  g0646(.A1(new_n641), .A2(new_n698), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n643), .A2(new_n644), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n384), .B(new_n847), .C1(new_n638), .C2(new_n642), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT103), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT103), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n381), .A2(new_n852), .A3(new_n384), .A4(new_n847), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n849), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n690), .B2(new_n698), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n698), .B1(new_n851), .B2(new_n853), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n680), .B2(new_n688), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n782), .B1(new_n858), .B2(new_n775), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n855), .A2(G330), .A3(new_n774), .A4(new_n857), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n795), .A2(new_n792), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT102), .Z(new_n863));
  OAI21_X1  g0663(.A(new_n782), .B1(new_n863), .B2(G77), .ZN(new_n864));
  INV_X1    g0664(.A(new_n826), .ZN(new_n865));
  INV_X1    g0665(.A(G303), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n835), .A2(new_n804), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(G116), .B2(new_n805), .ZN(new_n868));
  INV_X1    g0668(.A(G311), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n367), .B1(new_n821), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n812), .A2(new_n212), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n870), .B(new_n871), .C1(G107), .C2(new_n817), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n809), .A2(G294), .B1(new_n828), .B2(G97), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G137), .A2(new_n826), .B1(new_n803), .B2(G150), .ZN(new_n875));
  INV_X1    g0675(.A(G143), .ZN(new_n876));
  INV_X1    g0676(.A(new_n809), .ZN(new_n877));
  INV_X1    g0677(.A(G159), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n875), .B1(new_n876), .B2(new_n877), .C1(new_n878), .C2(new_n806), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT34), .Z(new_n880));
  AOI21_X1  g0680(.A(new_n390), .B1(G132), .B2(new_n822), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n201), .B2(new_n816), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n812), .A2(new_n203), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n828), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n202), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n874), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n864), .B1(new_n887), .B2(new_n795), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n849), .A2(new_n851), .A3(new_n853), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n793), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n861), .A2(new_n890), .ZN(G384));
  OR2_X1    g0691(.A1(new_n590), .A2(KEYINPUT35), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n590), .A2(KEYINPUT35), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(G116), .A3(new_n230), .A4(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT36), .Z(new_n895));
  OAI211_X1 g0695(.A(new_n227), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n201), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n265), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n652), .B1(new_n749), .B2(new_n445), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n313), .A2(new_n698), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n431), .A2(new_n696), .ZN(new_n902));
  INV_X1    g0702(.A(new_n696), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n439), .B1(new_n436), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n419), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n427), .A2(new_n430), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n437), .A2(new_n696), .B1(new_n906), .B2(new_n402), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT105), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n442), .A2(new_n902), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n904), .A2(new_n908), .A3(KEYINPUT37), .A4(new_n419), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n430), .A2(new_n298), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT16), .B1(new_n429), .B2(new_n425), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n402), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n903), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n649), .B2(new_n434), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n436), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT37), .A4(new_n419), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT37), .ZN(new_n920));
  INV_X1    g0720(.A(new_n419), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n907), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n917), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n912), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n924), .B1(new_n917), .B2(new_n923), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n429), .A2(new_n425), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n403), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n430), .A3(new_n298), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n696), .B1(new_n931), .B2(new_n402), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n442), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n419), .A2(KEYINPUT37), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n935), .A2(new_n918), .B1(new_n905), .B2(new_n920), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n936), .A3(KEYINPUT38), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n927), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n901), .B1(new_n926), .B2(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n381), .A2(new_n698), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n857), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n928), .A2(new_n937), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n311), .A2(new_n699), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n316), .B(new_n944), .C1(new_n292), .C2(new_n311), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT104), .B1(new_n292), .B2(new_n944), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT104), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n291), .A2(new_n287), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n947), .B(new_n943), .C1(new_n948), .C2(new_n285), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n941), .A2(new_n942), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n649), .A2(new_n903), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n939), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n900), .B(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(G330), .ZN(new_n956));
  XNOR2_X1  g0756(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n950), .A2(new_n889), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n772), .B1(new_n773), .B2(new_n634), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT107), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n762), .B2(new_n766), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n771), .A2(KEYINPUT107), .A3(new_n698), .A4(new_n765), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n750), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n958), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n957), .B1(new_n965), .B2(new_n942), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT40), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n420), .A2(new_n433), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n438), .A2(new_n441), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n902), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n909), .A2(new_n905), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n911), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n924), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n967), .B1(new_n973), .B2(new_n937), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n966), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n445), .B1(new_n960), .B2(new_n964), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n956), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n975), .B2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n955), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n265), .B2(new_n778), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n955), .A2(new_n978), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n899), .B1(new_n980), .B2(new_n981), .ZN(G367));
  INV_X1    g0782(.A(new_n242), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n796), .B1(new_n222), .B2(new_n552), .C1(new_n983), .C2(new_n789), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n984), .A2(new_n782), .ZN(new_n985));
  INV_X1    g0785(.A(new_n795), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n805), .A2(G283), .B1(new_n828), .B2(new_n371), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT113), .ZN(new_n988));
  INV_X1    g0788(.A(G317), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n390), .B1(new_n989), .B2(new_n821), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n812), .A2(new_n522), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(new_n826), .C2(G311), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n817), .A2(G116), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT46), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G294), .A2(new_n803), .B1(new_n809), .B2(G303), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n812), .A2(new_n210), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n367), .B(new_n997), .C1(G137), .C2(new_n822), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G150), .A2(new_n809), .B1(new_n803), .B2(G159), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n202), .C2(new_n816), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n828), .A2(G68), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n806), .B2(new_n201), .C1(new_n876), .C2(new_n865), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n988), .A2(new_n996), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT47), .Z(new_n1004));
  AOI21_X1  g0804(.A(new_n699), .B1(new_n572), .B2(new_n577), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT108), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n729), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n660), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n985), .B1(new_n986), .B2(new_n1004), .C1(new_n1009), .C2(new_n843), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n708), .B(new_n712), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(new_n703), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n776), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n736), .B1(new_n598), .B2(new_n699), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n731), .A2(new_n698), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1017), .A2(KEYINPUT110), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(KEYINPUT110), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n716), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT45), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n715), .ZN(new_n1023));
  XOR2_X1   g0823(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n715), .A3(new_n1024), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1021), .A2(new_n1028), .A3(new_n711), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT45), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1020), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1027), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1024), .B1(new_n1022), .B2(new_n715), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n710), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1014), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n776), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n719), .B(KEYINPUT41), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n780), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1009), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT43), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT109), .Z(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n627), .B1(new_n1022), .B2(new_n501), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n713), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1046), .A2(new_n699), .B1(KEYINPUT42), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT42), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n1047), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT111), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1045), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1044), .B(new_n1054), .C1(new_n1049), .C2(new_n1052), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n711), .A2(new_n1022), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1056), .A2(new_n1058), .B1(new_n711), .B2(new_n1022), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1010), .B1(new_n1040), .B2(new_n1063), .ZN(G387));
  NAND3_X1  g0864(.A1(new_n705), .A2(new_n707), .A3(new_n794), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n718), .A2(new_n785), .B1(G107), .B2(new_n222), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n237), .A2(G45), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n718), .ZN(new_n1068));
  AOI211_X1 g0868(.A(G45), .B(new_n1068), .C1(G68), .C2(G77), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n320), .A2(new_n201), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT50), .Z(new_n1071));
  AOI21_X1  g0871(.A(new_n789), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1066), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n782), .B1(new_n1073), .B2(new_n797), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n878), .A2(new_n865), .B1(new_n804), .B2(new_n401), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G68), .B2(new_n805), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n390), .B(new_n991), .C1(G150), .C2(new_n822), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n817), .A2(G77), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n809), .A2(G50), .B1(new_n828), .B2(new_n347), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n390), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n822), .B2(new_n838), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n885), .A2(new_n835), .B1(new_n490), .B2(new_n816), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G311), .A2(new_n803), .B1(new_n826), .B2(G322), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n866), .B2(new_n806), .C1(new_n989), .C2(new_n877), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT48), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT49), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1082), .B1(new_n527), .B2(new_n812), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1080), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1074), .B1(new_n1092), .B2(new_n795), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1012), .A2(new_n780), .B1(new_n1065), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1013), .A2(new_n781), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n776), .A2(new_n1012), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(G393));
  INV_X1    g0897(.A(new_n1035), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1031), .A2(new_n1034), .A3(new_n710), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n1013), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(new_n781), .A3(new_n1036), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n796), .B1(new_n522), .B2(new_n222), .C1(new_n249), .C2(new_n789), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1081), .B1(new_n876), .B2(new_n821), .C1(new_n812), .C2(new_n212), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n803), .A2(G50), .B1(new_n828), .B2(G77), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n401), .B2(new_n806), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G68), .C2(new_n817), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G150), .A2(new_n826), .B1(new_n809), .B2(G159), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT51), .Z(new_n1108));
  AOI21_X1  g0908(.A(new_n252), .B1(new_n822), .B2(G322), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n815), .B(new_n1109), .C1(new_n835), .C2(new_n816), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n490), .A2(new_n806), .B1(new_n804), .B2(new_n866), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G116), .C2(new_n828), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G311), .A2(new_n809), .B1(new_n826), .B2(G317), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT52), .Z(new_n1114));
  AOI22_X1  g0914(.A1(new_n1106), .A2(new_n1108), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n782), .B(new_n1102), .C1(new_n1115), .C2(new_n986), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1022), .B2(new_n794), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n780), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1101), .A2(new_n1119), .ZN(G390));
  NAND2_X1  g0920(.A1(new_n942), .A2(KEYINPUT39), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n973), .A2(new_n927), .A3(new_n937), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n857), .B2(new_n940), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1121), .B(new_n1122), .C1(new_n1124), .C2(new_n901), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n747), .A2(new_n699), .A3(new_n889), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1123), .B1(new_n1126), .B2(new_n940), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n912), .A2(new_n925), .B1(new_n313), .B2(new_n698), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n956), .B(new_n958), .C1(new_n960), .C2(new_n964), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n774), .A2(G330), .A3(new_n889), .A4(new_n950), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1125), .B(new_n1132), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1133), .A3(new_n780), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n522), .A2(new_n806), .B1(new_n877), .B2(new_n527), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G283), .B2(new_n826), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n818), .B(new_n367), .C1(new_n490), .C2(new_n821), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1137), .A2(new_n883), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n803), .A2(new_n371), .B1(new_n828), .B2(G77), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n817), .A2(G150), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT53), .Z(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT54), .B(G143), .Z(new_n1143));
  AOI22_X1  g0943(.A1(G137), .A2(new_n803), .B1(new_n805), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n809), .A2(G132), .B1(new_n828), .B2(G159), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n367), .B1(new_n822), .B2(G125), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n201), .B2(new_n812), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n826), .B2(G128), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n986), .B1(new_n1140), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n782), .B1(new_n863), .B2(new_n320), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n793), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1134), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n956), .B1(new_n960), .B2(new_n964), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n958), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n761), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n699), .B1(new_n1158), .B2(new_n769), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT31), .B1(new_n1159), .B2(new_n765), .ZN(new_n1160));
  OAI211_X1 g0960(.A(G330), .B(new_n889), .C1(new_n959), .C2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1156), .A2(new_n1157), .B1(new_n1161), .B2(new_n1123), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n941), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT114), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT114), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1161), .A2(new_n1123), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1165), .B(new_n941), .C1(new_n1166), .C2(new_n1130), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1126), .A2(new_n940), .A3(new_n1132), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n962), .A2(new_n750), .A3(new_n963), .ZN(new_n1170));
  OAI211_X1 g0970(.A(G330), .B(new_n889), .C1(new_n1170), .C2(new_n959), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1123), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT115), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1171), .A2(KEYINPUT115), .A3(new_n1123), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1169), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1168), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1156), .A2(new_n444), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n652), .B(new_n1178), .C1(new_n749), .C2(new_n445), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n719), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1177), .A2(new_n1131), .A3(new_n1180), .A4(new_n1133), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1155), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G378));
  NAND3_X1  g0986(.A1(new_n1126), .A2(new_n940), .A3(new_n1132), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT115), .B1(new_n1171), .B2(new_n1123), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1189), .A2(new_n1175), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1180), .B1(new_n1182), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n956), .B1(new_n974), .B2(new_n965), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n942), .B(new_n1157), .C1(new_n1170), .C2(new_n959), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n957), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n343), .A2(KEYINPUT118), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT118), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n338), .A2(new_n1199), .A3(new_n339), .A4(new_n342), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1198), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1202), .A2(new_n1203), .B1(new_n324), .B2(new_n696), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1203), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n324), .A2(new_n696), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1201), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1192), .A2(new_n1195), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n954), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1157), .B1(new_n1170), .B2(new_n959), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT40), .B1(new_n912), .B2(new_n925), .ZN(new_n1214));
  OAI21_X1  g1014(.A(G330), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1212), .B1(new_n1215), .B2(new_n966), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n952), .B1(new_n1153), .B2(new_n901), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1192), .A2(new_n1195), .A3(new_n1208), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1216), .A2(new_n951), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1191), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT57), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n719), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1184), .A2(new_n1180), .B1(new_n1219), .B2(new_n1211), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT57), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n781), .B(new_n780), .C1(new_n201), .C2(new_n862), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n805), .A2(G137), .B1(new_n817), .B2(new_n1143), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G128), .A2(new_n809), .B1(new_n803), .B2(G132), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n826), .A2(G125), .B1(new_n828), .B2(G150), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT116), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1228), .B(new_n1229), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(KEYINPUT59), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT117), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(G124), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(G124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n822), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n365), .A3(new_n272), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G159), .B2(new_n813), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1235), .A2(new_n1236), .A3(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1078), .B1(new_n835), .B2(new_n821), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n390), .A2(new_n272), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n812), .A2(new_n202), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(new_n1001), .C1(new_n527), .C2(new_n865), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G107), .A2(new_n809), .B1(new_n805), .B2(new_n347), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n522), .B2(new_n804), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT58), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1245), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1251), .A2(KEYINPUT58), .ZN(new_n1254));
  AND4_X1   g1054(.A1(new_n1243), .A2(new_n1252), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1227), .B1(new_n986), .B2(new_n1255), .C1(new_n1208), .C2(new_n793), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT119), .Z(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1220), .A2(new_n780), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1226), .A2(new_n1261), .ZN(G375));
  NAND2_X1  g1062(.A1(new_n1123), .A2(new_n792), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n782), .B1(new_n863), .B2(G68), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n527), .A2(new_n804), .B1(new_n806), .B2(new_n372), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G283), .B2(new_n809), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n367), .B1(new_n821), .B2(new_n866), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1267), .B(new_n997), .C1(G97), .C2(new_n817), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n826), .A2(G294), .B1(new_n828), .B2(new_n347), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G132), .A2(new_n826), .B1(new_n809), .B2(G137), .ZN(new_n1271));
  INV_X1    g1071(.A(G128), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1081), .B1(new_n1272), .B2(new_n821), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1246), .B(new_n1273), .C1(G159), .C2(new_n817), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(G150), .A2(new_n805), .B1(new_n803), .B2(new_n1143), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n828), .A2(G50), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1271), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1270), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1264), .B1(new_n1278), .B2(new_n795), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1263), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1190), .B2(new_n779), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1168), .A2(new_n1176), .A3(new_n1179), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT120), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1190), .A2(KEYINPUT120), .A3(new_n1179), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1181), .A2(new_n1039), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1282), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT121), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(G381));
  INV_X1    g1093(.A(G390), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1038), .B1(new_n1036), .B2(new_n776), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1061), .B(new_n1062), .C1(new_n1295), .C2(new_n780), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1296), .A3(new_n1010), .ZN(new_n1297));
  OR2_X1    g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1297), .A2(G384), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1292), .A3(new_n1291), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT122), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT122), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1299), .A2(new_n1302), .A3(new_n1292), .A4(new_n1291), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1226), .A2(new_n1185), .A3(new_n1261), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1301), .A2(new_n1303), .A3(new_n1305), .ZN(G407));
  INV_X1    g1106(.A(G213), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1305), .B2(new_n697), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(G407), .A2(new_n1308), .ZN(G409));
  OAI21_X1  g1109(.A(KEYINPUT60), .B1(new_n1190), .B2(new_n1179), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1168), .A2(new_n1176), .A3(new_n1179), .A4(KEYINPUT60), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1312), .A2(new_n781), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1282), .ZN(new_n1315));
  INV_X1    g1115(.A(G384), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1314), .A2(G384), .A3(new_n1282), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(KEYINPUT125), .A3(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G384), .B1(new_n1314), .B2(new_n1282), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1316), .B(new_n1281), .C1(new_n1311), .C2(new_n1313), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1320), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1191), .A2(new_n1039), .A3(new_n1220), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n779), .B1(new_n1220), .B2(KEYINPUT123), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT123), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1211), .A2(new_n1219), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1257), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT124), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1325), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1209), .A2(new_n1210), .A3(new_n954), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1216), .A2(new_n1218), .B1(new_n951), .B2(new_n1217), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT123), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(new_n780), .A3(new_n1328), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1258), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1336), .A2(KEYINPUT124), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1185), .B1(new_n1331), .B2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n781), .B1(new_n1224), .B2(KEYINPUT57), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1340));
  OAI211_X1 g1140(.A(G378), .B(new_n1261), .C1(new_n1339), .C2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1338), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n697), .A2(G213), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1324), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(KEYINPUT62), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n697), .A2(G213), .A3(G2897), .ZN(new_n1346));
  AOI21_X1  g1146(.A(KEYINPUT125), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1321), .A2(new_n1322), .A3(new_n1320), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1346), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  AOI211_X1 g1149(.A(new_n1185), .B(new_n1260), .C1(new_n1223), .C2(new_n1225), .ZN(new_n1350));
  AOI22_X1  g1150(.A1(new_n1336), .A2(KEYINPUT124), .B1(new_n1039), .B2(new_n1224), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1352));
  AOI21_X1  g1152(.A(G378), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1343), .B1(new_n1350), .B2(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1346), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1349), .A2(new_n1354), .A3(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT61), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1324), .A2(new_n1342), .A3(new_n1359), .A4(new_n1343), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1345), .A2(new_n1357), .A3(new_n1358), .A4(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(G387), .A2(G390), .ZN(new_n1362));
  AOI21_X1  g1162(.A(KEYINPUT126), .B1(new_n1362), .B2(new_n1297), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1363), .ZN(new_n1364));
  XNOR2_X1  g1164(.A(G393), .B(new_n845), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(G390), .A2(KEYINPUT126), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1365), .B1(G387), .B2(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT127), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(G387), .A2(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1365), .B1(new_n1370), .B2(G390), .ZN(new_n1371));
  AOI21_X1  g1171(.A(KEYINPUT127), .B1(new_n1296), .B2(new_n1010), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1372), .A2(new_n1294), .ZN(new_n1373));
  AOI22_X1  g1173(.A1(new_n1364), .A2(new_n1368), .B1(new_n1371), .B2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1361), .A2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1344), .A2(KEYINPUT63), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT63), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1324), .A2(new_n1342), .A3(new_n1377), .A4(new_n1343), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1376), .A2(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1365), .ZN(new_n1380));
  OAI21_X1  g1180(.A(new_n1380), .B1(new_n1372), .B2(new_n1294), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1370), .A2(G390), .ZN(new_n1382));
  OAI22_X1  g1182(.A1(new_n1363), .A2(new_n1367), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1355), .B1(new_n1324), .B2(new_n1346), .ZN(new_n1384));
  AOI21_X1  g1184(.A(KEYINPUT61), .B1(new_n1384), .B2(new_n1354), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1379), .A2(new_n1383), .A3(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1375), .A2(new_n1386), .ZN(G405));
  NAND2_X1  g1187(.A1(G375), .A2(new_n1185), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1388), .A2(new_n1341), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1389), .A2(new_n1324), .ZN(new_n1390));
  OAI211_X1 g1190(.A(new_n1388), .B(new_n1341), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1390), .A2(new_n1391), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1374), .A2(new_n1392), .ZN(new_n1393));
  NAND3_X1  g1193(.A1(new_n1383), .A2(new_n1390), .A3(new_n1391), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1393), .A2(new_n1394), .ZN(G402));
endmodule


