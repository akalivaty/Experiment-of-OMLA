//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT66), .B(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI22_X1  g0021(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n212), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n206), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(KEYINPUT64), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g0036(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n239), .A2(new_n204), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n213), .A2(new_n211), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  OR2_X1    g0042(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n243), .A2(G50), .A3(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  AOI211_X1 g0046(.A(new_n209), .B(new_n233), .C1(new_n240), .C2(new_n246), .ZN(G361));
  XNOR2_X1  g0047(.A(KEYINPUT2), .B(G226), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G232), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G238), .B(G244), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G250), .B(G257), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(G264), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(new_n221), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G358));
  XOR2_X1   g0055(.A(G68), .B(G77), .Z(new_n256));
  XNOR2_X1  g0056(.A(G50), .B(G58), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(G87), .B(G97), .ZN(new_n259));
  XNOR2_X1  g0059(.A(G107), .B(G116), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n258), .B(new_n261), .Z(G351));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n203), .A2(G13), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n204), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n236), .A2(new_n237), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n203), .B2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n267), .B1(new_n271), .B2(new_n264), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT16), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT7), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n211), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G58), .A2(G68), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n204), .B1(new_n241), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n204), .A2(new_n277), .ZN(new_n286));
  INV_X1    g0086(.A(G159), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n273), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n269), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT76), .B1(new_n277), .B2(KEYINPUT3), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT76), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(new_n279), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n278), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(new_n274), .A3(new_n204), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n279), .A2(G33), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n294), .B2(new_n296), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT7), .B1(new_n301), .B2(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n299), .A2(G68), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n289), .A2(KEYINPUT77), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT77), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n285), .B2(new_n288), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n303), .A2(new_n307), .A3(KEYINPUT16), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n272), .B1(new_n293), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n310));
  INV_X1    g0110(.A(G274), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G41), .ZN(new_n313));
  OAI211_X1 g0113(.A(G1), .B(G13), .C1(new_n277), .C2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n314), .A2(new_n310), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n315), .B2(G232), .ZN(new_n316));
  AND2_X1   g0116(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G223), .ZN(new_n320));
  INV_X1    g0120(.A(G1698), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n319), .A2(new_n320), .B1(new_n219), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n301), .B1(G33), .B2(G87), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n236), .A2(new_n237), .B1(G33), .B2(G41), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n316), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G200), .ZN(new_n327));
  INV_X1    g0127(.A(new_n316), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n301), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n277), .B2(new_n224), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n330), .B2(new_n324), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G190), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n309), .A2(KEYINPUT17), .A3(new_n327), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n308), .A2(new_n269), .A3(new_n291), .ZN(new_n334));
  INV_X1    g0134(.A(new_n272), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n332), .A2(new_n334), .A3(new_n327), .A4(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT17), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n303), .A2(KEYINPUT16), .A3(new_n307), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n335), .B1(new_n339), .B2(new_n292), .ZN(new_n340));
  OAI211_X1 g0140(.A(G179), .B(new_n316), .C1(new_n323), .C2(new_n325), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(new_n331), .B2(new_n342), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n340), .A2(KEYINPUT18), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT18), .B1(new_n340), .B2(new_n343), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n333), .B(new_n338), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n275), .B1(new_n210), .B2(new_n321), .C1(new_n214), .C2(new_n319), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n324), .C1(G107), .C2(new_n275), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n312), .B1(new_n315), .B2(G244), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G200), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n270), .A2(G77), .ZN(new_n354));
  INV_X1    g0154(.A(new_n266), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(G77), .ZN(new_n356));
  INV_X1    g0156(.A(new_n286), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n264), .A2(new_n357), .B1(G20), .B2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n204), .A2(G33), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n356), .B1(new_n362), .B2(new_n269), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n269), .ZN(new_n365));
  INV_X1    g0165(.A(new_n356), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n354), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n349), .B2(new_n350), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT71), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n349), .A2(G190), .A3(new_n350), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n351), .A2(new_n342), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n349), .A2(new_n374), .A3(new_n350), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n367), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n347), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G222), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n275), .B1(new_n320), .B2(new_n321), .C1(new_n319), .C2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(G77), .B2(new_n275), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT69), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT69), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n380), .B(new_n383), .C1(G77), .C2(new_n275), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n324), .A3(new_n384), .ZN(new_n385));
  OR2_X1    g0185(.A1(KEYINPUT67), .A2(G226), .ZN(new_n386));
  NAND2_X1  g0186(.A1(KEYINPUT67), .A2(G226), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n315), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n312), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(G179), .ZN(new_n391));
  OAI21_X1  g0191(.A(G20), .B1(new_n241), .B2(G50), .ZN(new_n392));
  INV_X1    g0192(.A(G150), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n392), .B1(new_n393), .B2(new_n286), .C1(new_n361), .C2(new_n263), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n269), .B1(new_n270), .B2(G50), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(G50), .B2(new_n355), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n390), .A2(new_n342), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT10), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT9), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n385), .A2(G190), .A3(new_n388), .A4(new_n389), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT73), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n396), .A2(new_n400), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n390), .A2(G200), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT73), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n399), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n408), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n399), .A4(new_n406), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n401), .A2(new_n402), .A3(new_n399), .A4(new_n404), .ZN(new_n414));
  INV_X1    g0214(.A(new_n406), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT72), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n398), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(G226), .B1(new_n317), .B2(new_n318), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G232), .A2(G1698), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n281), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n277), .A2(new_n226), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n324), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n312), .B1(new_n315), .B2(G238), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n324), .B(KEYINPUT74), .C1(new_n421), .C2(new_n422), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT13), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n425), .A2(new_n430), .A3(new_n426), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G169), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(G179), .A3(new_n431), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n436), .A3(G169), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n211), .A2(G20), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n439), .B1(new_n361), .B2(new_n215), .C1(new_n218), .C2(new_n286), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n440), .A2(new_n269), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT11), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n441), .A2(KEYINPUT11), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n265), .A2(new_n439), .ZN(new_n444));
  XOR2_X1   g0244(.A(new_n444), .B(KEYINPUT12), .Z(new_n445));
  NAND2_X1  g0245(.A1(new_n270), .A2(G68), .ZN(new_n446));
  AND4_X1   g0246(.A1(new_n442), .A2(new_n443), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n438), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n432), .A2(G200), .ZN(new_n450));
  INV_X1    g0250(.A(G190), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n447), .C1(new_n451), .C2(new_n432), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT75), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT75), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n449), .A2(new_n455), .A3(new_n452), .ZN(new_n456));
  AOI211_X1 g0256(.A(new_n378), .B(new_n418), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT83), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT82), .ZN(new_n460));
  OAI21_X1  g0260(.A(G257), .B1(new_n317), .B2(new_n318), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G264), .A2(G1698), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n301), .ZN(new_n464));
  INV_X1    g0264(.A(G303), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n278), .B2(new_n280), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n460), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  AOI211_X1 g0268(.A(KEYINPUT82), .B(new_n466), .C1(new_n463), .C2(new_n301), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n468), .A2(new_n469), .A3(new_n325), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n203), .B(G45), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n473), .A2(new_n311), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n314), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n221), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n459), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n464), .A2(new_n467), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT82), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n464), .A2(new_n460), .A3(new_n467), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n324), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n476), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(KEYINPUT83), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT84), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n220), .A2(G20), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n204), .C1(G33), .C2(new_n226), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n269), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n484), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n488), .A2(new_n489), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n484), .A3(new_n489), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n265), .A2(new_n485), .ZN(new_n495));
  INV_X1    g0295(.A(new_n269), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n496), .B(new_n355), .C1(G1), .C2(new_n277), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n220), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n477), .A2(G169), .A3(new_n483), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n470), .A2(new_n476), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G179), .A3(new_n500), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n477), .A2(G169), .A3(new_n483), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n500), .A2(KEYINPUT21), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(KEYINPUT85), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n318), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n225), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n227), .A2(new_n321), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n301), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G294), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n325), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n475), .A2(new_n230), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n474), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT90), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n521), .B2(new_n522), .ZN(new_n527));
  INV_X1    g0327(.A(new_n522), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n319), .A2(new_n225), .B1(new_n227), .B2(new_n321), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(new_n301), .B1(G33), .B2(G294), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n528), .B(KEYINPUT90), .C1(new_n530), .C2(new_n325), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n531), .A3(new_n474), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n525), .A2(new_n342), .B1(new_n532), .B2(new_n374), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT22), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n534), .A2(new_n224), .A3(G20), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n297), .A2(new_n278), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n278), .A2(new_n280), .A3(new_n204), .A4(G87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n229), .A2(G20), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n229), .A2(KEYINPUT23), .A3(G20), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n536), .A2(new_n538), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT88), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n537), .A2(new_n534), .B1(new_n541), .B2(new_n542), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n536), .A4(new_n544), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(KEYINPUT24), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n269), .A3(new_n552), .ZN(new_n553));
  OR2_X1    g0353(.A1(new_n265), .A2(new_n539), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(KEYINPUT89), .B2(KEYINPUT25), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(KEYINPUT89), .B2(KEYINPUT25), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(KEYINPUT89), .A3(KEYINPUT25), .ZN(new_n557));
  INV_X1    g0357(.A(new_n497), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G107), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n553), .A2(new_n556), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n533), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n470), .A2(new_n459), .A3(new_n476), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT83), .B1(new_n481), .B2(new_n482), .ZN(new_n563));
  OAI21_X1  g0363(.A(G190), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n500), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n477), .A2(G200), .A3(new_n483), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n564), .A2(KEYINPUT87), .A3(new_n565), .A4(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n355), .A2(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n276), .A2(new_n282), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G107), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n229), .A2(KEYINPUT6), .A3(G97), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n226), .A2(new_n229), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n580), .B2(KEYINPUT6), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(G20), .B1(G77), .B2(new_n357), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n573), .A2(KEYINPUT78), .A3(G107), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n576), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n572), .B1(new_n584), .B2(new_n269), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n497), .A2(new_n226), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n475), .A2(new_n227), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(G244), .B1(new_n317), .B2(new_n318), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT4), .B1(new_n592), .B2(new_n301), .ZN(new_n593));
  INV_X1    g0393(.A(new_n486), .ZN(new_n594));
  OAI211_X1 g0394(.A(KEYINPUT4), .B(G244), .C1(new_n317), .C2(new_n318), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G250), .A2(G1698), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n281), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n474), .B(new_n590), .C1(new_n598), .C2(new_n325), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n342), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT80), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n599), .B2(G179), .ZN(new_n602));
  INV_X1    g0402(.A(new_n597), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n298), .A2(new_n591), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n486), .C1(new_n604), .C2(KEYINPUT4), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n589), .B1(new_n605), .B2(new_n324), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT80), .A3(new_n374), .A4(new_n474), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n588), .A2(new_n600), .A3(new_n602), .A4(new_n607), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n572), .B(new_n586), .C1(new_n584), .C2(new_n269), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n599), .A2(G200), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n599), .B2(new_n451), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n606), .A2(KEYINPUT79), .A3(G190), .A4(new_n474), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n609), .A2(new_n610), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(G238), .B1(new_n317), .B2(new_n318), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G244), .A2(G1698), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n301), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n324), .ZN(new_n622));
  INV_X1    g0422(.A(G45), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n225), .B1(new_n623), .B2(G1), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n203), .A2(new_n311), .A3(G45), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n314), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT81), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT81), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n314), .A2(new_n624), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n368), .B1(new_n622), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n621), .A2(new_n324), .B1(new_n629), .B2(new_n627), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(G190), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n301), .A2(new_n204), .A3(G68), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n277), .A2(new_n226), .A3(G20), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT19), .ZN(new_n636));
  AOI21_X1  g0436(.A(G20), .B1(new_n422), .B2(KEYINPUT19), .ZN(new_n637));
  NOR3_X1   g0437(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n634), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n269), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n360), .A2(new_n266), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n558), .A2(G87), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n640), .B(new_n641), .C1(new_n360), .C2(new_n497), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n618), .A2(new_n301), .B1(G33), .B2(G116), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n630), .B(G179), .C1(new_n645), .C2(new_n325), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n632), .B2(new_n342), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n633), .A2(new_n643), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n451), .A2(new_n525), .B1(new_n532), .B2(new_n368), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n560), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n615), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n514), .A2(new_n561), .A3(new_n571), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n458), .A2(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n398), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n344), .A2(new_n345), .ZN(new_n655));
  INV_X1    g0455(.A(new_n449), .ZN(new_n656));
  INV_X1    g0456(.A(new_n376), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n452), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n333), .A2(new_n338), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n410), .A2(new_n417), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT21), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n488), .A2(new_n484), .A3(new_n489), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n490), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n498), .B1(new_n665), .B2(new_n492), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n495), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(G169), .A3(new_n477), .A4(new_n483), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n504), .A2(new_n561), .A3(new_n668), .A4(new_n507), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT91), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n510), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(KEYINPUT91), .A3(new_n561), .A4(new_n504), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n671), .A2(new_n651), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n608), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .A3(new_n648), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(new_n648), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n608), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n676), .A2(new_n679), .B1(new_n644), .B2(new_n647), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n662), .B1(new_n458), .B2(new_n682), .ZN(G369));
  OR3_X1    g0483(.A1(new_n265), .A2(KEYINPUT27), .A3(G20), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT27), .B1(new_n265), .B2(G20), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G213), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT92), .Z(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n514), .B(new_n571), .C1(new_n565), .C2(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n500), .B(new_n689), .C1(new_n505), .C2(new_n510), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n649), .A2(new_n560), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n560), .A2(new_n689), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n561), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n533), .A2(new_n560), .A3(new_n690), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n513), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT85), .B1(new_n668), .B2(new_n507), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n504), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(new_n561), .A3(new_n690), .A4(new_n697), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n698), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n207), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n638), .A2(new_n220), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(new_n203), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g0515(.A(new_n710), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n714), .B(new_n715), .C1(new_n245), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n561), .B(new_n504), .C1(new_n702), .C2(new_n703), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n651), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT95), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(KEYINPUT95), .A3(new_n651), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n680), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n719), .B1(new_n725), .B2(new_n690), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n681), .A2(new_n690), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(KEYINPUT29), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n606), .A2(new_n474), .A3(new_n531), .A4(new_n527), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n481), .A2(new_n632), .A3(G179), .A4(new_n482), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n470), .A2(new_n476), .A3(new_n646), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n527), .A2(new_n531), .A3(new_n474), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT30), .A4(new_n606), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n477), .A2(new_n483), .ZN(new_n737));
  INV_X1    g0537(.A(new_n632), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n532), .A2(new_n374), .A3(new_n599), .A4(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n733), .B(new_n736), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT31), .B1(new_n740), .B2(new_n689), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT94), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n689), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT94), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n743), .B(new_n749), .C1(new_n652), .C2(new_n689), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n729), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n718), .B1(new_n752), .B2(G1), .ZN(G364));
  XNOR2_X1  g0553(.A(new_n694), .B(KEYINPUT97), .ZN(new_n754));
  INV_X1    g0554(.A(G13), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n203), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n710), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G330), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n691), .A2(new_n761), .A3(new_n692), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT96), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n754), .A2(new_n760), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n204), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n693), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n239), .B1(G20), .B2(new_n342), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n374), .A2(new_n368), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n204), .A2(new_n451), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n218), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n204), .B1(new_n776), .B2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n226), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n374), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n281), .B(new_n778), .C1(G58), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n368), .A2(G179), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n773), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n204), .A2(G190), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n776), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n287), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n779), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n783), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G77), .A2(new_n792), .B1(new_n794), .B2(G107), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n782), .A2(new_n786), .A3(new_n790), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n772), .A2(new_n787), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n775), .B(new_n796), .C1(G68), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n774), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT101), .B(G326), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n800), .A2(new_n801), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n777), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G294), .ZN(new_n805));
  INV_X1    g0605(.A(new_n788), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G329), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n803), .A2(new_n281), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n792), .A2(G311), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n793), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G322), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n465), .A2(new_n784), .B1(new_n780), .B2(new_n812), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n808), .A2(new_n809), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n771), .B1(new_n799), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n246), .A2(new_n623), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n709), .A2(new_n301), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(new_n258), .C2(new_n623), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n207), .A2(G355), .A3(new_n275), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G116), .C2(new_n207), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT99), .Z(new_n821));
  INV_X1    g0621(.A(new_n771), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n769), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT100), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n770), .A2(new_n815), .A3(new_n759), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n767), .A2(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n689), .A2(new_n367), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n372), .A2(new_n376), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT103), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT103), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n372), .A2(new_n832), .A3(new_n376), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n376), .B2(new_n690), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n768), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n771), .A2(new_n768), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n215), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n281), .B1(new_n793), .B2(new_n224), .C1(new_n220), .C2(new_n791), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n778), .B1(G311), .B2(new_n806), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n810), .B2(new_n797), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n840), .B(new_n842), .C1(G303), .C2(new_n800), .ZN(new_n843));
  INV_X1    g0643(.A(G294), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n229), .B2(new_n784), .C1(new_n844), .C2(new_n780), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G143), .A2(new_n781), .B1(new_n792), .B2(G159), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n774), .C1(new_n393), .C2(new_n797), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT34), .Z(new_n849));
  OAI22_X1  g0649(.A1(new_n784), .A2(new_n218), .B1(new_n793), .B2(new_n211), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT102), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n850), .A2(new_n851), .B1(G132), .B2(new_n806), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n298), .B1(G58), .B2(new_n804), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(new_n851), .C2(new_n850), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n845), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n771), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n837), .A2(new_n759), .A3(new_n839), .A4(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n689), .B(new_n834), .C1(new_n674), .C2(new_n680), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n727), .B2(new_n836), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(new_n751), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n860), .B2(new_n759), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n756), .A2(new_n203), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n741), .A2(new_n742), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n652), .B2(new_n689), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n835), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n448), .A2(new_n689), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT105), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n438), .A2(new_n867), .A3(new_n448), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n438), .B2(new_n448), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n452), .B(new_n866), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n656), .A2(new_n689), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n865), .A2(new_n872), .A3(KEYINPUT40), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n687), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n303), .A2(new_n307), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n496), .B1(new_n876), .B2(new_n273), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT106), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n303), .B2(new_n307), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT106), .B1(new_n880), .B2(new_n496), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n308), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n335), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n346), .A2(new_n875), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n687), .B(new_n341), .C1(new_n331), .C2(new_n342), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n336), .B1(new_n886), .B2(new_n309), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n339), .B1(new_n877), .B2(new_n878), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n272), .B1(new_n889), .B2(new_n881), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n336), .B1(new_n890), .B2(new_n886), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n888), .B1(new_n891), .B2(KEYINPUT37), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n874), .B1(new_n884), .B2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(new_n336), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n883), .B2(new_n885), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n346), .A2(new_n875), .A3(new_n883), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n735), .A2(G200), .B1(G190), .B2(new_n524), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n553), .A2(new_n557), .A3(new_n559), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(new_n556), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(new_n608), .A3(new_n614), .A4(new_n648), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n569), .B2(new_n570), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n906), .A2(new_n561), .A3(new_n514), .A4(new_n690), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n836), .B1(new_n907), .B2(new_n863), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n346), .A2(new_n340), .A3(new_n875), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n887), .B(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n874), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n900), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n870), .A2(new_n871), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n908), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n873), .A2(new_n901), .B1(new_n915), .B2(KEYINPUT40), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n457), .A2(new_n864), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n916), .B(new_n917), .Z(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G330), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT107), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n457), .B1(new_n726), .B2(new_n728), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n662), .ZN(new_n922));
  INV_X1    g0722(.A(new_n834), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n681), .A2(new_n690), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n376), .A2(new_n689), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n872), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n901), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n900), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT39), .B1(new_n912), .B2(new_n900), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n868), .A2(new_n869), .A3(new_n689), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n655), .A2(new_n875), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n928), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n922), .B(new_n935), .Z(new_n936));
  AOI21_X1  g0736(.A(new_n862), .B1(new_n920), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT108), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n920), .B2(new_n936), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n246), .A2(G77), .A3(new_n284), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(G50), .B2(new_n211), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n755), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n220), .B1(new_n581), .B2(KEYINPUT35), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n943), .B(new_n240), .C1(KEYINPUT35), .C2(new_n581), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT104), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT36), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n942), .A3(new_n946), .ZN(G367));
  NOR3_X1   g0747(.A1(new_n254), .A2(new_n709), .A3(new_n301), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n825), .B1(new_n207), .B2(new_n360), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n791), .A2(new_n218), .B1(new_n788), .B2(new_n847), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n797), .A2(new_n287), .B1(new_n793), .B2(new_n215), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(G58), .C2(new_n785), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n804), .A2(G68), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n781), .A2(G150), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n281), .B1(new_n800), .B2(G143), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n777), .A2(new_n229), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n785), .A2(G116), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT46), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n793), .A2(new_n226), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n301), .B(new_n960), .C1(G303), .C2(new_n781), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n800), .A2(G311), .ZN(new_n962));
  XNOR2_X1  g0762(.A(KEYINPUT113), .B(G317), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n791), .A2(new_n810), .B1(new_n788), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G294), .B2(new_n798), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n959), .A2(new_n961), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n956), .B1(new_n957), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT47), .Z(new_n968));
  OAI221_X1 g0768(.A(new_n759), .B1(new_n948), .B2(new_n949), .C1(new_n968), .C2(new_n822), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT114), .Z(new_n970));
  NOR2_X1   g0770(.A1(new_n690), .A2(new_n643), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(new_n644), .A3(new_n647), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n678), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n970), .B1(new_n769), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n975));
  OAI211_X1 g0775(.A(new_n608), .B(new_n614), .C1(new_n609), .C2(new_n690), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT109), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT109), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n675), .A2(new_n689), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n975), .B1(new_n981), .B2(new_n706), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n981), .A2(new_n706), .A3(new_n975), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n698), .A3(new_n705), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n700), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT45), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n986), .B(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n990), .A2(new_n983), .A3(new_n701), .A4(new_n984), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n699), .B1(new_n514), .B2(new_n689), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT111), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT111), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n705), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n694), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n754), .B2(new_n996), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n752), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n710), .B(KEYINPUT41), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT112), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT112), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n758), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n700), .A2(new_n980), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n977), .A2(new_n978), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n705), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT42), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n608), .B1(new_n1011), .B2(new_n561), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1014), .A2(new_n690), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1010), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1009), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n974), .B1(new_n1006), .B2(new_n1017), .ZN(G387));
  OR2_X1    g0818(.A1(new_n752), .A2(new_n998), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n752), .A2(new_n998), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n710), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n769), .B1(new_n697), .B2(new_n698), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n791), .A2(new_n211), .B1(new_n788), .B2(new_n393), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n784), .A2(new_n215), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n780), .A2(new_n218), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n960), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n360), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n804), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n798), .A2(new_n264), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n298), .B1(G159), .B2(new_n800), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G311), .A2(new_n798), .B1(new_n792), .B2(G303), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n812), .B2(new_n774), .C1(new_n780), .C2(new_n963), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT48), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n810), .B2(new_n777), .C1(new_n844), .C2(new_n784), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT49), .Z(new_n1036));
  AOI21_X1  g0836(.A(new_n301), .B1(new_n806), .B2(new_n801), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n220), .B2(new_n793), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1031), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n760), .B1(new_n1039), .B2(new_n771), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n263), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n711), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(G68), .A2(G77), .ZN(new_n1043));
  OAI21_X1  g0843(.A(KEYINPUT50), .B1(new_n263), .B2(G50), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1042), .A2(new_n623), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n817), .B(new_n1045), .C1(new_n251), .C2(new_n623), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n207), .A2(new_n275), .A3(new_n711), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(G107), .C2(new_n207), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT115), .Z(new_n1049));
  OAI21_X1  g0849(.A(new_n1040), .B1(new_n824), .B2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT116), .Z(new_n1051));
  OAI221_X1 g0851(.A(new_n1021), .B1(new_n757), .B2(new_n999), .C1(new_n1022), .C2(new_n1051), .ZN(G393));
  AOI22_X1  g0852(.A1(G317), .A2(new_n800), .B1(new_n781), .B2(G311), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT52), .Z(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n465), .B2(new_n797), .C1(new_n812), .C2(new_n788), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G116), .B2(new_n804), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n275), .B1(new_n794), .B2(G107), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n792), .A2(G294), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n785), .A2(G283), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n793), .A2(new_n224), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n798), .A2(G50), .B1(new_n804), .B2(G77), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n263), .B2(new_n791), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT117), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1061), .B(new_n1064), .C1(G68), .C2(new_n785), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n806), .A2(G143), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n774), .A2(new_n393), .B1(new_n780), .B2(new_n287), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(new_n301), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n822), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n825), .B1(new_n226), .B2(new_n207), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n261), .B2(new_n817), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1070), .A2(new_n760), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n769), .B2(new_n980), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n992), .B2(new_n757), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1020), .A2(new_n992), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n716), .B1(new_n1020), .B2(new_n992), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G390));
  OR2_X1    g0879(.A1(new_n929), .A2(new_n930), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n927), .B2(new_n932), .ZN(new_n1081));
  AND4_X1   g0881(.A1(G330), .A2(new_n750), .A3(new_n835), .A4(new_n914), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n725), .A2(new_n690), .A3(new_n923), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n872), .B1(new_n1083), .B2(new_n926), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n932), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n913), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1081), .B(new_n1082), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n914), .B1(new_n858), .B2(new_n925), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n931), .B1(new_n1088), .B2(new_n1085), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1083), .A2(new_n926), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n914), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1086), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n908), .A2(G330), .A3(new_n914), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1087), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n758), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1080), .A2(new_n768), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n838), .A2(new_n263), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n780), .A2(new_n220), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n281), .B1(new_n777), .B2(new_n215), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n786), .B1(new_n211), .B2(new_n793), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(G107), .C2(new_n798), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n810), .B2(new_n774), .C1(new_n844), .C2(new_n788), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1100), .B(new_n1104), .C1(G97), .C2(new_n792), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n275), .B1(new_n793), .B2(new_n218), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT121), .Z(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT54), .B(G143), .Z(new_n1108));
  NAND2_X1  g0908(.A1(new_n792), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G128), .A2(new_n800), .B1(new_n781), .B2(G132), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n797), .A2(new_n847), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n785), .A2(G150), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT53), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1115), .A2(new_n788), .B1(new_n777), .B2(new_n287), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n771), .B1(new_n1105), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1098), .A2(new_n759), .A3(new_n1099), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1097), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT122), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT122), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1097), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n914), .B1(new_n908), .B2(G330), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1082), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1090), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n743), .A2(new_n749), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n571), .A2(new_n651), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1129), .A2(new_n720), .A3(new_n689), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n835), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n872), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1094), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n924), .A2(new_n926), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1126), .A2(new_n1127), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT118), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n457), .A2(new_n1136), .A3(G330), .A4(new_n864), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n418), .B1(new_n454), .B2(new_n456), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n378), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1138), .A2(new_n864), .A3(G330), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT118), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n921), .A3(new_n662), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1135), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1096), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1096), .A2(new_n1144), .A3(KEYINPUT119), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n710), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1096), .A2(new_n1144), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT120), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1124), .B1(new_n1150), .B2(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(KEYINPUT57), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1157));
  OR2_X1    g0957(.A1(new_n418), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n875), .A2(new_n396), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n418), .A2(new_n1157), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1160), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n916), .B2(new_n761), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n916), .A2(new_n761), .A3(new_n1164), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n935), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n935), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n1165), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1155), .B1(new_n1156), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1143), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1096), .A2(KEYINPUT119), .A3(new_n1144), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT119), .B1(new_n1096), .B2(new_n1144), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1172), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(KEYINPUT57), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1173), .A2(new_n710), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1168), .A2(new_n1171), .A3(new_n758), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n768), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1182));
  AOI21_X1  g0982(.A(G41), .B1(new_n1027), .B2(new_n792), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n793), .A2(new_n213), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G116), .B2(new_n800), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(new_n215), .C2(new_n784), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n788), .A2(new_n810), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n953), .B1(new_n226), .B2(new_n797), .C1(new_n229), .C2(new_n780), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(new_n1186), .A2(new_n301), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT58), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G128), .A2(new_n781), .B1(new_n792), .B2(G137), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n785), .A2(new_n1108), .B1(new_n804), .B2(G150), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n800), .A2(G125), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G132), .B2(new_n798), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT59), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G33), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G41), .B1(new_n806), .B2(G124), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n287), .C2(new_n793), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G41), .B1(new_n297), .B2(G33), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1199), .A2(new_n1200), .B1(G50), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n771), .B1(new_n1190), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n838), .A2(new_n218), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1182), .A2(new_n759), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1181), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1180), .A2(new_n1207), .ZN(G375));
  INV_X1    g1008(.A(new_n1135), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n215), .A2(new_n793), .B1(new_n791), .B2(new_n229), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n275), .B1(new_n806), .B2(G303), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1028), .B(new_n1211), .C1(new_n226), .C2(new_n784), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(G283), .C2(new_n781), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n220), .B2(new_n797), .C1(new_n844), .C2(new_n774), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n791), .A2(new_n393), .ZN(new_n1215));
  INV_X1    g1015(.A(G132), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n774), .A2(new_n1216), .B1(new_n784), .B2(new_n287), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(G50), .C2(new_n804), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n806), .A2(G128), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n798), .A2(new_n1108), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n298), .B(new_n1184), .C1(G137), .C2(new_n781), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n822), .B1(new_n1214), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n760), .B(new_n1223), .C1(new_n211), .C2(new_n838), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n872), .A2(new_n768), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT123), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1209), .A2(new_n758), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1001), .B1(new_n1209), .B2(new_n1174), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n1144), .ZN(G381));
  INV_X1    g1029(.A(new_n1120), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(G375), .A2(new_n1231), .ZN(new_n1232));
  OR3_X1    g1032(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1233), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(G407));
  OAI21_X1  g1035(.A(new_n1232), .B1(new_n1234), .B2(new_n688), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(G213), .ZN(G409));
  AOI21_X1  g1037(.A(new_n1172), .B1(new_n1149), .B2(new_n1174), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1206), .B1(new_n1238), .B2(new_n1001), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT124), .B1(new_n1239), .B2(new_n1231), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1179), .A2(new_n710), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G378), .B(new_n1207), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1177), .A2(new_n1001), .A3(new_n1178), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1207), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT124), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1151), .B(KEYINPUT120), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n716), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1120), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1240), .A2(new_n1243), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n688), .A2(G213), .ZN(new_n1252));
  XOR2_X1   g1052(.A(G384), .B(KEYINPUT125), .Z(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1209), .A2(new_n1174), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n716), .B1(new_n1255), .B2(KEYINPUT60), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1144), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(KEYINPUT60), .C2(new_n1255), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1254), .B1(new_n1258), .B2(new_n1227), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1258), .A2(new_n1227), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1251), .A2(new_n1252), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT62), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n688), .A2(G213), .A3(G2897), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1260), .A2(new_n1262), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1262), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1270), .B2(new_n1259), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1266), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1251), .A2(new_n1276), .A3(new_n1252), .A4(new_n1263), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1265), .A2(new_n1274), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(G393), .B(G396), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n974), .B(G390), .C1(new_n1006), .C2(new_n1017), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1279), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(new_n1078), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1280), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1284), .A2(new_n1282), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1278), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1272), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1264), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1251), .A2(KEYINPUT63), .A3(new_n1252), .A4(new_n1263), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1292), .A2(new_n1275), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1289), .A2(new_n1295), .ZN(G405));
  INV_X1    g1096(.A(new_n1243), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1231), .B1(new_n1180), .B2(new_n1207), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT127), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1263), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT127), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1293), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1293), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1301), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1303), .A2(new_n1302), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1288), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1309), .A2(new_n1300), .A3(new_n1299), .A4(new_n1304), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(G402));
endmodule


