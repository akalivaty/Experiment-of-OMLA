//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n221, new_n222, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n231, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1197, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND3_X1  g0009(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n210));
  OAI21_X1  g0010(.A(G50), .B1(G58), .B2(G68), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT64), .Z(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n218), .C2(KEYINPUT1), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0020(.A(G226), .B(G232), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n226), .B(new_n229), .ZN(G358));
  XNOR2_X1  g0030(.A(G50), .B(G68), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G58), .B(G77), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(G107), .B(G116), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G351));
  AND2_X1   g0037(.A1(G33), .A2(G41), .ZN(new_n238));
  NAND2_X1  g0038(.A1(G1), .A2(G13), .ZN(new_n239));
  OAI21_X1  g0039(.A(KEYINPUT67), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(G33), .A2(G41), .ZN(new_n241));
  INV_X1    g0041(.A(KEYINPUT67), .ZN(new_n242));
  NAND4_X1  g0042(.A1(new_n241), .A2(new_n242), .A3(G1), .A4(G13), .ZN(new_n243));
  AND2_X1   g0043(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n245), .B1(G41), .B2(G45), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n244), .A2(G226), .A3(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n246), .ZN(new_n248));
  NAND4_X1  g0048(.A1(new_n240), .A2(new_n248), .A3(G274), .A4(new_n243), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n238), .A2(new_n239), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G222), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G223), .A3(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(new_n256), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n250), .B1(new_n251), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G190), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT9), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT8), .ZN(new_n267));
  INV_X1    g0067(.A(G58), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(KEYINPUT8), .A3(G58), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G20), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n266), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n239), .B1(new_n206), .B2(new_n252), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n275), .A2(new_n278), .B1(new_n202), .B2(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n245), .A2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n263), .B1(new_n264), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n264), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n262), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT11), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n284), .A2(new_n285), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n274), .A2(new_n260), .B1(new_n273), .B2(G68), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  INV_X1    g0102(.A(new_n265), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n202), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n265), .A2(KEYINPUT73), .A3(G50), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n299), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n282), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT12), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n304), .A2(new_n305), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n278), .B(KEYINPUT11), .C1(new_n311), .C2(new_n301), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n286), .A2(G68), .A3(new_n287), .ZN(new_n313));
  AND4_X1   g0113(.A1(new_n307), .A2(new_n310), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G226), .A2(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G232), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n256), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G97), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n251), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n240), .A2(G238), .A3(new_n246), .A4(new_n243), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n249), .A4(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n256), .A2(new_n318), .B1(G33), .B2(G97), .ZN(new_n326));
  INV_X1    g0126(.A(new_n251), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n249), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G169), .ZN(new_n331));
  AND2_X1   g0131(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n331), .A2(new_n332), .B1(new_n333), .B2(new_n330), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n331), .A2(new_n332), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n315), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n286), .A2(G77), .A3(new_n287), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G20), .A2(G77), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT15), .B(G87), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n338), .B1(new_n339), .B2(new_n274), .C1(new_n303), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n278), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n282), .A2(new_n260), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n240), .A2(G244), .A3(new_n246), .A4(new_n243), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n249), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n253), .A2(new_n255), .A3(G238), .A4(G1698), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n253), .A2(new_n255), .A3(G232), .A4(new_n257), .ZN(new_n349));
  INV_X1    g0149(.A(G107), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n348), .B(new_n349), .C1(new_n256), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n251), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT71), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT71), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n347), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n345), .B1(new_n357), .B2(new_n333), .ZN(new_n358));
  INV_X1    g0158(.A(new_n356), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n355), .B1(new_n347), .B2(new_n352), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n262), .A2(new_n333), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n291), .C1(G169), .C2(new_n262), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n298), .A2(new_n336), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n272), .B1(new_n245), .B2(G20), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n286), .A2(new_n368), .B1(new_n282), .B2(new_n272), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n268), .A2(new_n308), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n371), .B2(new_n201), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n265), .A2(G159), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT76), .B1(new_n254), .B2(G33), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT76), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n252), .A3(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n378), .A3(new_n255), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n379), .A2(new_n273), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n379), .B2(new_n273), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT16), .B(new_n375), .C1(new_n387), .C2(new_n308), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n253), .A2(new_n255), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n389), .B2(new_n273), .ZN(new_n390));
  AOI211_X1 g0190(.A(new_n385), .B(G20), .C1(new_n253), .C2(new_n255), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n375), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n300), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n370), .B1(new_n388), .B2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n240), .A2(G232), .A3(new_n246), .A4(new_n243), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT78), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n249), .B1(new_n397), .B2(KEYINPUT78), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT79), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT78), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n244), .A2(new_n402), .A3(G232), .A4(new_n246), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT79), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(new_n398), .A4(new_n249), .ZN(new_n405));
  INV_X1    g0205(.A(G223), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n257), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(G226), .B2(new_n257), .ZN(new_n408));
  INV_X1    g0208(.A(G87), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n379), .A2(new_n408), .B1(new_n252), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(G190), .B1(new_n410), .B2(new_n251), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n401), .A2(new_n405), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n251), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n403), .A2(new_n413), .A3(new_n398), .A4(new_n249), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n294), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n396), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(G179), .B1(new_n410), .B2(new_n251), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n401), .A2(new_n405), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n414), .A2(new_n362), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n379), .A2(new_n273), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n380), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n379), .A2(new_n273), .A3(new_n381), .ZN(new_n426));
  INV_X1    g0226(.A(new_n386), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n394), .B(new_n374), .C1(new_n428), .C2(G68), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n385), .B1(new_n256), .B2(G20), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n389), .A2(KEYINPUT7), .A3(new_n273), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n374), .B1(new_n432), .B2(G68), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n278), .B1(new_n433), .B2(KEYINPUT16), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n369), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n423), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n396), .A2(new_n416), .A3(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n421), .A2(new_n422), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT18), .B1(new_n396), .B2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n419), .A2(new_n437), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n354), .A2(G200), .A3(new_n356), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n345), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT72), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n357), .A2(G190), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n442), .A2(KEYINPUT72), .A3(new_n345), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT74), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n325), .A2(new_n329), .A3(G190), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n314), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n294), .B1(new_n325), .B2(new_n329), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n452), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT74), .A3(new_n314), .A4(new_n450), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g0257(.A1(new_n367), .A2(new_n441), .A3(new_n448), .A4(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n281), .A2(G107), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT25), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n245), .A2(G33), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT80), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n300), .A2(new_n281), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n463), .B2(new_n350), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n274), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n256), .A2(new_n273), .A3(G87), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT22), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n376), .A2(new_n378), .A3(new_n273), .A4(new_n255), .ZN(new_n470));
  OR3_X1    g0270(.A1(new_n470), .A2(new_n468), .A3(new_n409), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT85), .B1(new_n350), .B2(G20), .ZN(new_n472));
  XOR2_X1   g0272(.A(new_n472), .B(KEYINPUT23), .Z(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT24), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT24), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n469), .A2(new_n471), .A3(new_n476), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n464), .B1(new_n478), .B2(new_n278), .ZN(new_n479));
  INV_X1    g0279(.A(G250), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n257), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G257), .B2(new_n257), .ZN(new_n482));
  INV_X1    g0282(.A(G294), .ZN(new_n483));
  OAI22_X1  g0283(.A1(new_n379), .A2(new_n482), .B1(new_n252), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n327), .B1(new_n484), .B2(KEYINPUT86), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT86), .ZN(new_n486));
  OAI221_X1 g0286(.A(new_n486), .B1(new_n252), .B2(new_n483), .C1(new_n379), .C2(new_n482), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n240), .A2(new_n243), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n245), .B(G45), .C1(new_n489), .C2(KEYINPUT5), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n490), .A2(new_n491), .B1(KEYINPUT5), .B2(new_n489), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n485), .A2(new_n487), .B1(G264), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n244), .A2(G274), .A3(new_n492), .A4(new_n493), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G190), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(new_n496), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G200), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n479), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT87), .B1(new_n497), .B2(new_n362), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT87), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n499), .A2(new_n503), .A3(G169), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n502), .B(new_n504), .C1(new_n333), .C2(new_n499), .ZN(new_n505));
  INV_X1    g0305(.A(new_n479), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  INV_X1    g0308(.A(G97), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n273), .C1(G33), .C2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n510), .B(new_n276), .C1(new_n273), .C2(G116), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT20), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n300), .A2(G116), .A3(new_n281), .A4(new_n462), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n280), .A2(G20), .A3(new_n465), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n494), .A2(G270), .ZN(new_n517));
  OR2_X1    g0317(.A1(G257), .A2(G1698), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G264), .B2(new_n257), .ZN(new_n519));
  INV_X1    g0319(.A(G303), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n379), .A2(new_n519), .B1(new_n256), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n251), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n517), .A2(new_n496), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n516), .A2(new_n523), .A3(G169), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(KEYINPUT84), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n523), .A2(KEYINPUT21), .A3(G169), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n517), .A2(new_n496), .A3(G179), .A4(new_n522), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n516), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n516), .B1(G200), .B2(new_n523), .ZN(new_n534));
  INV_X1    g0334(.A(G190), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n523), .ZN(new_n536));
  AND4_X1   g0336(.A1(new_n526), .A2(new_n529), .A3(new_n533), .A4(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G97), .A2(G107), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n273), .A2(new_n538), .B1(new_n539), .B2(new_n409), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT83), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n274), .A2(new_n509), .ZN(new_n543));
  OAI22_X1  g0343(.A1(new_n470), .A2(new_n308), .B1(KEYINPUT19), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n278), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n282), .A2(new_n339), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n286), .A2(G87), .A3(new_n462), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G244), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G1698), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(G238), .B2(G1698), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n379), .A2(new_n551), .B1(new_n252), .B2(new_n465), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n251), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n245), .A2(G45), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(G274), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n480), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n244), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n553), .A2(new_n557), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G190), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n548), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n545), .B(new_n546), .C1(new_n339), .C2(new_n463), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n333), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n362), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n432), .A2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n350), .A2(KEYINPUT6), .A3(G97), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n509), .A2(new_n350), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n539), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n571), .B2(KEYINPUT6), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(G20), .B1(G77), .B2(new_n265), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n278), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n282), .A2(G97), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n463), .B2(G97), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n509), .B1(new_n286), .B2(new_n462), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT81), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n579), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n575), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n549), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(new_n257), .A3(new_n253), .A4(new_n255), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n253), .A2(new_n255), .A3(G250), .A4(G1698), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n585), .A2(new_n508), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n257), .A2(G244), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n583), .B1(new_n379), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n251), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n494), .A2(G257), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n496), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n362), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n591), .A2(new_n333), .A3(new_n496), .A4(new_n592), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n582), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n580), .B1(new_n579), .B2(new_n576), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n278), .B2(new_n574), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(G200), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n591), .A2(new_n496), .A3(new_n592), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G190), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n567), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n458), .A2(new_n507), .A3(new_n537), .A4(new_n604), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n594), .A2(new_n595), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n607), .A2(new_n562), .A3(new_n582), .A4(new_n566), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT26), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT88), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n599), .A2(new_n606), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT88), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n567), .A2(new_n611), .A3(new_n612), .A4(KEYINPUT26), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(new_n609), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n504), .B1(new_n333), .B2(new_n499), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n503), .B1(new_n499), .B2(G169), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n506), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n529), .A2(new_n533), .A3(new_n526), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n479), .A2(new_n498), .A3(new_n500), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n621), .A2(new_n567), .A3(new_n596), .A4(new_n603), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n615), .A2(new_n623), .A3(new_n566), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n458), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n437), .A2(new_n440), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT89), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n437), .A2(new_n440), .A3(KEYINPUT89), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n419), .A2(new_n438), .ZN(new_n631));
  INV_X1    g0431(.A(new_n336), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n451), .A2(new_n452), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n364), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n631), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n298), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(new_n366), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n625), .A2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(KEYINPUT91), .ZN(new_n640));
  INV_X1    g0440(.A(new_n537), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n280), .A2(new_n273), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n516), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT90), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n529), .A2(new_n533), .A3(new_n526), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n649), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  INV_X1    g0454(.A(new_n647), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n507), .B1(new_n479), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n505), .A2(new_n506), .A3(new_n647), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n640), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n653), .A2(new_n658), .A3(KEYINPUT91), .A4(G330), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n651), .A2(new_n655), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n507), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n647), .B(KEYINPUT92), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n505), .A2(new_n506), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n662), .A2(new_n668), .ZN(G399));
  NAND3_X1  g0469(.A1(new_n539), .A2(new_n409), .A3(new_n465), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n207), .A2(new_n489), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(G1), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n211), .B2(new_n672), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  INV_X1    g0475(.A(new_n666), .ZN(new_n676));
  INV_X1    g0476(.A(new_n566), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n620), .B2(new_n622), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n678), .B2(new_n615), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT29), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n608), .B(new_n609), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n647), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT29), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT31), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n523), .A2(new_n333), .A3(new_n558), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n497), .A2(new_n685), .A3(new_n601), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n601), .A2(new_n532), .A3(new_n495), .A4(new_n560), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT30), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n560), .A2(new_n591), .A3(new_n496), .A4(new_n592), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(new_n495), .A4(new_n532), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n686), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n647), .B1(new_n693), .B2(KEYINPUT93), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n497), .A2(new_n601), .A3(new_n685), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n689), .A2(new_n531), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n691), .B1(new_n696), .B2(new_n495), .ZN(new_n697));
  INV_X1    g0497(.A(new_n495), .ZN(new_n698));
  NOR4_X1   g0498(.A1(new_n689), .A2(new_n698), .A3(new_n531), .A4(KEYINPUT30), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n695), .B(KEYINPUT93), .C1(new_n697), .C2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n684), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n507), .A2(new_n537), .A3(new_n604), .A4(new_n666), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n695), .B1(new_n697), .B2(new_n699), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n680), .A2(new_n683), .B1(G330), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n675), .B1(new_n707), .B2(G1), .ZN(G364));
  INV_X1    g0508(.A(G330), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n650), .A2(new_n709), .A3(new_n652), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n279), .A2(G20), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n245), .B1(new_n711), .B2(G45), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n672), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n654), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n713), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n256), .A2(new_n207), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(KEYINPUT94), .B2(G355), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(KEYINPUT94), .B2(G355), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(G116), .B2(new_n207), .ZN(new_n719));
  INV_X1    g0519(.A(G45), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n233), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n379), .A2(new_n207), .ZN(new_n722));
  INV_X1    g0522(.A(new_n211), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n719), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G13), .A2(G33), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n239), .B1(G20), .B2(new_n362), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n715), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G179), .A2(G200), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(G20), .A3(new_n535), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT95), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(KEYINPUT95), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G159), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT32), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n273), .A2(G179), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n273), .B1(new_n733), .B2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n743), .A2(G87), .B1(new_n745), .B2(G97), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n273), .A2(new_n333), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n294), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n746), .B1(new_n202), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n747), .A2(new_n535), .A3(new_n294), .ZN(new_n752));
  NOR4_X1   g0552(.A1(new_n273), .A2(new_n333), .A3(new_n294), .A4(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n256), .B1(new_n260), .B2(new_n752), .C1(new_n754), .C2(new_n308), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n748), .A2(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n741), .A2(new_n535), .A3(G200), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n268), .B1(new_n758), .B2(new_n350), .ZN(new_n759));
  OR4_X1    g0559(.A1(new_n740), .A2(new_n751), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n738), .A2(KEYINPUT98), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n738), .A2(KEYINPUT98), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n758), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n764), .A2(G329), .B1(G283), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT99), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n749), .B(KEYINPUT96), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n769), .A2(G326), .B1(G294), .B2(new_n745), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT97), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT97), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n389), .B1(new_n752), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n757), .A2(new_n775), .B1(new_n742), .B2(new_n520), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n774), .B(new_n776), .C1(new_n753), .C2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n771), .A2(new_n772), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n760), .B1(new_n767), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n732), .B1(new_n780), .B2(new_n729), .ZN(new_n781));
  INV_X1    g0581(.A(new_n728), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n653), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n714), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G396));
  NAND2_X1  g0585(.A1(new_n344), .A2(new_n647), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n364), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(KEYINPUT100), .B1(new_n448), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT100), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n789), .A2(new_n790), .A3(new_n364), .A4(new_n786), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n364), .A2(new_n655), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT101), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n679), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n706), .A2(G330), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n715), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n797), .B2(new_n796), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n729), .A2(new_n726), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n713), .B1(new_n260), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n729), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n379), .B1(G58), .B2(new_n745), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n803), .B1(new_n202), .B2(new_n742), .C1(new_n308), .C2(new_n758), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n764), .B2(G132), .ZN(new_n805));
  INV_X1    g0605(.A(new_n752), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G159), .B1(new_n753), .B2(G150), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n750), .B2(new_n808), .C1(new_n809), .C2(new_n757), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n764), .A2(G311), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n483), .A2(new_n757), .B1(new_n750), .B2(new_n520), .ZN(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n389), .B1(new_n465), .B2(new_n752), .C1(new_n754), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n758), .A2(new_n409), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n742), .A2(new_n350), .B1(new_n744), .B2(new_n509), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n813), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n805), .A2(new_n811), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n801), .B1(new_n802), .B2(new_n819), .C1(new_n795), .C2(new_n727), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n799), .A2(new_n820), .ZN(G384));
  NOR2_X1   g0621(.A1(new_n711), .A2(new_n245), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n386), .B1(new_n424), .B2(new_n380), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n308), .B1(new_n823), .B2(new_n426), .ZN(new_n824));
  OAI211_X1 g0624(.A(KEYINPUT103), .B(new_n394), .C1(new_n824), .C2(new_n374), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n394), .A2(KEYINPUT103), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n375), .B(new_n826), .C1(new_n387), .C2(new_n308), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n278), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n439), .B1(new_n828), .B2(new_n369), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n645), .B1(new_n828), .B2(new_n369), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n396), .A2(new_n416), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT37), .ZN(new_n833));
  INV_X1    g0633(.A(new_n645), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n435), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n417), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n423), .A2(new_n435), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n833), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n832), .A2(new_n833), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n441), .A2(KEYINPUT104), .A3(new_n830), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT104), .B1(new_n441), .B2(new_n830), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n839), .B(KEYINPUT38), .C1(new_n840), .C2(new_n841), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n844), .A2(KEYINPUT105), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT105), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n842), .A2(new_n847), .A3(new_n843), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(KEYINPUT39), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n836), .B2(new_n627), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n837), .A2(new_n835), .A3(new_n417), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n835), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n630), .A2(new_n631), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n845), .B(new_n850), .C1(new_n856), .C2(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n632), .A2(new_n655), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n624), .A2(new_n795), .A3(new_n666), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n364), .A2(new_n647), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n334), .A2(new_n335), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n456), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n314), .A2(new_n655), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n633), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n867), .A2(new_n868), .B1(new_n336), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n846), .A2(new_n865), .A3(new_n848), .A4(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n630), .A2(new_n834), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n861), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n680), .A2(new_n458), .A3(new_n683), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n638), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n875), .B(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT93), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n704), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n880), .A2(KEYINPUT31), .A3(new_n647), .A4(new_n700), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n702), .A2(new_n703), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n870), .B1(new_n792), .B2(new_n794), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n846), .A2(new_n848), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n845), .B1(new_n856), .B2(KEYINPUT38), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n882), .A2(new_n883), .A3(KEYINPUT40), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n885), .A2(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n458), .A2(new_n882), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n709), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n822), .B1(new_n878), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n878), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g0694(.A(G77), .B1(new_n268), .B2(new_n308), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n895), .A2(new_n211), .B1(G50), .B2(new_n308), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(G1), .A3(new_n279), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT102), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n465), .B(new_n210), .C1(new_n572), .C2(KEYINPUT35), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(KEYINPUT35), .B2(new_n572), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT36), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n901), .B2(new_n900), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n894), .A2(new_n903), .ZN(G367));
  INV_X1    g0704(.A(new_n712), .ZN(new_n905));
  INV_X1    g0705(.A(new_n662), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n596), .B(new_n603), .C1(new_n599), .C2(new_n666), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n596), .B2(new_n666), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n668), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT109), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(KEYINPUT44), .C1(new_n668), .C2(new_n908), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n668), .A2(KEYINPUT45), .A3(new_n908), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT45), .B1(new_n668), .B2(new_n908), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n911), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n906), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n662), .A2(KEYINPUT110), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n917), .A2(KEYINPUT110), .B1(new_n918), .B2(new_n916), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n665), .B1(new_n658), .B2(new_n664), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(new_n654), .Z(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n707), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n707), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n924));
  XNOR2_X1  g0724(.A(new_n672), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n905), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n908), .A2(new_n664), .A3(new_n507), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(KEYINPUT42), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n596), .B1(new_n907), .B2(new_n618), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n927), .A2(KEYINPUT42), .B1(new_n666), .B2(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n548), .A2(new_n655), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n567), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n566), .B2(new_n931), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n928), .A2(new_n930), .B1(KEYINPUT43), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n934), .B(new_n935), .Z(new_n936));
  NAND2_X1  g0736(.A1(new_n906), .A2(new_n908), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n936), .B(new_n937), .Z(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n926), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT112), .ZN(new_n941));
  INV_X1    g0741(.A(new_n229), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n730), .B1(new_n207), .B2(new_n339), .C1(new_n942), .C2(new_n722), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n943), .A2(new_n715), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n769), .A2(G143), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n758), .A2(new_n260), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n742), .A2(new_n268), .B1(new_n744), .B2(new_n308), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(G150), .C2(new_n756), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n738), .A2(G137), .ZN(new_n949));
  INV_X1    g0749(.A(G159), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n256), .B1(new_n754), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G50), .B2(new_n806), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n945), .A2(new_n948), .A3(new_n949), .A4(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n756), .A2(G303), .B1(G107), .B2(new_n745), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n509), .B2(new_n758), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n769), .B2(G311), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n379), .B1(new_n814), .B2(new_n752), .C1(new_n754), .C2(new_n483), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G317), .B2(new_n738), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n742), .A2(new_n465), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n956), .B(new_n958), .C1(KEYINPUT46), .C2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n743), .A2(KEYINPUT46), .A3(G116), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT111), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n953), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT47), .Z(new_n964));
  OAI221_X1 g0764(.A(new_n944), .B1(new_n782), .B2(new_n933), .C1(new_n964), .C2(new_n802), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n940), .A2(new_n941), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n926), .B2(new_n939), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT112), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(G387));
  OAI22_X1  g0770(.A1(new_n716), .A2(new_n671), .B1(G107), .B2(new_n207), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n226), .A2(G45), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n340), .A2(G50), .ZN(new_n973));
  XNOR2_X1  g0773(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  AOI211_X1 g0775(.A(G45), .B(new_n670), .C1(G68), .C2(G77), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n722), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n971), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n715), .B1(new_n978), .B2(new_n731), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n756), .A2(G317), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n806), .A2(G303), .B1(new_n753), .B2(G311), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(new_n768), .C2(new_n775), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT48), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n743), .A2(G294), .B1(new_n745), .B2(G283), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT49), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n379), .B1(new_n758), .B2(new_n465), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n738), .B2(G326), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n743), .A2(G77), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n509), .B2(new_n758), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n379), .B(new_n995), .C1(G68), .C2(new_n806), .ZN(new_n996));
  INV_X1    g0796(.A(new_n272), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n749), .A2(G159), .B1(new_n997), .B2(new_n753), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n744), .A2(new_n339), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n756), .B2(G50), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n738), .A2(G150), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n802), .B1(new_n993), .B2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n979), .B(new_n1003), .C1(new_n659), .C2(new_n728), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n921), .B2(new_n905), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n672), .B(KEYINPUT114), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n922), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n921), .A2(new_n707), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G393));
  AOI21_X1  g0809(.A(KEYINPUT115), .B1(new_n906), .B2(new_n916), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n906), .A2(new_n916), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n906), .A2(KEYINPUT115), .A3(new_n916), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n905), .A4(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n730), .B1(new_n509), .B2(new_n207), .C1(new_n236), .C2(new_n722), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n715), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n389), .B1(new_n483), .B2(new_n752), .C1(new_n754), .C2(new_n520), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n737), .A2(new_n775), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n765), .A2(G107), .B1(new_n745), .B2(G116), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n814), .C2(new_n742), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n756), .A2(G311), .B1(new_n749), .B2(G317), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT52), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n744), .A2(new_n260), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1024), .B(new_n816), .C1(G68), .C2(new_n743), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n754), .A2(new_n202), .B1(new_n340), .B2(new_n752), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n379), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(new_n809), .C2(new_n737), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n756), .A2(G159), .B1(new_n749), .B2(G150), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1021), .A2(new_n1023), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1016), .B1(new_n1032), .B2(new_n729), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n908), .B2(new_n782), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1014), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n919), .A2(new_n922), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1006), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n922), .B1(new_n1039), .B2(new_n1010), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1035), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(G390));
  AOI21_X1  g0842(.A(new_n863), .B1(new_n679), .B2(new_n795), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n859), .B1(new_n1043), .B2(new_n870), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n849), .A2(new_n1044), .A3(new_n857), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n863), .B1(new_n682), .B2(new_n795), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n887), .B(new_n859), .C1(new_n870), .C2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n882), .A2(G330), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n883), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n706), .A2(G330), .A3(new_n795), .A4(new_n871), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1045), .A2(new_n1047), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1049), .A2(new_n458), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n876), .A2(new_n638), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n882), .A2(G330), .A3(new_n795), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(new_n870), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1053), .A2(new_n1046), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n795), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n870), .B1(new_n797), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1043), .B1(new_n1050), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1057), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1055), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n876), .A2(new_n638), .A3(new_n1056), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1050), .A2(new_n1063), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n865), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1052), .A2(new_n1071), .A3(new_n1054), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1066), .A2(new_n1072), .A3(new_n1006), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1045), .A2(new_n1047), .A3(new_n1053), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1050), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n905), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n800), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n715), .B1(new_n1078), .B2(new_n997), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n764), .A2(G125), .ZN(new_n1080));
  INV_X1    g0880(.A(G150), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n742), .A2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT54), .B(G143), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n256), .B1(new_n752), .B2(new_n1085), .C1(new_n754), .C2(new_n808), .ZN(new_n1086));
  INV_X1    g0886(.A(G132), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n757), .A2(new_n1087), .B1(new_n744), .B2(new_n950), .ZN(new_n1088));
  INV_X1    g0888(.A(G128), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n750), .A2(new_n1089), .B1(new_n758), .B2(new_n202), .ZN(new_n1090));
  OR4_X1    g0890(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n763), .A2(new_n483), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n389), .B1(new_n754), .B2(new_n350), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G97), .B2(new_n806), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n756), .A2(G116), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1024), .B1(new_n749), .B2(G283), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n743), .A2(G87), .B1(new_n765), .B2(G68), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1080), .A2(new_n1091), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1079), .B1(new_n1099), .B2(new_n729), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n858), .B2(new_n727), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT118), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1101), .B(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1073), .A2(new_n1077), .A3(new_n1103), .ZN(G378));
  NAND2_X1  g0904(.A1(new_n885), .A2(new_n886), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n709), .B1(new_n887), .B2(new_n888), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n298), .A2(new_n366), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n291), .A2(new_n834), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1107), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT123), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1105), .A2(new_n1106), .A3(new_n1114), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n859), .B1(new_n849), .B2(new_n857), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n872), .A2(new_n873), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n875), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1072), .A2(new_n1057), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT57), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1064), .A2(new_n1061), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1067), .B1(new_n1076), .B2(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1105), .A2(new_n1106), .A3(new_n1114), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1114), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n875), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1116), .A2(new_n1122), .A3(new_n1118), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(KEYINPUT57), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1006), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1127), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1114), .A2(new_n726), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n715), .B1(new_n1078), .B2(G50), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n994), .B1(new_n339), .B2(new_n752), .C1(new_n509), .C2(new_n754), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n757), .A2(new_n350), .B1(new_n758), .B2(new_n268), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n379), .A2(new_n489), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n749), .A2(G116), .B1(G68), .B2(new_n745), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(new_n763), .C2(new_n814), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT120), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G50), .B1(new_n252), .B2(new_n489), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1147), .A2(KEYINPUT58), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n749), .A2(G125), .B1(G150), .B2(new_n745), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT121), .Z(new_n1151));
  AOI22_X1  g0951(.A1(new_n806), .A2(G137), .B1(new_n753), .B2(G132), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n742), .B2(new_n1085), .C1(new_n1089), .C2(new_n757), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT122), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n738), .A2(G124), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G33), .B(G41), .C1(new_n765), .C2(G159), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1155), .A2(KEYINPUT122), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1149), .B1(KEYINPUT58), .B2(new_n1147), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1139), .B1(new_n1161), .B2(new_n729), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1138), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n1125), .B2(new_n905), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1137), .A2(new_n1165), .ZN(G375));
  NAND3_X1  g0966(.A1(new_n1069), .A2(new_n1070), .A3(new_n1067), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT124), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT124), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1128), .A2(new_n1169), .A3(new_n1067), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n1170), .A3(new_n925), .A4(new_n1065), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT125), .Z(new_n1172));
  AOI21_X1  g0972(.A(new_n713), .B1(new_n308), .B2(new_n800), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n750), .A2(new_n1087), .B1(new_n758), .B2(new_n268), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n754), .A2(new_n1085), .B1(new_n752), .B2(new_n1081), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1174), .A2(new_n1175), .A3(new_n379), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n756), .A2(G137), .B1(new_n743), .B2(G159), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n202), .C2(new_n744), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G128), .B2(new_n764), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n763), .A2(new_n520), .B1(new_n509), .B2(new_n742), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT126), .Z(new_n1181));
  OAI22_X1  g0981(.A1(new_n814), .A2(new_n757), .B1(new_n750), .B2(new_n483), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n389), .B1(new_n350), .B2(new_n752), .C1(new_n754), .C2(new_n465), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1182), .A2(new_n1183), .A3(new_n946), .A4(new_n999), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1179), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1173), .B1(new_n802), .B2(new_n1185), .C1(new_n871), .C2(new_n727), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1129), .B2(new_n905), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1172), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(G381));
  NAND2_X1  g0990(.A1(new_n1077), .A2(new_n1103), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1037), .B1(new_n1055), .B2(new_n1065), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1072), .B2(new_n1192), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n969), .A2(new_n1189), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1195), .A2(G375), .ZN(G407));
  NAND2_X1  g0996(.A1(new_n646), .A2(G213), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(G407), .B(G213), .C1(G375), .C2(new_n1199), .ZN(G409));
  XNOR2_X1  g1000(.A(G393), .B(new_n784), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n940), .A2(G390), .A3(new_n965), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n967), .A2(new_n1041), .A3(KEYINPUT127), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT127), .B1(new_n967), .B2(new_n1041), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1201), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n966), .A2(new_n968), .A3(new_n1041), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n967), .A2(new_n1041), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(new_n1201), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT63), .ZN(new_n1212));
  OAI211_X1 g1012(.A(G378), .B(new_n1165), .C1(new_n1127), .C2(new_n1136), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n875), .B1(new_n1214), .B2(new_n1117), .ZN(new_n1215));
  AND4_X1   g1015(.A1(new_n1117), .A2(new_n875), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n925), .B(new_n1126), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1133), .A2(new_n1134), .A3(new_n905), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1218), .A2(new_n1163), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1193), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1213), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1197), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1065), .A2(KEYINPUT60), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1167), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1037), .B1(new_n1226), .B2(KEYINPUT60), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1228), .A2(G384), .A3(new_n1188), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G384), .B1(new_n1228), .B2(new_n1188), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1212), .B1(new_n1223), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1198), .A2(G2897), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1228), .A2(new_n1188), .ZN(new_n1237));
  INV_X1    g1037(.A(G384), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1228), .A2(G384), .A3(new_n1188), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1234), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT61), .B1(new_n1223), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1198), .B1(new_n1213), .B2(new_n1221), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(KEYINPUT63), .A3(new_n1231), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1211), .A2(new_n1233), .A3(new_n1243), .A4(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT62), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1244), .A2(new_n1247), .A3(new_n1231), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT61), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1244), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1247), .B1(new_n1244), .B2(new_n1231), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1248), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1246), .B1(new_n1253), .B2(new_n1211), .ZN(G405));
  AOI21_X1  g1054(.A(G378), .B1(new_n1137), .B2(new_n1165), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n1232), .A3(new_n1213), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n967), .A2(new_n1041), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1203), .A3(new_n1202), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1261), .A2(new_n1201), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1213), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1231), .B1(new_n1255), .B2(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1257), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1262), .B1(new_n1257), .B2(new_n1264), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(G402));
endmodule


