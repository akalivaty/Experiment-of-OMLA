//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT96), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g003(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT86), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT15), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT86), .A3(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(KEYINPUT15), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  MUX2_X1   g014(.A(new_n214), .B(new_n213), .S(new_n215), .Z(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(new_n212), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(new_n212), .B2(new_n216), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT87), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g021(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT95), .B(G85gat), .ZN(new_n224));
  INV_X1    g023(.A(G92gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n223), .B1(new_n226), .B2(KEYINPUT7), .ZN(new_n227));
  AND3_X1   g026(.A1(KEYINPUT94), .A2(G99gat), .A3(G106gat), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT94), .B1(G99gat), .B2(G106gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(KEYINPUT7), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G99gat), .B(G106gat), .Z(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n235), .A3(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n222), .B(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n205), .B(new_n240), .C1(new_n242), .C2(new_n239), .ZN(new_n243));
  INV_X1    g042(.A(G162gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n202), .A2(new_n203), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n243), .B2(new_n246), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n204), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n246), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G162gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n204), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n247), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G134gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n250), .A2(new_n254), .A3(new_n257), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G15gat), .B(G22gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT16), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT89), .B(G1gat), .Z(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT90), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n262), .B(KEYINPUT88), .ZN(new_n270));
  INV_X1    g069(.A(G1gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n273), .A3(G8gat), .ZN(new_n274));
  INV_X1    g073(.A(G8gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n267), .B(new_n272), .C1(new_n268), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G64gat), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G71gat), .B(G78gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n277), .B1(KEYINPUT21), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(KEYINPUT21), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(G127gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n283), .B(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n287));
  XNOR2_X1  g086(.A(G155gat), .B(G183gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n286), .B(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(G211gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n290), .B(new_n293), .Z(new_n294));
  NAND3_X1  g093(.A1(new_n261), .A2(KEYINPUT97), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT97), .B1(new_n261), .B2(new_n294), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(KEYINPUT0), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(G57gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(G85gat), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT2), .ZN(new_n305));
  OR2_X1    g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G155gat), .B(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(KEYINPUT74), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n309), .B1(new_n308), .B2(new_n310), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G113gat), .B(G120gat), .ZN(new_n314));
  OAI21_X1  g113(.A(G127gat), .B1(new_n314), .B2(KEYINPUT1), .ZN(new_n315));
  INV_X1    g114(.A(G120gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G113gat), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G120gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321));
  INV_X1    g120(.A(G127gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n315), .A2(new_n323), .A3(G134gat), .ZN(new_n324));
  AOI21_X1  g123(.A(G134gat), .B1(new_n315), .B2(new_n323), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n313), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n310), .ZN(new_n327));
  INV_X1    g126(.A(new_n309), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G134gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n322), .B1(new_n320), .B2(new_n321), .ZN(new_n333));
  AOI211_X1 g132(.A(KEYINPUT1), .B(G127gat), .C1(new_n317), .C2(new_n319), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n323), .A3(G134gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n326), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT5), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n335), .A2(new_n336), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT3), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n311), .B2(new_n312), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n311), .B2(new_n312), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT76), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n348), .B1(new_n352), .B2(new_n343), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n324), .A2(new_n325), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n331), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n347), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n342), .B1(new_n339), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n348), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n354), .A2(new_n351), .A3(new_n350), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n347), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n340), .A2(KEYINPUT5), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n303), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n340), .B(new_n347), .C1(new_n353), .C2(new_n356), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n367), .B(new_n302), .C1(new_n368), .C2(new_n342), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(KEYINPUT6), .B(new_n303), .C1(new_n358), .C2(new_n364), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  INV_X1    g172(.A(G169gat), .ZN(new_n374));
  INV_X1    g173(.A(G176gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT23), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT67), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT67), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT23), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n373), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n383), .A2(KEYINPUT24), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(KEYINPUT23), .ZN(new_n385));
  NOR2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(KEYINPUT24), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n384), .B(new_n385), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT25), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n380), .B1(new_n379), .B2(KEYINPUT23), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n377), .B(KEYINPUT67), .C1(G169gat), .C2(G176gat), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n390), .A2(new_n391), .B1(G169gat), .B2(G176gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n383), .A2(KEYINPUT24), .ZN(new_n393));
  INV_X1    g192(.A(new_n387), .ZN(new_n394));
  INV_X1    g193(.A(new_n386), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n375), .A2(KEYINPUT66), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT66), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G176gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT65), .B(G169gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT23), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT25), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n392), .A2(new_n396), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G190gat), .ZN(new_n405));
  AND2_X1   g204(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT68), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT28), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT69), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT26), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT26), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n379), .A2(KEYINPUT69), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n373), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT27), .B(G183gat), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n409), .A2(KEYINPUT28), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n409), .A2(KEYINPUT28), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n416), .A2(new_n405), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n410), .A2(new_n415), .A3(new_n419), .A4(new_n383), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n389), .A2(new_n404), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT73), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT73), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n389), .A2(new_n420), .A3(new_n404), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G197gat), .B(G204gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT22), .ZN(new_n430));
  INV_X1    g229(.A(G218gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n292), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G211gat), .B(G218gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n427), .B(KEYINPUT72), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n421), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n428), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n427), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n422), .A2(new_n442), .A3(new_n425), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n421), .A2(new_n423), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n437), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n435), .B(KEYINPUT71), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G8gat), .B(G36gat), .Z(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(G64gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(new_n225), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n441), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n439), .B1(new_n426), .B2(new_n427), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n455), .A2(new_n436), .B1(new_n446), .B2(new_n448), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT37), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT38), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT82), .B(KEYINPUT37), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n449), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n452), .A4(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n372), .A2(KEYINPUT83), .A3(new_n454), .A4(new_n461), .ZN(new_n462));
  AOI211_X1 g261(.A(new_n435), .B(new_n439), .C1(new_n426), .C2(new_n427), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n447), .B1(new_n443), .B2(new_n445), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n460), .A2(new_n452), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT38), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n461), .A2(new_n370), .A3(new_n371), .A4(new_n454), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n462), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT80), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n345), .B1(new_n435), .B2(KEYINPUT29), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n313), .ZN(new_n476));
  NAND2_X1  g275(.A1(G228gat), .A2(G233gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT29), .B1(new_n331), .B2(new_n345), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n476), .B(new_n478), .C1(new_n447), .C2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  OR3_X1    g280(.A1(new_n479), .A2(KEYINPUT79), .A3(new_n436), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n475), .A2(new_n352), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n475), .A2(new_n352), .A3(KEYINPUT78), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT79), .B1(new_n479), .B2(new_n436), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n482), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n477), .B(KEYINPUT77), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G22gat), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n474), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(G78gat), .B(G106gat), .Z(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G50gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n490), .A2(new_n491), .ZN(new_n497));
  AOI211_X1 g296(.A(G22gat), .B(new_n481), .C1(new_n488), .C2(new_n489), .ZN(new_n498));
  OAI22_X1  g297(.A1(new_n492), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n490), .A2(new_n491), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n490), .A2(new_n491), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n500), .A2(new_n474), .A3(new_n501), .A4(new_n495), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n452), .B1(new_n463), .B2(new_n464), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(KEYINPUT30), .A3(new_n454), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n465), .A2(new_n506), .A3(new_n453), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n505), .A2(KEYINPUT81), .A3(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR3_X1    g311(.A1(new_n362), .A2(KEYINPUT39), .A3(new_n339), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n326), .A2(new_n337), .A3(new_n339), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT39), .B(new_n514), .C1(new_n362), .C2(new_n339), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n302), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT40), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n518), .A2(new_n365), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n503), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n473), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT84), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n421), .B(new_n343), .ZN(new_n524));
  NAND2_X1  g323(.A1(G227gat), .A2(G233gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT64), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT32), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT33), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G43gat), .ZN(new_n531));
  INV_X1    g330(.A(G71gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G99gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n528), .B1(new_n530), .B2(new_n534), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n524), .A2(new_n526), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n530), .A2(new_n534), .ZN(new_n543));
  INV_X1    g342(.A(new_n528), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n542), .B1(new_n545), .B2(new_n535), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n538), .A2(new_n539), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n541), .A2(new_n546), .B1(KEYINPUT34), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n540), .B1(new_n536), .B2(new_n537), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n547), .A2(KEYINPUT34), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n542), .A3(new_n535), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n548), .A2(KEYINPUT36), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT36), .B1(new_n548), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n370), .A2(new_n371), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n499), .A2(new_n502), .B1(new_n555), .B2(new_n508), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT84), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n473), .A2(new_n521), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n523), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n548), .A2(new_n552), .ZN(new_n561));
  INV_X1    g360(.A(new_n503), .ZN(new_n562));
  AND4_X1   g361(.A1(new_n555), .A2(new_n561), .A3(new_n508), .A4(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT35), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n561), .A2(new_n564), .A3(new_n562), .A4(new_n555), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n563), .A2(new_n564), .B1(new_n565), .B2(new_n512), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n277), .A2(new_n222), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n222), .B(KEYINPUT17), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n274), .A2(new_n276), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(KEYINPUT18), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n573), .B(KEYINPUT13), .Z(new_n576));
  NOR2_X1   g375(.A1(new_n277), .A2(new_n222), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n578), .A2(KEYINPUT91), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(new_n571), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n580), .A2(KEYINPUT18), .A3(new_n573), .A4(new_n568), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(KEYINPUT91), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT11), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(new_n374), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT12), .Z(new_n588));
  NOR3_X1   g387(.A1(new_n575), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(KEYINPUT92), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n574), .A2(KEYINPUT18), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT92), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n579), .A2(new_n581), .A3(new_n592), .A4(new_n582), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n588), .B(KEYINPUT85), .Z(new_n595));
  AOI21_X1  g394(.A(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n232), .A2(new_n233), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n282), .B1(new_n597), .B2(KEYINPUT98), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(new_n239), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n239), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT10), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n239), .A2(KEYINPUT10), .A3(new_n282), .ZN(new_n602));
  INV_X1    g401(.A(G230gat), .ZN(new_n603));
  INV_X1    g402(.A(G233gat), .ZN(new_n604));
  OAI22_X1  g403(.A1(new_n601), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(new_n606), .A3(new_n600), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT99), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n375), .ZN(new_n611));
  INV_X1    g410(.A(G204gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n605), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n596), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n298), .A2(new_n567), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n555), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n271), .ZN(G1324gat));
  INV_X1    g420(.A(new_n619), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n512), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n623), .A2(KEYINPUT100), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(KEYINPUT100), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(G8gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT16), .B(G8gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT101), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n626), .ZN(new_n630));
  OR3_X1    g429(.A1(new_n623), .A2(new_n626), .A3(new_n629), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n631), .A2(KEYINPUT102), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(KEYINPUT102), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n627), .B(new_n630), .C1(new_n632), .C2(new_n633), .ZN(G1325gat));
  INV_X1    g433(.A(new_n561), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n553), .A2(new_n554), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(G15gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT103), .ZN(new_n640));
  OAI22_X1  g439(.A1(new_n636), .A2(G15gat), .B1(new_n619), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT104), .Z(G1326gat));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643));
  OR3_X1    g442(.A1(new_n619), .A2(KEYINPUT105), .A3(new_n562), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT105), .B1(new_n619), .B2(new_n562), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(new_n643), .A3(new_n645), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G22gat), .ZN(G1327gat));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n652));
  INV_X1    g451(.A(new_n260), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n257), .B1(new_n250), .B2(new_n254), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n259), .A2(KEYINPUT107), .A3(new_n260), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n567), .A2(new_n651), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n261), .B1(new_n560), .B2(new_n566), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n651), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662));
  INV_X1    g461(.A(new_n294), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n618), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT106), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n662), .B1(new_n661), .B2(new_n665), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G29gat), .B1(new_n669), .B2(new_n555), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n660), .A2(new_n618), .A3(new_n663), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n671), .A2(G29gat), .A3(new_n555), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT45), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(G1328gat));
  INV_X1    g473(.A(new_n512), .ZN(new_n675));
  OAI21_X1  g474(.A(G36gat), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n671), .A2(G36gat), .A3(new_n675), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT46), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(G1329gat));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n665), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n681), .B2(new_n637), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n661), .A2(KEYINPUT109), .A3(new_n638), .A4(new_n665), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(G43gat), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n671), .A2(G43gat), .A3(new_n635), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(KEYINPUT47), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n638), .B1(new_n667), .B2(new_n668), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n688), .B2(G43gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g489(.A(KEYINPUT48), .ZN(new_n691));
  OAI21_X1  g490(.A(G50gat), .B1(new_n681), .B2(new_n562), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n671), .A2(G50gat), .A3(new_n562), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n691), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n691), .B(G50gat), .C1(new_n669), .C2(new_n562), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n693), .B1(new_n694), .B2(KEYINPUT48), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(G1331gat));
  NAND2_X1  g498(.A1(new_n594), .A2(new_n595), .ZN(new_n700));
  INV_X1    g499(.A(new_n589), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n296), .A2(new_n702), .A3(new_n297), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n617), .A3(new_n567), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT113), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n555), .B(KEYINPUT111), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT113), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT112), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g515(.A1(new_n704), .A2(KEYINPUT114), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n704), .A2(KEYINPUT114), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n675), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT115), .Z(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n722), .B(new_n723), .Z(G1333gat));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n719), .A2(new_n638), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G71gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n705), .A2(new_n532), .A3(new_n561), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n637), .B1(new_n717), .B2(new_n718), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n725), .B(new_n728), .C1(new_n730), .C2(new_n532), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n729), .A2(new_n732), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n719), .A2(new_n503), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  INV_X1    g534(.A(new_n261), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n702), .A2(new_n294), .ZN(new_n737));
  AND4_X1   g536(.A1(KEYINPUT51), .A2(new_n567), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT51), .B1(new_n660), .B2(new_n737), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n740), .A2(new_n372), .A3(new_n224), .A4(new_n617), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n651), .B1(new_n567), .B2(new_n736), .ZN(new_n742));
  AOI211_X1 g541(.A(KEYINPUT44), .B(new_n657), .C1(new_n560), .C2(new_n566), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n617), .B(new_n737), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n555), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n224), .B2(new_n745), .ZN(G1336gat));
  NOR2_X1   g545(.A1(new_n744), .A2(new_n675), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT117), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n744), .B2(new_n675), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(G92gat), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n740), .A2(new_n225), .A3(new_n617), .A4(new_n512), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n747), .B2(new_n225), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT52), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1337gat));
  XOR2_X1   g556(.A(KEYINPUT118), .B(G99gat), .Z(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n744), .B2(new_n637), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n617), .A3(new_n561), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n758), .ZN(G1338gat));
  NAND4_X1  g560(.A1(new_n661), .A2(new_n617), .A3(new_n503), .A4(new_n737), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT121), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(new_n765), .A3(G106gat), .ZN(new_n766));
  INV_X1    g565(.A(new_n617), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n562), .A2(new_n767), .A3(G106gat), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT53), .B1(new_n740), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G106gat), .B1(new_n744), .B2(new_n562), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n738), .B2(new_n739), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT119), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(new_n768), .C1(new_n738), .C2(new_n739), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n771), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n776), .A2(KEYINPUT120), .A3(KEYINPUT53), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT120), .B1(new_n776), .B2(KEYINPUT53), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n770), .B1(new_n777), .B2(new_n778), .ZN(G1339gat));
  NOR2_X1   g578(.A1(new_n572), .A2(new_n573), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n569), .A2(new_n577), .A3(new_n576), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n587), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n701), .A2(new_n617), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n605), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n615), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n601), .A2(new_n602), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n606), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(KEYINPUT54), .A3(new_n605), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(KEYINPUT55), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n616), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n786), .A2(new_n789), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n783), .B1(new_n795), .B2(new_n596), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n657), .A2(new_n796), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n701), .A2(new_n791), .A3(new_n794), .A4(new_n782), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n656), .A3(new_n655), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n294), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n298), .A2(new_n596), .A3(new_n767), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n512), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n635), .A2(new_n503), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n709), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n318), .A3(new_n702), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n805), .A2(new_n555), .A3(new_n596), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n318), .ZN(G1340gat));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n316), .A3(new_n617), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n805), .A2(new_n555), .A3(new_n767), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(new_n316), .ZN(G1341gat));
  AOI21_X1  g611(.A(G127gat), .B1(new_n806), .B2(new_n294), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n805), .A2(new_n555), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n663), .A2(new_n322), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(G1342gat));
  NAND3_X1  g615(.A1(new_n806), .A2(new_n332), .A3(new_n736), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n806), .A2(new_n819), .A3(new_n332), .A4(new_n736), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n555), .A3(new_n261), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n818), .B(new_n820), .C1(new_n332), .C2(new_n821), .ZN(G1343gat));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n296), .A2(new_n297), .A3(new_n702), .A4(new_n617), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n823), .B(new_n503), .C1(new_n824), .C2(new_n800), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n638), .A2(new_n555), .A3(new_n512), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n794), .A2(KEYINPUT122), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n794), .A2(KEYINPUT122), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n702), .B(new_n791), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n736), .B1(new_n829), .B2(new_n783), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n798), .A2(new_n656), .A3(new_n655), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n663), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n562), .B1(new_n832), .B2(new_n802), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n825), .B(new_n826), .C1(new_n833), .C2(new_n823), .ZN(new_n834));
  OAI21_X1  g633(.A(G141gat), .B1(new_n834), .B2(new_n596), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n803), .A2(new_n707), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n638), .A2(new_n562), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n596), .A2(G141gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT58), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n835), .A2(new_n842), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1344gat));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(G148gat), .C1(new_n834), .C2(new_n767), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n830), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n798), .A2(new_n736), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n294), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n823), .B(new_n503), .C1(new_n850), .C2(new_n824), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n503), .B1(new_n824), .B2(new_n800), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT57), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n851), .A2(new_n853), .A3(new_n617), .A4(new_n826), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n845), .B1(new_n854), .B2(G148gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n803), .A2(new_n707), .A3(new_n837), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n767), .A2(G148gat), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n847), .A2(new_n855), .B1(new_n856), .B2(new_n857), .ZN(G1345gat));
  OAI21_X1  g657(.A(G155gat), .B1(new_n834), .B2(new_n663), .ZN(new_n859));
  INV_X1    g658(.A(G155gat), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n836), .A2(new_n860), .A3(new_n294), .A4(new_n837), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n859), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n834), .B2(new_n657), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n856), .A2(new_n261), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n867), .A2(KEYINPUT124), .A3(new_n244), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT124), .B1(new_n867), .B2(new_n244), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(G1347gat));
  NAND2_X1  g669(.A1(new_n801), .A2(new_n802), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n804), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n675), .A2(new_n372), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n702), .A3(new_n401), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n707), .A2(new_n675), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n871), .A2(new_n804), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n596), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n875), .A2(new_n878), .ZN(G1348gat));
  NOR3_X1   g678(.A1(new_n877), .A2(new_n767), .A3(new_n400), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n874), .A2(new_n617), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n375), .ZN(G1349gat));
  NAND4_X1  g681(.A1(new_n872), .A2(new_n294), .A3(new_n416), .A4(new_n873), .ZN(new_n883));
  OAI21_X1  g682(.A(G183gat), .B1(new_n877), .B2(new_n663), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g685(.A1(new_n872), .A2(new_n736), .A3(new_n876), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G190gat), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(KEYINPUT125), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n405), .A3(new_n658), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n889), .A2(KEYINPUT125), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n889), .A2(KEYINPUT125), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n887), .A2(G190gat), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(G1351gat));
  AND2_X1   g694(.A1(new_n851), .A2(new_n853), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n637), .A2(new_n876), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n702), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(KEYINPUT126), .B(G197gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n871), .A2(new_n837), .A3(new_n873), .ZN(new_n902));
  INV_X1    g701(.A(new_n900), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n702), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1352gat));
  NAND3_X1  g704(.A1(new_n902), .A2(new_n612), .A3(new_n617), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT62), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(KEYINPUT62), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n896), .A2(new_n617), .A3(new_n898), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n907), .B(new_n908), .C1(new_n909), .C2(new_n612), .ZN(G1353gat));
  NAND3_X1  g709(.A1(new_n902), .A2(new_n292), .A3(new_n294), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n851), .A2(new_n853), .A3(new_n294), .A4(new_n898), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT63), .B1(new_n912), .B2(G211gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1354gat));
  AOI21_X1  g714(.A(G218gat), .B1(new_n902), .B2(new_n658), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n896), .A2(new_n898), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n736), .A2(G218gat), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT127), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(G1355gat));
endmodule


