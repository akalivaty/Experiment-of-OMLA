//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n635, new_n638, new_n640,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n461), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n464), .A2(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  OR2_X1    g055(.A1(new_n469), .A2(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n469), .A2(KEYINPUT66), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n477), .B(new_n480), .C1(new_n483), .C2(G136), .ZN(G162));
  NAND2_X1  g059(.A1(new_n469), .A2(G138), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT4), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n475), .B2(G126), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  AND2_X1   g067(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n494));
  OAI21_X1  g069(.A(G651), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(KEYINPUT6), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n495), .A2(G50), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(G62), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n495), .A2(new_n507), .A3(G50), .A4(new_n498), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(new_n496), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n495), .A2(new_n512), .A3(G88), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n500), .A2(new_n506), .A3(new_n508), .A4(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  AND2_X1   g091(.A1(new_n495), .A2(new_n498), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G51), .ZN(new_n518));
  OR2_X1    g093(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n497), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n513), .B1(new_n501), .B2(new_n502), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n512), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n518), .A2(new_n524), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  XOR2_X1   g106(.A(KEYINPUT70), .B(G52), .Z(new_n532));
  NAND2_X1  g107(.A1(new_n517), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT71), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n540));
  OR3_X1    g115(.A1(new_n539), .A2(new_n540), .A3(new_n497), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n539), .B2(new_n497), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n537), .A2(new_n538), .A3(new_n541), .A4(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  OAI21_X1  g120(.A(G56), .B1(new_n501), .B2(new_n502), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n545), .B1(new_n548), .B2(G651), .ZN(new_n549));
  AOI211_X1 g124(.A(KEYINPUT72), .B(new_n497), .C1(new_n546), .C2(new_n547), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n517), .A2(G43), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT73), .B(G81), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n523), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n495), .A2(G53), .A3(new_n498), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n495), .A2(new_n564), .A3(G53), .A4(new_n498), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT75), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G65), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n572), .B1(new_n501), .B2(new_n502), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n510), .A2(KEYINPUT74), .A3(new_n511), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(G78), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n523), .A2(G91), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n566), .A2(new_n577), .A3(new_n578), .ZN(G299));
  NAND4_X1  g154(.A1(new_n495), .A2(new_n512), .A3(G87), .A4(new_n513), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n495), .A2(G49), .A3(new_n498), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n510), .B2(new_n511), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n588), .A2(G73), .A3(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n495), .A2(G48), .A3(new_n498), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n495), .A2(new_n512), .A3(G86), .A4(new_n513), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G305));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n510), .B2(new_n511), .ZN(new_n596));
  AND2_X1   g171(.A1(G72), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n495), .A2(new_n512), .A3(G85), .A4(new_n513), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n495), .A2(G47), .A3(new_n498), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT77), .A4(new_n600), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n495), .A2(new_n512), .A3(G92), .A4(new_n513), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n573), .B2(new_n574), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n495), .A2(G54), .A3(new_n498), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(KEYINPUT78), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(KEYINPUT78), .B1(new_n614), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(KEYINPUT79), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n622));
  NOR3_X1   g197(.A1(new_n501), .A2(new_n502), .A3(new_n572), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT74), .B1(new_n510), .B2(new_n511), .ZN(new_n624));
  OAI21_X1  g199(.A(G66), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n497), .B1(new_n625), .B2(new_n612), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n622), .B1(new_n626), .B2(new_n615), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n608), .B1(new_n627), .B2(new_n617), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n606), .B1(new_n631), .B2(G868), .ZN(G284));
  OAI21_X1  g207(.A(new_n606), .B1(new_n631), .B2(G868), .ZN(G321));
  NAND2_X1  g208(.A1(G286), .A2(G868), .ZN(new_n634));
  INV_X1    g209(.A(G299), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G868), .ZN(G297));
  OAI21_X1  g211(.A(new_n634), .B1(new_n635), .B2(G868), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n631), .B1(new_n638), .B2(G860), .ZN(G148));
  NOR3_X1   g214(.A1(new_n551), .A2(new_n555), .A3(G868), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n631), .A2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT80), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n640), .B1(new_n642), .B2(G868), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g219(.A1(new_n475), .A2(G123), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n461), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n481), .A2(new_n482), .ZN(new_n648));
  INV_X1    g223(.A(G135), .ZN(new_n649));
  OAI221_X1 g224(.A(new_n645), .B1(new_n646), .B2(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n650), .A2(G2096), .ZN(new_n651));
  INV_X1    g226(.A(G2100), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n465), .A2(new_n471), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT12), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT13), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(G2096), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n656), .B(new_n657), .C1(new_n652), .C2(new_n655), .ZN(G156));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2451), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT16), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n664), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  AND3_X1   g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(G401));
  INV_X1    g248(.A(KEYINPUT18), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT17), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n652), .ZN(new_n681));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n677), .B2(KEYINPUT18), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(G2096), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n691), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n702));
  NOR2_X1   g277(.A1(G16), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n704));
  NAND2_X1  g279(.A1(G288), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n580), .A2(new_n582), .A3(new_n581), .A4(KEYINPUT85), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n703), .B1(new_n708), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G166), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G1971), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G6), .A2(G16), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT32), .B(G1981), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n719), .B(new_n720), .Z(new_n721));
  AND3_X1   g296(.A1(new_n711), .A2(new_n716), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G25), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G107), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n475), .B2(G119), .ZN(new_n731));
  INV_X1    g306(.A(G131), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n648), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT81), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(new_n726), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT82), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n702), .B(new_n724), .C1(new_n725), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(new_n725), .ZN(new_n741));
  MUX2_X1   g316(.A(G24), .B(G290), .S(G16), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1986), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT84), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n741), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n722), .A2(new_n723), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n740), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n740), .A2(new_n747), .A3(KEYINPUT36), .A4(new_n748), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n631), .B2(G16), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n726), .A2(G33), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n758));
  NAND3_X1  g333(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n760), .B1(new_n461), .B2(new_n761), .C1(new_n648), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT89), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n757), .B1(new_n765), .B2(new_n726), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G2072), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n712), .A2(G5), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G171), .B2(new_n712), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G1961), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G19), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n556), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1341), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n767), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(G162), .A2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G29), .B2(G35), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2090), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n726), .A2(G27), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n726), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(G2078), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(G2078), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT24), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G34), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G160), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G29), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G28), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT30), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n794), .B2(KEYINPUT30), .ZN(new_n796));
  OR2_X1    g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  NAND2_X1  g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n793), .B(new_n799), .C1(new_n776), .C2(new_n778), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n650), .A2(new_n801), .A3(new_n726), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n650), .B2(new_n726), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n792), .B2(new_n791), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n784), .A2(new_n800), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n766), .A2(G2072), .B1(G1961), .B2(new_n769), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n774), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n726), .A2(G32), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n483), .A2(G141), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT90), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT92), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT91), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT26), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n475), .A2(G129), .B1(G105), .B2(new_n471), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n811), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n808), .B1(new_n817), .B2(G29), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT27), .B(G1996), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT93), .Z(new_n821));
  OR2_X1    g396(.A1(new_n818), .A2(new_n819), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n726), .A2(G26), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT28), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n483), .A2(G140), .ZN(new_n825));
  OR2_X1    g400(.A1(G104), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT87), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G128), .B2(new_n475), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n824), .B1(new_n830), .B2(G29), .ZN(new_n831));
  INV_X1    g406(.A(G2067), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(G168), .A2(G16), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n834), .B(KEYINPUT94), .C1(G16), .C2(G21), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(KEYINPUT94), .B2(new_n834), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(G1966), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n712), .A2(G20), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT23), .Z(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G299), .B2(G16), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1956), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n836), .A2(G1966), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n822), .A2(new_n837), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n807), .A2(new_n821), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n751), .A2(new_n752), .A3(new_n756), .A4(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(G311));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(G150));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n510), .B2(new_n511), .ZN(new_n850));
  AND2_X1   g425(.A1(G80), .A2(G543), .ZN(new_n851));
  OAI21_X1  g426(.A(G651), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n495), .A2(new_n512), .A3(G93), .A4(new_n513), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n495), .A2(G55), .A3(new_n498), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT99), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n621), .A2(new_n630), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n638), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT98), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT38), .Z(new_n862));
  NOR3_X1   g437(.A1(new_n551), .A2(new_n555), .A3(new_n855), .ZN(new_n863));
  INV_X1    g438(.A(new_n855), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n548), .A2(G651), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT72), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n548), .A2(new_n545), .A3(G651), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI22_X1  g443(.A1(G43), .A2(new_n517), .B1(new_n523), .B2(new_n553), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n862), .B(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  INV_X1    g448(.A(G860), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n872), .B2(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n858), .B1(new_n873), .B2(new_n875), .ZN(G145));
  XNOR2_X1  g451(.A(new_n650), .B(G160), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n490), .A2(KEYINPUT100), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n490), .A2(KEYINPUT100), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n486), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n817), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n817), .A2(new_n882), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n830), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n764), .A2(KEYINPUT101), .ZN(new_n887));
  INV_X1    g462(.A(new_n830), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n888), .A3(new_n884), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n764), .A2(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n475), .A2(G130), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n461), .A2(G118), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n483), .B2(G142), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(new_n654), .Z(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n735), .ZN(new_n899));
  INV_X1    g474(.A(new_n891), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n886), .A2(new_n900), .A3(new_n887), .A4(new_n889), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n892), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n892), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n879), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n899), .ZN(new_n905));
  AOI211_X1 g480(.A(KEYINPUT101), .B(new_n764), .C1(new_n886), .C2(new_n889), .ZN(new_n906));
  INV_X1    g481(.A(new_n901), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n892), .A2(new_n899), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n878), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n904), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g488(.A(new_n642), .B(new_n871), .ZN(new_n914));
  AOI211_X1 g489(.A(new_n608), .B(G299), .C1(new_n627), .C2(new_n617), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n627), .A2(new_n617), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n635), .B1(new_n916), .B2(new_n609), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT41), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n620), .A2(G299), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n628), .A2(new_n635), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n915), .A2(new_n917), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(KEYINPUT102), .A3(new_n922), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n914), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n914), .B1(new_n917), .B2(new_n915), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  NAND2_X1  g505(.A1(G290), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n603), .A2(KEYINPUT103), .A3(new_n604), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G303), .A2(new_n718), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n523), .A2(G88), .B1(new_n505), .B2(G651), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n935), .A2(G305), .A3(new_n508), .A4(new_n500), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n707), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n707), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n708), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n707), .A2(new_n934), .A3(new_n936), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n931), .A3(new_n932), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n944), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n933), .A2(new_n937), .A3(new_n938), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n941), .A2(new_n942), .B1(new_n931), .B2(new_n932), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n939), .A2(new_n943), .A3(KEYINPUT104), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n949), .B(new_n950), .C1(new_n951), .C2(new_n944), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n945), .B1(new_n952), .B2(KEYINPUT42), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n928), .A2(new_n929), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n928), .B2(new_n929), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G868), .B2(new_n864), .ZN(G295));
  OAI21_X1  g532(.A(new_n956), .B1(G868), .B2(new_n864), .ZN(G331));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n855), .B1(new_n551), .B2(new_n555), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n868), .A2(new_n864), .A3(new_n869), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n961), .A2(new_n962), .A3(G286), .ZN(new_n963));
  AOI21_X1  g538(.A(G286), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g539(.A(G301), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(G168), .B1(new_n863), .B2(new_n870), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(new_n962), .A3(G286), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(G171), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n949), .A2(new_n950), .B1(new_n969), .B2(new_n925), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n963), .A2(new_n964), .A3(G301), .ZN(new_n971));
  AOI21_X1  g546(.A(G171), .B1(new_n966), .B2(new_n967), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n924), .A2(new_n926), .A3(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n970), .A2(new_n974), .A3(KEYINPUT107), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT107), .B1(new_n970), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n969), .A2(new_n925), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n939), .A2(new_n943), .A3(KEYINPUT104), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT104), .B1(new_n939), .B2(new_n943), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n949), .A2(KEYINPUT106), .A3(new_n950), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n911), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n960), .B1(new_n977), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n970), .A2(new_n974), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n970), .A2(new_n974), .A3(KEYINPUT107), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n981), .A2(new_n982), .A3(new_n980), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT106), .B1(new_n949), .B2(new_n950), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n918), .A2(new_n923), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n978), .B1(new_n996), .B2(new_n969), .ZN(new_n997));
  AOI21_X1  g572(.A(G37), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(new_n998), .A3(KEYINPUT43), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n959), .B1(new_n987), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT43), .B1(new_n977), .B2(new_n986), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n974), .A2(new_n978), .ZN(new_n1003));
  AOI21_X1  g578(.A(G37), .B1(new_n995), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n960), .B1(new_n992), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n992), .A2(new_n998), .A3(new_n960), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI211_X1 g584(.A(KEYINPUT109), .B(new_n1000), .C1(new_n1009), .C2(new_n959), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1012));
  AOI211_X1 g587(.A(KEYINPUT108), .B(new_n960), .C1(new_n992), .C2(new_n1004), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n959), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1000), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1010), .A2(new_n1016), .ZN(G397));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n882), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G160), .A2(G40), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n817), .A2(new_n1023), .A3(G1996), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT111), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n830), .B(G2067), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1996), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g604(.A(new_n1029), .B(KEYINPUT110), .Z(new_n1030));
  OAI211_X1 g605(.A(new_n1025), .B(new_n1027), .C1(new_n1030), .C2(new_n817), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n734), .B(new_n738), .Z(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1023), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G290), .B(G1986), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1023), .A2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n491), .A2(new_n1018), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1022), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n882), .A2(new_n1041), .A3(new_n1018), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1019), .A2(G2067), .A3(new_n1022), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1043), .A2(new_n755), .B1(new_n1044), .B2(KEYINPUT116), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1044), .A2(KEYINPUT116), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n859), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1956), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n882), .A2(new_n1018), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(new_n1041), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1040), .B1(new_n1038), .B2(KEYINPUT50), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n1018), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1053), .A2(new_n1040), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1038), .A2(new_n1020), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT56), .B(G2072), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(G299), .B(KEYINPUT57), .Z(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1060));
  XOR2_X1   g635(.A(new_n1058), .B(KEYINPUT117), .Z(new_n1061));
  AOI22_X1  g636(.A1(new_n1047), .A2(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1054), .A2(new_n1028), .A3(new_n1055), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1049), .A2(new_n1040), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT58), .B(G1341), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1064), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(new_n1064), .A3(new_n1068), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1063), .B1(new_n1072), .B2(new_n556), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1071), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n556), .B(new_n1063), .C1(new_n1074), .C2(new_n1069), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT61), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1059), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1079), .B2(new_n1059), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1059), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1058), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1045), .A2(new_n859), .A3(new_n1046), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT60), .B1(new_n1085), .B2(new_n1047), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n859), .A2(KEYINPUT60), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1045), .A2(new_n1087), .A3(new_n1046), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1081), .A2(new_n1084), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1062), .B1(new_n1077), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT125), .B(G1961), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1043), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1040), .B1(new_n1038), .B2(new_n1020), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT45), .B1(new_n882), .B2(new_n1018), .ZN(new_n1095));
  OR4_X1    g670(.A1(new_n1093), .A2(new_n1094), .A3(G2078), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G2078), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1054), .A2(new_n1097), .A3(new_n1055), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1098), .A2(KEYINPUT126), .A3(new_n1093), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT126), .B1(new_n1098), .B2(new_n1093), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1092), .B(new_n1096), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1054), .A2(KEYINPUT53), .A3(new_n1097), .A4(new_n1021), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1092), .B(new_n1102), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1103), .A2(new_n1104), .A3(G171), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1103), .B2(G171), .ZN(new_n1106));
  OAI221_X1 g681(.A(KEYINPUT54), .B1(G171), .B2(new_n1101), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1101), .A2(G171), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(G171), .B2(new_n1103), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G8), .ZN(new_n1112));
  INV_X1    g687(.A(G1966), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1039), .A2(new_n792), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT112), .B(G8), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(G286), .A2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT121), .Z(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT122), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT51), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1122), .A2(KEYINPUT123), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1118), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1120), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(KEYINPUT51), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1122), .A2(KEYINPUT123), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1123), .A2(new_n1128), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n708), .A2(G1976), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1066), .A2(new_n1118), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT52), .ZN(new_n1132));
  INV_X1    g707(.A(G1976), .ZN(new_n1133));
  AND2_X1   g708(.A1(G288), .A2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1134), .A2(KEYINPUT52), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1066), .A2(new_n1118), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n718), .B(G1981), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT49), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(KEYINPUT113), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(KEYINPUT113), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1136), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(G303), .A2(G8), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT55), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1050), .A2(G2090), .A3(new_n1051), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n715), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1145), .B1(new_n1148), .B2(new_n1117), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n715), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1043), .ZN(new_n1151));
  INV_X1    g726(.A(G2090), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1112), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1145), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1143), .A2(new_n1149), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1129), .A2(new_n1157), .ZN(new_n1158));
  AND4_X1   g733(.A1(new_n1090), .A2(new_n1107), .A3(new_n1111), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1143), .A2(new_n1155), .A3(new_n1154), .ZN(new_n1160));
  NOR2_X1   g735(.A1(G305), .A2(G1981), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1162));
  NOR2_X1   g737(.A1(G288), .A2(G1976), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1160), .B1(new_n1164), .B2(new_n1137), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT114), .B(KEYINPUT63), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1124), .A2(G168), .A3(new_n1118), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1157), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT115), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1169), .B1(new_n1170), .B2(new_n1112), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1154), .A2(KEYINPUT115), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1145), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1167), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1173), .A2(new_n1156), .A3(new_n1143), .A4(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1165), .B1(new_n1168), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1129), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1157), .A2(new_n1108), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1180), .B1(new_n1129), .B2(new_n1178), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1177), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1037), .B1(new_n1159), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1023), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1184), .A2(G1986), .A3(G290), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT48), .Z(new_n1186));
  NAND2_X1  g761(.A1(new_n1034), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1030), .B(KEYINPUT46), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1023), .B1(new_n817), .B2(new_n1026), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1190), .A2(KEYINPUT47), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(KEYINPUT47), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1187), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OR3_X1    g768(.A1(new_n1031), .A2(new_n738), .A3(new_n734), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n888), .A2(new_n832), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1184), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1183), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g773(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n1200), .A2(new_n912), .A3(new_n1009), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


