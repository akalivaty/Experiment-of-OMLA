//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n204), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT0), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n213), .A2(new_n215), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(new_n219), .B2(new_n218), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  AND2_X1   g0026(.A1(new_n226), .A2(new_n216), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n227), .A2(new_n228), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n221), .A2(new_n230), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G97), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(G223), .A3(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n250), .B(new_n251), .C1(new_n252), .C2(new_n248), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G41), .A2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n257), .A2(G1), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n257), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n254), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n259), .B1(new_n266), .B2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n255), .A2(new_n256), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n256), .B1(new_n255), .B2(new_n267), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G200), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n212), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT69), .A2(G58), .ZN(new_n275));
  XOR2_X1   g0075(.A(new_n275), .B(KEYINPUT8), .Z(new_n276));
  NAND2_X1  g0076(.A1(new_n211), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n276), .A2(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n201), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G58), .A2(G68), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n207), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n274), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n274), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT67), .B(G1), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n207), .ZN(new_n289));
  MUX2_X1   g0089(.A(new_n286), .B(new_n289), .S(G50), .Z(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT9), .ZN(new_n292));
  OAI21_X1  g0092(.A(G190), .B1(new_n269), .B2(new_n270), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n272), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n272), .A2(new_n292), .A3(new_n296), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n211), .A2(G33), .A3(G77), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n279), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n287), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT11), .ZN(new_n302));
  INV_X1    g0102(.A(G13), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n288), .A2(new_n303), .A3(new_n207), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT70), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n286), .A2(KEYINPUT70), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n287), .B(new_n305), .C1(new_n288), .C2(new_n207), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT12), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT12), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n311), .A2(G68), .B1(new_n312), .B2(new_n286), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT72), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT72), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n302), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n248), .A2(G232), .A3(G1698), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n248), .A2(G226), .A3(new_n249), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n254), .ZN(new_n323));
  INV_X1    g0123(.A(G33), .ZN(new_n324));
  INV_X1    g0124(.A(G41), .ZN(new_n325));
  OAI211_X1 g0125(.A(G1), .B(G13), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n326), .B(G238), .C1(new_n288), .C2(new_n257), .ZN(new_n327));
  INV_X1    g0127(.A(new_n259), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n327), .A2(KEYINPUT71), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT71), .B1(new_n327), .B2(new_n328), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT13), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n323), .B(new_n333), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(G190), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n318), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n332), .B2(new_n334), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n271), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n269), .B2(new_n270), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n291), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n248), .A2(G238), .A3(G1698), .ZN(new_n346));
  INV_X1    g0146(.A(G107), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n345), .B(new_n346), .C1(new_n347), .C2(new_n248), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n254), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n259), .B1(new_n266), .B2(G244), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G200), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n308), .A2(new_n252), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n310), .A2(new_n252), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT8), .B(G58), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT65), .B(G20), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n356), .A2(new_n279), .B1(new_n357), .B2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n277), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n354), .B1(new_n360), .B2(new_n274), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n349), .A2(new_n350), .A3(G190), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n352), .A2(new_n353), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n344), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n298), .A2(new_n339), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n302), .ZN(new_n366));
  INV_X1    g0166(.A(new_n317), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT72), .B1(new_n309), .B2(new_n313), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n332), .A2(G179), .A3(new_n334), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT73), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n340), .B1(new_n332), .B2(new_n334), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n370), .B(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n361), .A2(new_n353), .B1(new_n351), .B2(new_n340), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n349), .A2(new_n342), .A3(new_n350), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT18), .ZN(new_n382));
  INV_X1    g0182(.A(new_n276), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n289), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n276), .A2(new_n286), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT76), .ZN(new_n387));
  AND2_X1   g0187(.A1(G58), .A2(G68), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n283), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n279), .A2(G159), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n389), .A2(KEYINPUT75), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT75), .B1(new_n389), .B2(new_n390), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT3), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(G33), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n394), .B(new_n207), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(G33), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n208), .A2(new_n210), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(G68), .B(new_n398), .C1(new_n401), .C2(new_n394), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n387), .B(KEYINPUT16), .C1(new_n393), .C2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G58), .A2(G68), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n207), .B1(new_n204), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n390), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n389), .A2(KEYINPUT75), .A3(new_n390), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT76), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(new_n409), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n399), .A2(new_n400), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT74), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n394), .B1(new_n357), .B2(new_n248), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n415), .A2(new_n419), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n414), .B1(new_n421), .B2(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n287), .B1(new_n422), .B2(KEYINPUT16), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n386), .B1(new_n413), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n248), .A2(G226), .A3(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n248), .A2(G223), .A3(new_n249), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n254), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n259), .B1(new_n266), .B2(G232), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n340), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n429), .A2(new_n430), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(G179), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n382), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT7), .B1(new_n357), .B2(new_n248), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n435), .A2(G68), .A3(new_n398), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n411), .B1(new_n436), .B2(new_n414), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n387), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n418), .A2(new_n420), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n248), .A2(G20), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n419), .B1(new_n440), .B2(KEYINPUT7), .ZN(new_n441));
  OAI21_X1  g0241(.A(G68), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(KEYINPUT16), .A3(new_n393), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n410), .A2(KEYINPUT76), .A3(new_n411), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n438), .A2(new_n274), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n386), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n382), .B(new_n433), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n434), .B1(new_n447), .B2(KEYINPUT77), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n433), .B1(new_n445), .B2(new_n446), .ZN(new_n449));
  OR3_X1    g0249(.A1(new_n449), .A2(KEYINPUT77), .A3(KEYINPUT18), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n429), .A2(new_n430), .ZN(new_n451));
  INV_X1    g0251(.A(G190), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(G200), .B2(new_n451), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n424), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT17), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n454), .A2(new_n445), .A3(new_n446), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT17), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n448), .A2(new_n450), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n365), .B(new_n381), .C1(KEYINPUT78), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n456), .A2(new_n459), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT77), .B1(new_n449), .B2(KEYINPUT18), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n449), .A2(KEYINPUT18), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n449), .A2(KEYINPUT77), .A3(KEYINPUT18), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT78), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n287), .B1(new_n288), .B2(new_n324), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(new_n306), .A3(new_n307), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n286), .A2(KEYINPUT70), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n207), .B1(new_n261), .B2(new_n263), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n305), .B1(new_n475), .B2(G13), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n471), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n324), .A2(G97), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n211), .A2(KEYINPUT86), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT86), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n479), .B1(new_n483), .B2(G33), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n357), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n273), .A2(new_n212), .B1(G20), .B2(new_n471), .ZN(new_n486));
  AND4_X1   g0286(.A1(KEYINPUT20), .A2(new_n481), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n481), .A2(new_n485), .A3(new_n486), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n490), .B2(KEYINPUT87), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n478), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n248), .A2(G257), .A3(new_n249), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n248), .A2(G264), .A3(G1698), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n415), .A2(G303), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n254), .ZN(new_n499));
  INV_X1    g0299(.A(G45), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n261), .B2(new_n263), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT5), .B(G41), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(G274), .A3(new_n326), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n254), .B1(new_n501), .B2(new_n502), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G270), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n499), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n506), .A2(new_n342), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT88), .B1(new_n494), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n490), .A2(KEYINPUT87), .ZN(new_n509));
  INV_X1    g0309(.A(new_n487), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n493), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n478), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT88), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n506), .A2(new_n342), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT89), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n506), .A2(G169), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n518), .B(new_n519), .C1(new_n494), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n520), .B1(new_n511), .B2(new_n512), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n518), .A2(new_n519), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n470), .A2(new_n304), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n347), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT25), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n286), .B2(G107), .ZN(new_n529));
  AOI22_X1  g0329(.A1(G107), .A2(new_n526), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(KEYINPUT23), .A2(G107), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n357), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT23), .A2(G107), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(G20), .C2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G87), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(KEYINPUT90), .B2(KEYINPUT22), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n211), .A2(new_n248), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(KEYINPUT90), .B2(KEYINPUT22), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n415), .A2(new_n357), .ZN(new_n540));
  NOR2_X1   g0340(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(new_n537), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n535), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n274), .B1(new_n543), .B2(KEYINPUT24), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n530), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n399), .A2(new_n400), .A3(G257), .A4(G1698), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(KEYINPUT91), .B1(G33), .B2(G294), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n248), .A2(KEYINPUT92), .A3(G250), .A4(new_n249), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT91), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n248), .A2(new_n551), .A3(G257), .A4(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n399), .A2(new_n400), .A3(G250), .A4(new_n249), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT92), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n549), .A2(new_n550), .A3(new_n552), .A4(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n254), .B1(G264), .B2(new_n504), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n342), .A3(new_n503), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n254), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n504), .A2(G264), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n503), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n340), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n547), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n517), .A2(new_n521), .A3(new_n525), .A4(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(G257), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n565), .B(new_n254), .C1(new_n501), .C2(new_n502), .ZN(new_n566));
  INV_X1    g0366(.A(new_n503), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT80), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n399), .A2(new_n400), .A3(G244), .A4(new_n249), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT4), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n479), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n569), .A2(new_n570), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n254), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n504), .A2(G257), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT80), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n577), .A3(new_n503), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n568), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n579), .A2(G200), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n452), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT79), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n347), .A2(G97), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n483), .A2(G107), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT6), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n347), .A2(KEYINPUT6), .A3(G97), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n211), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n280), .A2(new_n252), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n582), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n589), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n347), .A2(KEYINPUT6), .A3(G97), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n245), .B2(new_n585), .ZN(new_n593));
  OAI211_X1 g0393(.A(KEYINPUT79), .B(new_n591), .C1(new_n593), .C2(new_n211), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n435), .A2(G107), .A3(new_n398), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n274), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n286), .A2(G97), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n526), .B2(G97), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n580), .A2(new_n581), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n579), .A2(new_n340), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n568), .A2(new_n575), .A3(new_n578), .A4(new_n342), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n340), .A2(new_n579), .B1(new_n597), .B2(new_n599), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(KEYINPUT81), .A3(new_n603), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT24), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n539), .A2(new_n542), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(new_n535), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n274), .A3(new_n544), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n561), .A2(G200), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n557), .A2(G190), .A3(new_n503), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n530), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n248), .A2(G244), .A3(G1698), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G33), .A2(G116), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n399), .A2(new_n400), .A3(G238), .A4(new_n249), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT83), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n617), .A2(KEYINPUT83), .A3(new_n618), .A4(new_n619), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n326), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT82), .ZN(new_n626));
  INV_X1    g0426(.A(new_n501), .ZN(new_n627));
  INV_X1    g0427(.A(G250), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n254), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n626), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NOR4_X1   g0430(.A1(new_n501), .A2(new_n254), .A3(KEYINPUT82), .A4(new_n628), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n326), .A2(G274), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n630), .A2(new_n631), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n625), .A2(new_n634), .A3(G190), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n536), .A2(new_n483), .A3(new_n347), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT19), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n321), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n357), .B2(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(KEYINPUT84), .B1(new_n540), .B2(G68), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n639), .A2(KEYINPUT84), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT85), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n357), .A2(new_n324), .A3(new_n483), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(KEYINPUT19), .ZN(new_n644));
  OAI211_X1 g0444(.A(KEYINPUT85), .B(new_n637), .C1(new_n277), .C2(new_n483), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n640), .A2(new_n641), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n646), .A2(new_n274), .B1(new_n308), .B2(new_n359), .ZN(new_n647));
  OAI21_X1  g0447(.A(G200), .B1(new_n624), .B2(new_n633), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n526), .A2(G87), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n635), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n274), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n308), .A2(new_n359), .ZN(new_n652));
  INV_X1    g0452(.A(new_n359), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n526), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n625), .A2(new_n634), .A3(new_n342), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n340), .B1(new_n624), .B2(new_n633), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n616), .A2(new_n650), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n506), .A2(G200), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n494), .B(new_n660), .C1(new_n452), .C2(new_n506), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n609), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  NOR4_X1   g0462(.A1(new_n461), .A2(new_n469), .A3(new_n564), .A4(new_n662), .ZN(G372));
  NOR2_X1   g0463(.A1(new_n461), .A2(new_n469), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n564), .A2(new_n609), .A3(new_n659), .ZN(new_n665));
  INV_X1    g0465(.A(new_n658), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n606), .A2(new_n608), .A3(new_n658), .A4(new_n650), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n650), .A2(new_n658), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n602), .A2(new_n600), .A3(KEYINPUT93), .A4(new_n603), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT93), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n604), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n669), .A2(new_n670), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n665), .A2(new_n668), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n344), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n449), .A2(KEYINPUT18), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n434), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n462), .A2(new_n339), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n381), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT94), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n298), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n295), .A2(KEYINPUT94), .A3(new_n297), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n677), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n676), .A2(new_n686), .ZN(G369));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n211), .A2(G13), .ZN(new_n689));
  OR3_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .A3(new_n288), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT27), .B1(new_n689), .B2(new_n288), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n547), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n613), .A2(new_n530), .B1(new_n340), .B2(new_n561), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n616), .A2(new_n695), .B1(new_n696), .B2(new_n558), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n563), .A2(new_n694), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT96), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n616), .A2(new_n695), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n563), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT96), .ZN(new_n702));
  INV_X1    g0502(.A(new_n694), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n696), .A2(new_n558), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n517), .A2(new_n521), .A3(new_n525), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n494), .A2(new_n703), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n661), .B1(new_n494), .B2(new_n703), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT95), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT95), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n709), .B(new_n714), .C1(new_n707), .C2(new_n711), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n688), .B(new_n706), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n707), .A2(new_n703), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n699), .A3(new_n705), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT97), .B1(new_n719), .B2(new_n704), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n719), .A2(KEYINPUT97), .A3(new_n704), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n717), .B1(new_n720), .B2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n217), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n636), .A2(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n214), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n669), .A2(new_n670), .A3(new_n606), .A4(new_n608), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n673), .A2(new_n658), .A3(new_n650), .A4(new_n671), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n666), .B1(new_n731), .B2(KEYINPUT26), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n665), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .A3(new_n703), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT100), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT100), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n733), .A2(new_n736), .A3(KEYINPUT29), .A4(new_n703), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AOI211_X1 g0538(.A(KEYINPUT99), .B(KEYINPUT29), .C1(new_n675), .C2(new_n703), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT99), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n675), .A2(new_n703), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n738), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n662), .A2(new_n564), .A3(new_n694), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n579), .A2(new_n342), .A3(new_n506), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT98), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n624), .B2(new_n633), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n624), .A2(new_n633), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT98), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n746), .A2(new_n561), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n579), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n752), .A2(new_n749), .A3(new_n515), .A4(new_n557), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n579), .A2(new_n624), .A3(new_n633), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n756), .A2(KEYINPUT30), .A3(new_n515), .A4(new_n557), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n751), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n694), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT31), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(G330), .B1(new_n745), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n744), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n729), .B1(new_n766), .B2(G1), .ZN(G364));
  INV_X1    g0567(.A(new_n689), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n260), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n724), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n713), .A2(new_n715), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(new_n772), .B2(G330), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n248), .A2(new_n217), .ZN(new_n775));
  INV_X1    g0575(.A(G355), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n776), .B1(G116), .B2(new_n217), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n415), .A2(new_n217), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT101), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n500), .B2(new_n215), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n243), .A2(G45), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n212), .B1(G20), .B2(new_n340), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n771), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G179), .A2(G200), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n357), .A2(new_n452), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n792), .A2(KEYINPUT32), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G50), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n211), .A2(new_n342), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n337), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(new_n452), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n795), .A2(new_n799), .B1(new_n802), .B2(new_n252), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n797), .A2(G200), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n794), .B(new_n803), .C1(G58), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n337), .A2(G179), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n806), .A2(G20), .A3(G190), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT102), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT102), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G87), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT32), .B1(new_n792), .B2(new_n793), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n791), .A2(G190), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n357), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n415), .B1(new_n815), .B2(G97), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n812), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n357), .A2(new_n452), .A3(new_n806), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT103), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n347), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  OR3_X1    g0621(.A1(new_n800), .A2(KEYINPUT104), .A3(new_n337), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT104), .B1(new_n800), .B2(new_n337), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n805), .B(new_n821), .C1(new_n203), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n819), .ZN(new_n827));
  INV_X1    g0627(.A(new_n792), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n827), .A2(G283), .B1(G329), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT105), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  INV_X1    g0631(.A(new_n815), .ZN(new_n832));
  INV_X1    g0632(.A(G303), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n415), .B1(new_n831), .B2(new_n832), .C1(new_n810), .C2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G322), .B2(new_n804), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G311), .A2(new_n801), .B1(new_n798), .B2(G326), .ZN(new_n836));
  XOR2_X1   g0636(.A(KEYINPUT33), .B(G317), .Z(new_n837));
  OAI211_X1 g0637(.A(new_n835), .B(new_n836), .C1(new_n825), .C2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n826), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n790), .B1(new_n839), .B2(new_n787), .ZN(new_n840));
  INV_X1    g0640(.A(new_n786), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n772), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n774), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  NAND2_X1  g0644(.A1(new_n361), .A2(new_n353), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n694), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n363), .A2(new_n846), .B1(new_n378), .B2(new_n379), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n378), .A2(new_n379), .A3(new_n703), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT107), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n363), .A2(new_n846), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n380), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT107), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(new_n853), .A3(new_n848), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n675), .A2(new_n703), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT108), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n850), .A2(new_n854), .A3(KEYINPUT108), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n675), .B2(new_n703), .ZN(new_n862));
  OR3_X1    g0662(.A1(new_n857), .A2(new_n862), .A3(new_n764), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n764), .B1(new_n857), .B2(new_n862), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n863), .B(new_n864), .C1(new_n724), .C2(new_n770), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n787), .A2(new_n784), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n771), .B1(G77), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n248), .B1(new_n815), .B2(G97), .ZN(new_n869));
  INV_X1    g0669(.A(G311), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n869), .B1(new_n870), .B2(new_n792), .C1(new_n810), .C2(new_n347), .ZN(new_n871));
  AOI22_X1  g0671(.A1(G116), .A2(new_n801), .B1(new_n798), .B2(G303), .ZN(new_n872));
  INV_X1    g0672(.A(new_n804), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n831), .B2(new_n873), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n871), .B(new_n874), .C1(G87), .C2(new_n827), .ZN(new_n875));
  INV_X1    g0675(.A(G283), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n824), .B(KEYINPUT106), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G137), .A2(new_n798), .B1(new_n804), .B2(G143), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n879), .B1(new_n793), .B2(new_n802), .C1(new_n825), .C2(new_n278), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT34), .Z(new_n881));
  OAI221_X1 g0681(.A(new_n248), .B1(new_n202), .B2(new_n832), .C1(new_n810), .C2(new_n795), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G132), .B2(new_n828), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n819), .A2(new_n203), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n878), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n868), .B1(new_n887), .B2(new_n787), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n785), .B2(new_n855), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n865), .A2(new_n889), .ZN(G384));
  INV_X1    g0690(.A(new_n593), .ZN(new_n891));
  OAI211_X1 g0691(.A(G116), .B(new_n213), .C1(new_n891), .C2(KEYINPUT35), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(KEYINPUT35), .B2(new_n891), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT36), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n215), .A2(G77), .A3(new_n405), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n282), .A2(G68), .ZN(new_n896));
  AOI211_X1 g0696(.A(G13), .B(new_n264), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n369), .B(new_n703), .C1(new_n375), .C2(new_n376), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n423), .B1(KEYINPUT16), .B2(new_n422), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n446), .ZN(new_n904));
  INV_X1    g0704(.A(new_n692), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n448), .A2(new_n450), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n907), .B2(new_n462), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n445), .A2(new_n446), .B1(new_n433), .B2(new_n692), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n911), .A3(new_n455), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n433), .A2(new_n692), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n457), .B1(new_n913), .B2(new_n904), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n914), .B2(new_n911), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n902), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(KEYINPUT38), .B(new_n915), .C1(new_n460), .C2(new_n906), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n901), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n920));
  OR2_X1    g0720(.A1(new_n424), .A2(new_n692), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n462), .B2(new_n679), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT37), .B1(new_n457), .B2(new_n909), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n912), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n918), .A2(new_n925), .A3(new_n901), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n900), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n679), .A2(new_n905), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n917), .A2(new_n918), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n336), .A2(new_n338), .B1(new_n318), .B2(new_n703), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n377), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n899), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n856), .B2(new_n848), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n928), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n738), .B(new_n664), .C1(new_n739), .C2(new_n743), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n686), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(new_n855), .A3(new_n899), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n609), .A2(new_n659), .ZN(new_n940));
  INV_X1    g0740(.A(new_n564), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n940), .A2(new_n941), .A3(new_n661), .A4(new_n703), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT110), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(KEYINPUT31), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n758), .A2(new_n694), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n758), .B2(new_n694), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n939), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n929), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT40), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n918), .A2(new_n925), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(KEYINPUT40), .A3(new_n950), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n469), .B(new_n461), .C1(new_n942), .C2(new_n949), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n931), .A2(new_n855), .A3(new_n899), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n759), .A2(new_n944), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n946), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n958), .B1(new_n745), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n917), .B2(new_n918), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n955), .B(G330), .C1(new_n962), .C2(KEYINPUT40), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n688), .B1(new_n942), .B2(new_n949), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n664), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n956), .A2(new_n957), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n938), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n264), .B2(new_n768), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n938), .A2(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n898), .B1(new_n968), .B2(new_n969), .ZN(G367));
  NAND2_X1  g0770(.A1(new_n600), .A2(new_n694), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n609), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n719), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(KEYINPUT42), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n606), .A2(new_n608), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n607), .A2(new_n603), .A3(new_n694), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n975), .B1(new_n978), .B2(new_n563), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n973), .A2(KEYINPUT42), .B1(new_n979), .B2(new_n703), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n647), .A2(new_n649), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n694), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n669), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(new_n658), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT43), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n981), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n974), .A2(new_n980), .A3(new_n988), .A4(new_n987), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n717), .A2(new_n978), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n724), .B(KEYINPUT41), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n977), .B1(new_n721), .B2(new_n720), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(KEYINPUT45), .B(new_n977), .C1(new_n721), .C2(new_n720), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n719), .A2(new_n704), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT97), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n719), .A2(KEYINPUT97), .A3(new_n704), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n1006), .A3(new_n978), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1005), .A2(new_n1006), .A3(KEYINPUT44), .A4(new_n978), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1002), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n716), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n772), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n706), .B1(new_n1014), .B2(new_n688), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n717), .A3(new_n718), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n718), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n772), .A2(G330), .B1(new_n699), .B2(new_n705), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n716), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n1019), .A3(new_n744), .A4(new_n764), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1002), .A2(new_n1011), .A3(new_n717), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1013), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n997), .B1(new_n1023), .B2(new_n766), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n995), .B1(new_n1024), .B2(new_n770), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n788), .B1(new_n217), .B2(new_n359), .C1(new_n780), .C2(new_n239), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n771), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n828), .A2(G137), .B1(G68), .B2(new_n815), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n818), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n415), .B1(new_n1029), .B2(G77), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1028), .B1(new_n810), .B2(new_n202), .C1(new_n1030), .C2(KEYINPUT112), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G143), .A2(new_n798), .B1(new_n801), .B2(new_n201), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n278), .B2(new_n873), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1031), .B(new_n1033), .C1(KEYINPUT112), .C2(new_n1030), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n793), .B2(new_n877), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n811), .A2(G116), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT46), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1036), .A2(new_n1037), .B1(new_n801), .B2(G283), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n833), .B2(new_n873), .ZN(new_n1039));
  XOR2_X1   g0839(.A(KEYINPUT111), .B(G317), .Z(new_n1040));
  NAND2_X1  g0840(.A1(new_n828), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n248), .B1(new_n815), .B2(G107), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n483), .C2(new_n818), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1036), .A2(new_n1037), .B1(new_n870), .B2(new_n799), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1039), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n877), .B2(new_n831), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT47), .B1(new_n1035), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n787), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1035), .A2(KEYINPUT47), .A3(new_n1046), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1027), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n841), .B2(new_n986), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1025), .A2(new_n1052), .ZN(G387));
  NAND2_X1  g0853(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n765), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1055), .A2(new_n724), .A3(new_n1020), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1016), .A2(new_n1019), .A3(new_n770), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n779), .B1(new_n236), .B2(new_n500), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n726), .B2(new_n775), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n356), .A2(new_n795), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT50), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(KEYINPUT50), .ZN(new_n1062));
  AOI21_X1  g0862(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1061), .A2(new_n726), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1059), .A2(new_n1064), .B1(new_n347), .B2(new_n723), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n771), .B1(new_n1065), .B2(new_n789), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n706), .B2(new_n786), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n811), .A2(G77), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n415), .B1(new_n815), .B2(new_n653), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n278), .C2(new_n792), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G97), .B2(new_n827), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G50), .A2(new_n804), .B1(new_n798), .B2(G159), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n203), .C2(new_n802), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n383), .B2(new_n824), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G303), .A2(new_n801), .B1(new_n804), .B2(new_n1040), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n877), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1076), .A2(G311), .B1(G322), .B2(new_n798), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1077), .A2(KEYINPUT113), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(KEYINPUT113), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n811), .A2(G294), .B1(G283), .B2(new_n815), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT49), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n248), .B1(new_n828), .B2(G326), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n471), .B2(new_n818), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1074), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1067), .B1(new_n1091), .B2(new_n1048), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1056), .A2(new_n1057), .A3(new_n1092), .ZN(G393));
  AND2_X1   g0893(.A1(new_n1023), .A2(new_n724), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1013), .A2(new_n1022), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n1021), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G311), .A2(new_n804), .B1(new_n798), .B2(G317), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n828), .A2(G322), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n248), .B1(new_n815), .B2(G116), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n810), .C2(new_n876), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1101), .B(new_n820), .C1(G294), .C2(new_n801), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1098), .B(new_n1102), .C1(new_n877), .C2(new_n833), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n815), .A2(G77), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n355), .B2(new_n802), .C1(new_n877), .C2(new_n282), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G150), .A2(new_n798), .B1(new_n804), .B2(G159), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT115), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1108), .A2(KEYINPUT51), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(KEYINPUT51), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n415), .B1(new_n828), .B2(G143), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n810), .B2(new_n203), .C1(new_n819), .C2(new_n536), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT116), .Z(new_n1113));
  NOR4_X1   g0913(.A1(new_n1106), .A2(new_n1109), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n787), .B1(new_n1104), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n788), .B1(new_n483), .B2(new_n217), .C1(new_n780), .C2(new_n246), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n771), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n786), .B2(new_n978), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1095), .B2(new_n770), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1096), .A2(new_n1119), .ZN(G390));
  OAI211_X1 g0920(.A(G330), .B(new_n861), .C1(new_n745), .C2(new_n960), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(KEYINPUT118), .A3(new_n932), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n733), .A2(new_n703), .A3(new_n855), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n848), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n958), .C1(new_n745), .C2(new_n763), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(KEYINPUT118), .A2(new_n1127), .B1(new_n1121), .B2(new_n932), .ZN(new_n1128));
  OAI211_X1 g0928(.A(G330), .B(new_n855), .C1(new_n745), .C2(new_n763), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1129), .A2(new_n932), .B1(new_n964), .B2(new_n958), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n856), .A2(new_n848), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1126), .A2(new_n1128), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1133), .A2(new_n686), .A3(new_n965), .A4(new_n936), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n906), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n467), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT38), .B1(new_n1136), .B2(new_n915), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n918), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT39), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n918), .A2(new_n925), .A3(new_n901), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n900), .C2(new_n933), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1124), .A2(new_n931), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n900), .B1(new_n918), .B2(new_n925), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1141), .A2(new_n1144), .A3(new_n1127), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n964), .A2(new_n958), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1134), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1146), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n932), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n900), .B1(new_n1131), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1151), .A2(new_n919), .A3(new_n926), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1144), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n936), .A2(new_n686), .A3(new_n965), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1144), .B(new_n1127), .C1(new_n1156), .C2(new_n1151), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .A4(new_n1133), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1148), .A2(new_n1158), .A3(new_n724), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n919), .A2(new_n926), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1151), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1160), .A2(new_n1161), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1157), .B(new_n770), .C1(new_n1162), .C2(new_n1146), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n771), .B1(new_n383), .B2(new_n867), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1076), .A2(G137), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n810), .A2(new_n278), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1167), .A2(KEYINPUT53), .B1(new_n798), .B2(G128), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT54), .B(G143), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n801), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT53), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1166), .A2(new_n1171), .B1(G132), .B2(new_n804), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n248), .B1(new_n818), .B2(new_n282), .C1(new_n832), .C2(new_n793), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G125), .B2(new_n828), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1168), .A2(new_n1170), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n877), .A2(new_n347), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n812), .A2(new_n415), .A3(new_n1105), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G294), .B2(new_n828), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n801), .A2(G97), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G116), .A2(new_n804), .B1(new_n798), .B2(G283), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1178), .A2(new_n885), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n1165), .A2(new_n1175), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1164), .B1(new_n1182), .B2(new_n787), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1156), .B2(new_n785), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1163), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1159), .A2(new_n1185), .ZN(G378));
  NAND2_X1  g0986(.A1(new_n291), .A2(new_n905), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n685), .B2(new_n344), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n685), .A2(new_n344), .A3(new_n1187), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1191), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1187), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n677), .B(new_n1194), .C1(new_n683), .C2(new_n684), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1188), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n953), .A2(G330), .A3(new_n1197), .A4(new_n955), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n963), .A2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n935), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1198), .A2(new_n1200), .B1(new_n927), .B2(new_n934), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n770), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1197), .A2(new_n785), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n248), .A2(G41), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G50), .B(new_n1205), .C1(new_n324), .C2(new_n325), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n818), .A2(new_n202), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G283), .B2(new_n828), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1068), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n653), .B2(new_n801), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n804), .A2(G107), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT119), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n799), .A2(new_n471), .B1(new_n203), .B2(new_n832), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT120), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1213), .A2(KEYINPUT120), .B1(new_n824), .B2(G97), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1210), .A2(new_n1212), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT58), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1206), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n811), .A2(new_n1169), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT121), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1219), .A2(new_n1220), .B1(new_n278), .B2(new_n832), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1219), .A2(new_n1220), .B1(new_n804), .B2(G128), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G125), .A2(new_n798), .B1(new_n801), .B2(G137), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1221), .B(new_n1224), .C1(G132), .C2(new_n824), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT59), .Z(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n828), .C2(G124), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n793), .B2(new_n818), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1218), .B1(new_n1217), .B2(new_n1216), .C1(new_n1226), .C2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n787), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1230), .B(new_n771), .C1(new_n201), .C2(new_n867), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1204), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1203), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1158), .A2(new_n1155), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n927), .A2(new_n934), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n963), .A2(new_n1199), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n963), .A2(new_n1199), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n935), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT57), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n724), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1158), .A2(new_n1155), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(KEYINPUT57), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1235), .B1(new_n1245), .B2(new_n1247), .ZN(G375));
  AOI21_X1  g1048(.A(new_n248), .B1(new_n815), .B2(new_n653), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n833), .B2(new_n792), .C1(new_n810), .C2(new_n483), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G107), .A2(new_n801), .B1(new_n798), .B2(G294), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n876), .B2(new_n873), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1250), .B(new_n1252), .C1(G77), .C2(new_n827), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1076), .A2(G116), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1076), .A2(new_n1169), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n415), .B(new_n1207), .C1(G50), .C2(new_n815), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n811), .A2(G159), .B1(G128), .B2(new_n828), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G132), .A2(new_n798), .B1(new_n804), .B2(G137), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n801), .A2(G150), .ZN(new_n1259));
  AND4_X1   g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1253), .A2(new_n1254), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n771), .B1(G68), .B2(new_n867), .C1(new_n1261), .C2(new_n1048), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT122), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n785), .B2(new_n1150), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1121), .A2(new_n932), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1127), .A2(KEYINPUT118), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1129), .A2(new_n932), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1146), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1265), .A2(new_n1268), .B1(new_n1131), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1264), .B1(new_n1271), .B2(new_n769), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1134), .A2(new_n996), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n936), .A2(new_n686), .A3(new_n965), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1271), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1272), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(G381));
  INV_X1    g1078(.A(G390), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1277), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT123), .Z(new_n1282));
  AOI21_X1  g1082(.A(new_n725), .B1(new_n1246), .B2(KEYINPUT57), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1234), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G378), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G387), .A2(new_n1280), .A3(new_n1282), .A4(new_n1287), .ZN(G407));
  INV_X1    g1088(.A(G213), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(G343), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1285), .A2(new_n1286), .A3(new_n1290), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1291), .A2(KEYINPUT124), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(KEYINPUT124), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(G407), .A2(G213), .A3(new_n1292), .A4(new_n1293), .ZN(G409));
  XNOR2_X1  g1094(.A(G393), .B(new_n843), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1295), .B1(G387), .B2(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G393), .B(G396), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(new_n1052), .B2(new_n1025), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1279), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G387), .A2(new_n1295), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT126), .B1(new_n1025), .B2(new_n1052), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1301), .B(G390), .C1(new_n1302), .C2(new_n1295), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1290), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1243), .A2(new_n997), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1159), .A2(new_n1203), .A3(new_n1185), .A4(new_n1233), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(G375), .B2(G378), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT60), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1276), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n725), .B1(new_n1155), .B2(new_n1133), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1271), .A2(new_n1275), .A3(KEYINPUT60), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1272), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G384), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n865), .A2(KEYINPUT125), .A3(new_n889), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1317), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1320), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1315), .A2(new_n1316), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1290), .A2(G2897), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1327), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1323), .A2(new_n1329), .A3(new_n1325), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1305), .B1(new_n1310), .B2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1304), .A2(new_n1332), .ZN(new_n1333));
  AND4_X1   g1133(.A1(new_n1159), .A2(new_n1203), .A3(new_n1185), .A4(new_n1233), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1246), .A2(new_n996), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1290), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1336), .B(new_n1326), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1337), .B(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1336), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1325), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1321), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1327), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1329), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT61), .B1(new_n1340), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1337), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G375), .A2(G378), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1349), .A2(KEYINPUT63), .A3(new_n1336), .A4(new_n1326), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1346), .A2(new_n1348), .A3(new_n1350), .ZN(new_n1351));
  AOI22_X1  g1151(.A1(new_n1333), .A2(new_n1339), .B1(new_n1351), .B2(new_n1304), .ZN(G405));
  NAND2_X1  g1152(.A1(new_n1349), .A2(new_n1287), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1326), .A2(KEYINPUT127), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1349), .A2(new_n1287), .A3(new_n1354), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1304), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1356), .A2(new_n1300), .A3(new_n1303), .A4(new_n1357), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(G402));
endmodule


