//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n206), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n212), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n211), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT64), .Z(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n221), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n217), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT66), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT67), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT8), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT68), .B1(new_n212), .B2(KEYINPUT8), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(new_n254), .A3(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT69), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n206), .A2(KEYINPUT69), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G150), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR3_X1   g0070(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n268), .A2(new_n270), .B1(new_n271), .B2(new_n206), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n252), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n205), .A2(G20), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n251), .A2(G50), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n274), .A2(new_n206), .A3(G1), .ZN(new_n279));
  INV_X1    g0079(.A(G50), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n278), .A2(KEYINPUT70), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT70), .B1(new_n278), .B2(new_n281), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n273), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT9), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT9), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n286), .B(new_n273), .C1(new_n282), .C2(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n262), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n293), .A2(G223), .B1(new_n296), .B2(G77), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1698), .B1(new_n291), .B2(new_n292), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G222), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G1), .A3(G13), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  INV_X1    g0105(.A(G45), .ZN(new_n306));
  AOI21_X1  g0106(.A(G1), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(new_n302), .A3(G274), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n303), .A2(new_n307), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(G226), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n304), .B2(new_n311), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n288), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT75), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT74), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n285), .A2(new_n322), .A3(new_n287), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n314), .A2(KEYINPUT10), .A3(new_n316), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n285), .B2(new_n287), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n321), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n326), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n328), .A2(KEYINPUT75), .A3(new_n323), .A4(new_n324), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n320), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n284), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n312), .A2(G179), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT71), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  AOI211_X1 g0134(.A(new_n331), .B(new_n333), .C1(new_n334), .C2(new_n312), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n277), .B1(new_n255), .B2(new_n259), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n248), .A2(new_n217), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n250), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n249), .A2(KEYINPUT66), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n276), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n260), .A2(new_n279), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT83), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n345), .B(KEYINPUT83), .C1(new_n342), .C2(new_n337), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT82), .ZN(new_n350));
  AND2_X1   g0150(.A1(KEYINPUT67), .A2(G58), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT67), .A2(G58), .ZN(new_n352));
  OAI21_X1  g0152(.A(G68), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n206), .B1(new_n353), .B2(new_n214), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  INV_X1    g0155(.A(G159), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n270), .A2(new_n356), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n292), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n294), .A2(new_n295), .A3(G20), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT79), .B1(new_n361), .B2(KEYINPUT7), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n291), .A2(new_n206), .A3(new_n292), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT79), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n360), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n358), .B1(new_n367), .B2(new_n213), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n249), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(new_n365), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(KEYINPUT81), .A3(new_n359), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT81), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n361), .A2(new_n374), .A3(KEYINPUT7), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(G68), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n354), .A2(new_n357), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n350), .B1(new_n369), .B2(new_n378), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n364), .B1(new_n363), .B2(new_n365), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n359), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G68), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n339), .B1(new_n383), .B2(new_n358), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n376), .A2(new_n377), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n370), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(KEYINPUT82), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n349), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n298), .A2(G223), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n291), .A2(new_n292), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(G226), .A3(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(G179), .B1(new_n393), .B2(new_n303), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n302), .A2(G232), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT84), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n302), .A2(new_n395), .A3(KEYINPUT84), .A4(G232), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n308), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT85), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n398), .A2(KEYINPUT85), .A3(new_n308), .A4(new_n399), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n394), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n293), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n302), .B1(new_n405), .B2(new_n389), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n334), .B1(new_n406), .B2(new_n400), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT18), .B1(new_n388), .B2(new_n408), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n346), .A2(new_n348), .ZN(new_n410));
  AOI21_X1  g0210(.A(G190), .B1(new_n393), .B2(new_n303), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(new_n402), .A3(new_n403), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n315), .B1(new_n406), .B2(new_n400), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n369), .A2(new_n350), .A3(new_n378), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT82), .B1(new_n384), .B2(new_n386), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n410), .B(new_n415), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n410), .B1(new_n416), .B2(new_n417), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(new_n408), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n388), .A2(KEYINPUT17), .A3(new_n415), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n409), .A2(new_n420), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n427));
  INV_X1    g0227(.A(G77), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n266), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n252), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT11), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n252), .A2(KEYINPUT11), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n339), .A2(new_n276), .ZN(new_n434));
  INV_X1    g0234(.A(new_n277), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n434), .A2(new_n213), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT12), .B1(new_n276), .B2(G68), .ZN(new_n437));
  OR3_X1    g0237(.A1(new_n276), .A2(KEYINPUT12), .A3(G68), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n432), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n298), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n390), .A2(G232), .A3(G1698), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n302), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n307), .A2(new_n302), .A3(new_n446), .A4(G274), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n302), .A2(G238), .A3(new_n395), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT13), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n390), .A2(G226), .A3(new_n289), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G97), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n443), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n303), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT13), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n334), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT14), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n450), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n450), .A2(new_n461), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(G179), .A4(new_n457), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n450), .A2(new_n457), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n459), .A3(G169), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT78), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n441), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n462), .A2(new_n463), .A3(G190), .A4(new_n457), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n440), .B1(new_n466), .B2(G200), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G179), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n293), .A2(G238), .B1(new_n296), .B2(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n390), .A2(G232), .A3(new_n289), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n303), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT72), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n309), .B1(G244), .B2(new_n310), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n474), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n483), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(new_n334), .A3(new_n481), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n434), .A2(new_n428), .A3(new_n435), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT73), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n279), .A2(new_n428), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT15), .B(G87), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n266), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT8), .B(G58), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n492), .A2(new_n270), .B1(new_n206), .B2(new_n428), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n249), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n488), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n484), .A2(new_n486), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(G190), .B1(new_n482), .B2(new_n483), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n485), .A2(G200), .A3(new_n481), .ZN(new_n498));
  INV_X1    g0298(.A(new_n495), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NOR4_X1   g0301(.A1(new_n426), .A2(new_n469), .A3(new_n473), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n336), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(new_n206), .C1(G33), .C2(new_n222), .ZN(new_n505));
  INV_X1    g0305(.A(G116), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n249), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n275), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n507), .ZN(new_n512));
  INV_X1    g0312(.A(new_n434), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n506), .B1(new_n205), .B2(G33), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT89), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n298), .A2(new_n517), .A3(G257), .ZN(new_n518));
  OAI211_X1 g0318(.A(G257), .B(new_n289), .C1(new_n294), .C2(new_n295), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT89), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n293), .A2(G264), .B1(new_n296), .B2(G303), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n302), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT5), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT87), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(G41), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n305), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n306), .A2(G1), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n530), .A2(G270), .A3(new_n302), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n302), .A2(G274), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n516), .A2(new_n524), .A3(G179), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n390), .A2(G264), .A3(G1698), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n296), .A2(G303), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n518), .B2(new_n520), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n534), .B1(new_n539), .B2(new_n302), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n334), .B1(new_n510), .B2(new_n515), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n535), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n206), .B(G87), .C1(new_n294), .C2(new_n295), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT22), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n390), .A2(new_n548), .A3(new_n206), .A4(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n206), .B2(G107), .ZN(new_n553));
  INV_X1    g0353(.A(G107), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(KEYINPUT23), .A3(G20), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n262), .A2(new_n506), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n553), .A2(new_n555), .B1(new_n556), .B2(new_n206), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n550), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n551), .B1(new_n550), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n249), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT90), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT90), .B(new_n249), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n251), .B(new_n276), .C1(G1), .C2(new_n262), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n554), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n279), .A2(new_n554), .ZN(new_n567));
  XNOR2_X1  g0367(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G250), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n223), .B2(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n390), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G294), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n302), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n530), .A2(G264), .A3(new_n302), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n576), .A2(new_n577), .A3(new_n533), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n474), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n530), .A2(new_n532), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n530), .A2(G264), .A3(new_n302), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n573), .A2(new_n390), .B1(G33), .B2(G294), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n581), .C1(new_n302), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n334), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n545), .B1(new_n571), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(new_n289), .C1(new_n294), .C2(new_n295), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT86), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT4), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(KEYINPUT86), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n293), .A2(G250), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n590), .A2(new_n592), .A3(new_n504), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n303), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n530), .A2(new_n302), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G257), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n580), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n279), .A2(new_n222), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n565), .B2(new_n222), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n373), .A2(G107), .A3(new_n375), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n554), .A2(KEYINPUT6), .A3(G97), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n222), .A2(new_n554), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n202), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n605), .B2(KEYINPUT6), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G20), .B1(G77), .B2(new_n269), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n339), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n599), .B(new_n609), .C1(new_n313), .C2(new_n598), .ZN(new_n610));
  INV_X1    g0410(.A(new_n609), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n598), .A2(new_n334), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n594), .A2(new_n303), .B1(G257), .B2(new_n596), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n474), .A3(new_n580), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n556), .B1(new_n293), .B2(G244), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n298), .A2(G238), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n303), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT88), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n529), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n205), .A2(G45), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT88), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n622), .A2(new_n624), .A3(G250), .A4(new_n302), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n302), .A2(G274), .A3(new_n529), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G200), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n390), .A2(new_n206), .A3(G68), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT19), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n206), .B1(new_n453), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(G87), .B2(new_n203), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT19), .B1(new_n265), .B2(G97), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n249), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n490), .A2(new_n279), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G87), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n565), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n627), .B1(new_n619), .B2(new_n303), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G190), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n630), .A2(new_n639), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n629), .A2(new_n334), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n637), .B(new_n638), .C1(new_n565), .C2(new_n490), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n474), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n570), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n562), .B2(new_n563), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n583), .A2(new_n313), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(G200), .B2(new_n583), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n516), .B1(new_n540), .B2(G200), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n313), .B2(new_n540), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n587), .A2(new_n616), .A3(new_n654), .A4(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n503), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT92), .Z(G372));
  INV_X1    g0459(.A(new_n496), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n469), .B1(new_n660), .B2(new_n472), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n420), .A2(new_n425), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n409), .B(new_n424), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n330), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n335), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n648), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n644), .A2(new_n648), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n609), .B1(new_n334), .B2(new_n598), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT26), .A4(new_n614), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n615), .B2(new_n649), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n666), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n651), .A2(new_n585), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n545), .A2(KEYINPUT93), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n545), .A2(KEYINPUT93), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n616), .A2(new_n654), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n665), .B1(new_n503), .B2(new_n679), .ZN(G369));
  INV_X1    g0480(.A(new_n535), .ZN(new_n681));
  INV_X1    g0481(.A(new_n544), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n510), .ZN(new_n685));
  INV_X1    g0485(.A(new_n515), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OR3_X1    g0487(.A1(new_n511), .A2(KEYINPUT27), .A3(G20), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT27), .B1(new_n511), .B2(G20), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(G213), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n656), .B1(new_n684), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n674), .A2(new_n675), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT94), .Z(new_n698));
  NAND2_X1  g0498(.A1(new_n673), .A2(new_n693), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n673), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n651), .A2(new_n653), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n651), .B2(new_n693), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n700), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n698), .A2(G330), .A3(new_n704), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n684), .A2(new_n692), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n700), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n209), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n215), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n678), .A2(new_n693), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n587), .A2(KEYINPUT97), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n616), .B(new_n654), .C1(new_n587), .C2(KEYINPUT97), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT96), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n723), .A2(new_n724), .B1(new_n725), .B2(new_n672), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n672), .A2(new_n725), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n693), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n721), .B1(new_n728), .B2(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n531), .A2(new_n474), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n524), .A2(new_n642), .A3(new_n578), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n595), .A2(new_n597), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n578), .A2(new_n642), .A3(G179), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(new_n598), .A3(new_n540), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n531), .A2(new_n474), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n523), .A2(new_n738), .A3(new_n583), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(KEYINPUT30), .A3(new_n613), .A4(new_n642), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT31), .B1(new_n741), .B2(new_n692), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n657), .B2(new_n692), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n730), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n719), .B1(new_n747), .B2(G1), .ZN(G364));
  NAND2_X1  g0548(.A1(new_n698), .A2(G330), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT98), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n698), .A2(KEYINPUT98), .A3(G330), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n274), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n205), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n714), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n698), .A2(G330), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n753), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n697), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n217), .B1(G20), .B2(new_n334), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n206), .A2(G179), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G190), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT32), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n771), .A3(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n206), .A2(new_n474), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n313), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n773), .B(KEYINPUT99), .Z(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n768), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n772), .B1(new_n280), .B2(new_n776), .C1(new_n779), .C2(new_n428), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n313), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(new_n253), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n767), .A2(new_n313), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n554), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n767), .A2(G190), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n640), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n786), .A2(new_n788), .A3(new_n296), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT100), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n206), .B1(new_n781), .B2(new_n474), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n222), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n771), .B1(new_n770), .B2(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n774), .A2(G190), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(G68), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n784), .A2(new_n790), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  INV_X1    g0598(.A(G329), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n785), .A2(new_n798), .B1(new_n769), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n779), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(new_n801), .B2(G311), .ZN(new_n802));
  INV_X1    g0602(.A(G294), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(KEYINPUT33), .A2(G317), .ZN(new_n805));
  NAND2_X1  g0605(.A1(KEYINPUT33), .A2(G317), .ZN(new_n806));
  AOI211_X1 g0606(.A(G190), .B(new_n774), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(G326), .C2(new_n775), .ZN(new_n808));
  INV_X1    g0608(.A(G303), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n296), .B1(new_n787), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT101), .Z(new_n811));
  NAND2_X1  g0611(.A1(new_n783), .A2(G322), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n802), .A2(new_n808), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n766), .B1(new_n797), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n713), .A2(new_n390), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n306), .B2(new_n216), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n306), .B2(new_n243), .ZN(new_n818));
  INV_X1    g0618(.A(G355), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n209), .A2(new_n390), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(G116), .B2(new_n209), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n762), .A2(new_n765), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n757), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n764), .A2(new_n814), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n759), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n495), .A2(new_n692), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n496), .A2(new_n500), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT105), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n496), .A2(new_n500), .A3(KEYINPUT105), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n678), .A2(new_n693), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n720), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n660), .A2(new_n692), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n832), .A2(new_n837), .A3(new_n833), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT106), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n835), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n745), .A2(G330), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n757), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n766), .A2(new_n761), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n757), .B1(G77), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n801), .A2(G116), .B1(new_n783), .B2(G294), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n785), .A2(new_n640), .ZN(new_n848));
  INV_X1    g0648(.A(G311), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n793), .B1(new_n849), .B2(new_n769), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n848), .B(new_n850), .C1(G303), .C2(new_n775), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n795), .A2(KEYINPUT102), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n795), .A2(KEYINPUT102), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n787), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n390), .B1(new_n856), .B2(G107), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n855), .A2(G283), .B1(KEYINPUT103), .B2(new_n857), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n847), .A2(new_n851), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n795), .A2(G150), .B1(new_n775), .B2(G137), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n779), .B2(new_n356), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G143), .B2(new_n783), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT34), .Z(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(KEYINPUT104), .ZN(new_n866));
  INV_X1    g0666(.A(G132), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n390), .B1(new_n769), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n253), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n869), .A2(new_n791), .B1(new_n787), .B2(new_n280), .ZN(new_n870));
  INV_X1    g0670(.A(new_n785), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n868), .B(new_n870), .C1(G68), .C2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n865), .B2(KEYINPUT104), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n860), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n846), .B1(new_n874), .B2(new_n765), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n761), .B2(new_n838), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n844), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(G384));
  OAI211_X1 g0678(.A(G116), .B(new_n218), .C1(new_n606), .C2(KEYINPUT35), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n879), .A2(KEYINPUT107), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(KEYINPUT107), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT36), .Z(new_n884));
  NAND3_X1  g0684(.A1(new_n216), .A2(G77), .A3(new_n353), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n280), .A2(G68), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n205), .B(G13), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n665), .ZN(new_n889));
  INV_X1    g0689(.A(new_n503), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n730), .B2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT111), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n354), .A2(new_n357), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n382), .B2(G68), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n252), .B(new_n368), .C1(new_n894), .C2(new_n371), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n344), .A2(new_n345), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n895), .A2(new_n896), .B1(new_n408), .B2(new_n690), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n388), .B2(new_n415), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT109), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n421), .A2(new_n423), .ZN(new_n901));
  INV_X1    g0701(.A(new_n690), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n421), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n901), .A2(new_n903), .A3(new_n899), .A4(new_n418), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT109), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n414), .B(new_n349), .C1(new_n379), .C2(new_n387), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n905), .B(KEYINPUT37), .C1(new_n906), .C2(new_n897), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n900), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n690), .B1(new_n895), .B2(new_n896), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n409), .A2(new_n424), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(new_n662), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n908), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n908), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n908), .A2(new_n911), .A3(KEYINPUT38), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n418), .B1(new_n388), .B2(new_n408), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n388), .A2(new_n690), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT37), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n904), .A2(new_n919), .B1(new_n426), .B2(new_n918), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n915), .B(new_n916), .C1(KEYINPUT38), .C2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(KEYINPUT110), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT78), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n458), .A2(new_n923), .A3(new_n459), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n458), .B2(new_n459), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n460), .B(new_n464), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n440), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n692), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT110), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(KEYINPUT39), .C1(new_n912), .C2(new_n913), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n922), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n908), .A2(new_n911), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n915), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n441), .A2(new_n693), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n927), .A2(new_n472), .A3(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n440), .B(new_n692), .C1(new_n926), .C2(new_n473), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n660), .A2(new_n693), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT108), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n835), .B2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n935), .A2(new_n943), .B1(new_n910), .B2(new_n690), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n931), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n892), .B(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n919), .A2(new_n904), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n426), .A2(new_n918), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT38), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT112), .B1(new_n912), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT112), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n915), .B(new_n952), .C1(KEYINPUT38), .C2(new_n920), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n938), .A2(new_n939), .ZN(new_n954));
  AND4_X1   g0754(.A1(KEYINPUT40), .A2(new_n745), .A3(new_n954), .A4(new_n838), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n745), .A2(new_n954), .A3(new_n838), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n912), .B2(new_n913), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n890), .A2(new_n745), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(G330), .A3(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT113), .Z(new_n966));
  OR2_X1    g0766(.A1(new_n947), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT114), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n947), .A2(new_n966), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n205), .C2(new_n754), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n967), .A2(KEYINPUT114), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n888), .B1(new_n970), .B2(new_n971), .ZN(G367));
  INV_X1    g0772(.A(new_n490), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n824), .B1(new_n713), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n815), .A2(new_n238), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n714), .B(new_n756), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n693), .B1(new_n641), .B2(new_n639), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n666), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n649), .B2(new_n977), .ZN(new_n979));
  INV_X1    g0779(.A(G137), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n390), .B1(new_n769), .B2(new_n980), .C1(new_n869), .C2(new_n787), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n783), .B2(G150), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n855), .A2(G159), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n801), .A2(G50), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n785), .A2(new_n428), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n791), .A2(new_n213), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G143), .C2(new_n775), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n776), .A2(new_n849), .B1(new_n554), .B2(new_n791), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n801), .B2(G283), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n785), .A2(new_n222), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n390), .B(new_n991), .C1(G317), .C2(new_n770), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT119), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(KEYINPUT119), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n855), .A2(G294), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n856), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT46), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n787), .B2(new_n506), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(new_n782), .C2(new_n809), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n988), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT47), .Z(new_n1002));
  OAI221_X1 g0802(.A(new_n976), .B1(new_n979), .B2(new_n763), .C1(new_n1002), .C2(new_n766), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n616), .B1(new_n609), .B2(new_n693), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n668), .A2(new_n614), .A3(new_n692), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n711), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT45), .Z(new_n1008));
  NOR2_X1   g0808(.A1(new_n711), .A2(new_n1006), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT44), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n708), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n706), .A3(new_n1010), .A4(new_n707), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n751), .A2(new_n752), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n704), .B(new_n709), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT117), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n749), .A2(new_n1017), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT118), .Z(new_n1021));
  INV_X1    g0821(.A(KEYINPUT117), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1022), .A3(new_n1017), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1021), .A3(new_n747), .A4(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n747), .B1(new_n1015), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n714), .B(KEYINPUT41), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n756), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n710), .A2(new_n1006), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n615), .B1(new_n1004), .B2(new_n701), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1029), .A2(KEYINPUT42), .B1(new_n693), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT115), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1029), .A2(KEYINPUT42), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1031), .B2(KEYINPUT115), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT116), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n979), .B(KEYINPUT43), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1038), .B(new_n1039), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n708), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1042), .B(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1003), .B1(new_n1028), .B2(new_n1045), .ZN(G387));
  NAND3_X1  g0846(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n755), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n704), .A2(new_n763), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n820), .A2(new_n716), .B1(G107), .B2(new_n209), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n235), .A2(new_n306), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n716), .ZN(new_n1052));
  AOI211_X1 g0852(.A(G45), .B(new_n1052), .C1(G68), .C2(G77), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n492), .A2(G50), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT50), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n816), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1050), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n757), .B1(new_n1057), .B2(new_n824), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n801), .A2(G68), .B1(new_n783), .B2(G50), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n787), .A2(new_n428), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n791), .A2(new_n490), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(G159), .C2(new_n775), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n260), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n795), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n296), .B(new_n991), .C1(G150), .C2(new_n770), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1059), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n390), .B1(new_n770), .B2(G326), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n791), .A2(new_n798), .B1(new_n787), .B2(new_n803), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n801), .A2(G303), .B1(G322), .B2(new_n775), .ZN(new_n1069));
  INV_X1    g0869(.A(G317), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1069), .B1(new_n849), .B2(new_n854), .C1(new_n1070), .C2(new_n782), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1068), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1067), .B1(new_n506), .B2(new_n785), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1066), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT120), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n766), .B1(new_n1078), .B2(KEYINPUT120), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1058), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1048), .B1(new_n1049), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1047), .B1(new_n746), .B2(new_n730), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(new_n714), .A3(new_n1024), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(G393));
  NAND2_X1  g0885(.A1(new_n1014), .A2(new_n756), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n823), .B1(new_n222), .B2(new_n209), .C1(new_n816), .C2(new_n246), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n757), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n782), .A2(new_n849), .B1(new_n1070), .B2(new_n776), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT52), .Z(new_n1090));
  AOI211_X1 g0890(.A(new_n390), .B(new_n786), .C1(G322), .C2(new_n770), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n791), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1092), .A2(G116), .B1(new_n856), .B2(G283), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n803), .B2(new_n779), .C1(new_n809), .C2(new_n854), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n782), .A2(new_n356), .B1(new_n268), .B2(new_n776), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT51), .Z(new_n1097));
  AOI211_X1 g0897(.A(new_n296), .B(new_n848), .C1(G143), .C2(new_n770), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1092), .A2(G77), .B1(new_n856), .B2(G68), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n280), .B2(new_n854), .C1(new_n492), .C2(new_n779), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1090), .A2(new_n1095), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1088), .B1(new_n1102), .B2(new_n765), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1006), .B2(new_n763), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1014), .A2(new_n747), .A3(new_n1105), .A4(new_n1019), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n714), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1086), .B(new_n1104), .C1(new_n1107), .C2(new_n1108), .ZN(G390));
  OAI21_X1  g0909(.A(new_n757), .B1(new_n1063), .B2(new_n845), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n390), .B1(new_n769), .B2(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n791), .A2(new_n356), .B1(new_n785), .B2(new_n280), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(G128), .C2(new_n775), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1114), .B1(new_n867), .B2(new_n782), .C1(new_n779), .C2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n787), .A2(new_n268), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT53), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n854), .B2(new_n980), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n390), .B(new_n788), .C1(G294), .C2(new_n770), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n782), .B2(new_n506), .C1(new_n222), .C2(new_n779), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1092), .A2(G77), .B1(new_n871), .B2(G68), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n798), .B2(new_n776), .C1(new_n854), .C2(new_n554), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1116), .A2(new_n1119), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1110), .B1(new_n1124), .B2(new_n765), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n930), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n929), .B1(new_n935), .B2(KEYINPUT39), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n921), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1125), .B1(new_n1128), .B2(new_n761), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n746), .A2(new_n838), .A3(new_n954), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n693), .B(new_n834), .C1(new_n726), .C2(new_n727), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n941), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n954), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n928), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1133), .A2(new_n951), .A3(new_n953), .A4(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n943), .A2(new_n928), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1130), .B(new_n1135), .C1(new_n1128), .C2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n838), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n842), .A2(new_n1138), .A3(new_n940), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1136), .B1(new_n922), .B2(new_n930), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n951), .A2(new_n953), .A3(new_n1134), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n940), .B1(new_n1131), .B2(new_n941), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1139), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1137), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1129), .B1(new_n1145), .B2(new_n755), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT121), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1137), .A2(KEYINPUT121), .A3(new_n1144), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n840), .A2(new_n746), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1139), .B1(new_n940), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1132), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n940), .B1(new_n842), .B2(new_n1138), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1130), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n835), .A2(new_n942), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n890), .A2(new_n746), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n665), .B(new_n1159), .C1(new_n729), .C2(new_n503), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1148), .A2(new_n1149), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT122), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1151), .A2(new_n1152), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1165), .A2(new_n1160), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT122), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n1149), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1137), .A2(new_n1144), .A3(new_n1166), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n714), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1146), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(G378));
  INV_X1    g0975(.A(KEYINPUT124), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n956), .A2(new_n960), .A3(G330), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n331), .A2(new_n690), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n330), .B2(new_n335), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n330), .A2(new_n335), .A3(new_n1180), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1185), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1177), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n956), .A3(G330), .A4(new_n960), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n945), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n931), .A3(new_n944), .A4(new_n1190), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1171), .A2(new_n1161), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1176), .B1(new_n1194), .B2(KEYINPUT57), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n715), .B1(new_n1194), .B2(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1171), .A2(new_n1161), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(KEYINPUT124), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1195), .A2(new_n1196), .A3(new_n1201), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n776), .A2(new_n506), .B1(new_n869), .B2(new_n785), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1060), .B(new_n1203), .C1(G97), .C2(new_n795), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n801), .A2(new_n973), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n783), .A2(G107), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n296), .A2(new_n305), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1207), .B(new_n986), .C1(G283), .C2(new_n770), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G50), .B1(new_n262), .B2(new_n305), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1209), .A2(new_n1210), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n801), .A2(G137), .B1(new_n783), .B2(G128), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n795), .A2(G132), .B1(new_n1092), .B2(G150), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n1111), .C2(new_n776), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n787), .A2(new_n1115), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT123), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n871), .A2(G159), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1212), .B1(new_n1210), .B2(new_n1209), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n765), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n757), .C1(G50), .C2(new_n845), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1188), .B2(new_n760), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1198), .B2(new_n756), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1202), .A2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n940), .A2(new_n760), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n757), .B1(G68), .B2(new_n845), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n869), .A2(new_n785), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n296), .B(new_n1233), .C1(G128), .C2(new_n770), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n782), .B2(new_n980), .C1(new_n268), .C2(new_n779), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1092), .A2(G50), .B1(new_n856), .B2(G159), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n867), .B2(new_n776), .C1(new_n854), .C2(new_n1115), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n390), .B(new_n985), .C1(G303), .C2(new_n770), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n782), .B2(new_n798), .C1(new_n554), .C2(new_n779), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1061), .B1(G294), .B2(new_n775), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n222), .B2(new_n787), .C1(new_n854), .C2(new_n506), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1235), .A2(new_n1237), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1232), .B1(new_n1242), .B2(new_n765), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1158), .A2(new_n756), .B1(new_n1231), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1162), .A2(new_n1027), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(G381));
  NOR2_X1   g1047(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1086), .A2(new_n1104), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n877), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1082), .A2(new_n827), .A3(new_n1084), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1251), .A2(G387), .A3(new_n1252), .A4(G381), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1253), .A2(new_n1174), .A3(new_n1229), .A4(new_n1202), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n691), .A2(G213), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1174), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G375), .C2(new_n1257), .ZN(G409));
  NAND2_X1  g1058(.A1(G393), .A2(G396), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1252), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G387), .A2(new_n1250), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1042), .B(new_n1043), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1026), .B1(new_n1106), .B2(new_n747), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n756), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G390), .B1(new_n1264), .B2(new_n1003), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1260), .B1(new_n1261), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G387), .A2(new_n1250), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1264), .A2(new_n1003), .A3(G390), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1252), .A4(new_n1259), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1172), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1202), .B(new_n1229), .C1(new_n1271), .C2(new_n1146), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1167), .A2(new_n1168), .A3(new_n1149), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1168), .B1(new_n1167), .B2(new_n1149), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1173), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1146), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1229), .B1(new_n1199), .B2(new_n1026), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1256), .B1(new_n1272), .B2(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1162), .A2(KEYINPUT60), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n715), .B1(new_n1280), .B2(new_n1246), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1246), .B2(new_n1280), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1244), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n877), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(G384), .A3(new_n1244), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT62), .B1(new_n1279), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT125), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1289), .B(new_n1256), .C1(new_n1272), .C2(new_n1278), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1278), .B1(G375), .B2(new_n1174), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT125), .B1(new_n1291), .B2(new_n1255), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1287), .A2(KEYINPUT62), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1288), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1256), .A2(G2897), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1286), .B(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1270), .B1(new_n1295), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1293), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1270), .A2(KEYINPUT61), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1279), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(new_n1286), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1297), .A2(new_n1305), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1302), .A2(new_n1303), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1301), .A2(new_n1308), .ZN(G405));
  NAND2_X1  g1109(.A1(G375), .A2(new_n1174), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(G375), .A2(new_n1174), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(KEYINPUT126), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1287), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1286), .B1(new_n1311), .B2(KEYINPUT126), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1310), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1310), .A3(new_n1314), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1316), .A2(new_n1269), .A3(new_n1266), .A4(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1317), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1270), .B1(new_n1319), .B2(new_n1315), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(G402));
endmodule


