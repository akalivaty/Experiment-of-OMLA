//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n456));
  NAND3_X1  g031(.A1(new_n456), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n457));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n456), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n459), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n458), .A2(G2105), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n467), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(G160));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n464), .A2(G2105), .A3(new_n457), .A4(new_n459), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI221_X1 g057(.A(new_n479), .B1(new_n480), .B2(new_n481), .C1(new_n465), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n480), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT69), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(new_n488), .C1(new_n480), .C2(new_n489), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n461), .A2(G138), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n464), .A2(new_n457), .A3(new_n459), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n460), .A2(new_n497), .A3(new_n464), .A4(new_n494), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n494), .A2(new_n500), .A3(new_n462), .A4(new_n459), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n491), .A2(new_n493), .B1(new_n499), .B2(new_n501), .ZN(G164));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n506), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT71), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n503), .B(new_n505), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n504), .B2(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n506), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(new_n513), .B1(new_n504), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(new_n503), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n503), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G651), .B1(G50), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n518), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n503), .A2(new_n529), .A3(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n531), .A2(G51), .B1(new_n514), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n510), .A2(G89), .A3(new_n516), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n534), .A2(KEYINPUT74), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(KEYINPUT74), .B1(new_n534), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g116(.A(KEYINPUT75), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n517), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n520), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(G52), .A2(new_n531), .B1(new_n547), .B2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n531), .A2(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n510), .A2(new_n516), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n554), .A2(KEYINPUT76), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(KEYINPUT76), .ZN(new_n556));
  OAI221_X1 g131(.A(new_n551), .B1(new_n552), .B2(new_n553), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT77), .Z(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g136(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n562));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n520), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n517), .A2(G91), .B1(G651), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n523), .A2(KEYINPUT9), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n523), .B2(new_n571), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n572), .A2(new_n570), .A3(new_n573), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n569), .B1(new_n574), .B2(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(new_n534), .A2(new_n536), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n534), .A2(KEYINPUT74), .A3(new_n536), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT75), .B1(new_n581), .B2(new_n533), .ZN(new_n582));
  INV_X1    g157(.A(new_n542), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(G286));
  NAND2_X1  g159(.A1(new_n517), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n524), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n517), .A2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n520), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n531), .A2(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n553), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT81), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G651), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(new_n602), .ZN(G290));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(G301), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n553), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n520), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(G54), .A2(new_n531), .B1(new_n613), .B2(G651), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT82), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n605), .B1(new_n616), .B2(new_n604), .ZN(G284));
  AOI21_X1  g192(.A(new_n605), .B1(new_n616), .B2(new_n604), .ZN(G321));
  NOR2_X1   g193(.A1(G299), .A2(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g195(.A(new_n619), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n557), .A2(new_n604), .ZN(new_n624));
  AND2_X1   g199(.A1(new_n616), .A2(new_n622), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g202(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n633));
  INV_X1    g208(.A(G123), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n480), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(G135), .B2(new_n466), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n631), .A2(new_n638), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(G14), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n651), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(G2100), .Z(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n637), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n671), .A2(new_n677), .A3(new_n675), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n677), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n680));
  AOI211_X1 g255(.A(new_n676), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1981), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT85), .B(KEYINPUT86), .Z(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(G32), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n466), .A2(G141), .ZN(new_n693));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT26), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n696), .A2(new_n697), .B1(G105), .B2(new_n473), .ZN(new_n698));
  INV_X1    g273(.A(G129), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n480), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT95), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n692), .B1(new_n703), .B2(G29), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G1996), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT96), .Z(new_n707));
  NAND2_X1  g282(.A1(G160), .A2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G34), .ZN(new_n709));
  AOI21_X1  g284(.A(G29), .B1(new_n709), .B2(KEYINPUT24), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(KEYINPUT24), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G2084), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n691), .A2(G26), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G116), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G2105), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT91), .ZN(new_n720));
  INV_X1    g295(.A(new_n480), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G128), .ZN(new_n722));
  INV_X1    g297(.A(G140), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n722), .C1(new_n723), .C2(new_n465), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n716), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G2067), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G5), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G171), .B2(new_n727), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(G1961), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(G1961), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n714), .A2(new_n726), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n704), .A2(new_n705), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n691), .A2(G35), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G162), .B2(new_n691), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT29), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G2090), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(G2090), .ZN(new_n738));
  NOR2_X1   g313(.A1(G164), .A2(new_n691), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G27), .B2(new_n691), .ZN(new_n740));
  INV_X1    g315(.A(G2078), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n733), .A2(new_n737), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G11), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT30), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n744), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n636), .B2(G29), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n752), .B1(new_n741), .B2(new_n740), .C1(new_n712), .C2(new_n713), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n707), .A2(new_n732), .A3(new_n743), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n727), .A2(G19), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n558), .B2(new_n727), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n727), .A2(G20), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT23), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G299), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G33), .ZN(new_n762));
  INV_X1    g337(.A(G139), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n465), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT92), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT25), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  INV_X1    g343(.A(G127), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n469), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n767), .B1(G2105), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT93), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n762), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT94), .B(G2072), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n761), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n757), .B(new_n776), .C1(new_n774), .C2(new_n775), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n754), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G16), .A2(G21), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G168), .B2(G16), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT97), .Z(new_n781));
  INV_X1    g356(.A(G1966), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n727), .A2(G4), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n616), .B2(new_n727), .ZN(new_n787));
  INV_X1    g362(.A(G1348), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n778), .A2(new_n783), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(KEYINPUT36), .ZN(new_n792));
  MUX2_X1   g367(.A(G23), .B(G288), .S(G16), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT89), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT33), .B(G1976), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G6), .B(G305), .S(G16), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT32), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G1981), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(G1981), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n727), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n727), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1971), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n796), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n727), .A2(G24), .ZN(new_n807));
  INV_X1    g382(.A(G290), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n727), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT88), .ZN(new_n810));
  INV_X1    g385(.A(G1986), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n691), .A2(G25), .ZN(new_n814));
  INV_X1    g389(.A(G131), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n465), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT87), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(G107), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G2105), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n721), .B2(G119), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n814), .B1(new_n823), .B2(new_n691), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT35), .B(G1991), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n791), .A2(KEYINPUT36), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n812), .A2(new_n813), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n792), .B1(new_n806), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n806), .A2(new_n792), .A3(new_n828), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n790), .B1(new_n830), .B2(new_n831), .ZN(G311));
  INV_X1    g407(.A(new_n790), .ZN(new_n833));
  INV_X1    g408(.A(new_n831), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n829), .ZN(G150));
  NAND2_X1  g410(.A1(new_n616), .A2(G559), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT99), .B(G55), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n531), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n510), .A2(G93), .A3(new_n516), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n520), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G651), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n838), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT100), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n838), .A2(new_n839), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n557), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n555), .A2(new_n556), .ZN(new_n849));
  INV_X1    g424(.A(new_n844), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n517), .A2(G81), .B1(G43), .B2(new_n531), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n846), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n836), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n844), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(G160), .B(new_n483), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT102), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n636), .ZN(new_n865));
  OR3_X1    g440(.A1(new_n461), .A2(KEYINPUT104), .A3(G118), .ZN(new_n866));
  OAI21_X1  g441(.A(KEYINPUT104), .B1(new_n461), .B2(G118), .ZN(new_n867));
  OR2_X1    g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n866), .A2(G2104), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G130), .ZN(new_n870));
  INV_X1    g445(.A(G142), .ZN(new_n871));
  OAI221_X1 g446(.A(new_n869), .B1(new_n480), .B2(new_n870), .C1(new_n465), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT105), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n629), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n823), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n701), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n773), .A2(KEYINPUT95), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(KEYINPUT103), .B2(new_n773), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n499), .A2(new_n501), .ZN(new_n879));
  INV_X1    g454(.A(new_n490), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n724), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n878), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n876), .A2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n865), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(new_n865), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n884), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g468(.A(G288), .B(G305), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n808), .A2(G303), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n599), .A2(G303), .A3(new_n602), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(G290), .A2(G166), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n897), .A3(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n848), .A2(new_n852), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n625), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n616), .A2(new_n622), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n853), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n615), .A2(G299), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n575), .A2(new_n574), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(new_n610), .A3(new_n569), .A4(new_n614), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n908), .B2(new_n910), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n908), .A2(KEYINPUT41), .A3(new_n910), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n904), .B(new_n906), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n913), .B1(new_n912), .B2(new_n916), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n902), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n915), .A2(new_n914), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n907), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n911), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n904), .B2(new_n906), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n902), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n917), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n604), .B1(new_n920), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n850), .A2(G868), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT106), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n918), .A2(new_n919), .A3(new_n902), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n926), .B1(new_n925), .B2(new_n917), .ZN(new_n932));
  OAI21_X1  g507(.A(G868), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n934));
  INV_X1    g509(.A(new_n929), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n935), .ZN(G331));
  AND3_X1   g513(.A1(new_n541), .A2(new_n542), .A3(G301), .ZN(new_n939));
  AOI21_X1  g514(.A(G301), .B1(new_n541), .B2(new_n542), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(new_n853), .ZN(new_n941));
  OAI21_X1  g516(.A(G171), .B1(new_n582), .B2(new_n583), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n541), .A2(new_n542), .A3(G301), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n903), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n921), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n853), .B1(new_n939), .B2(new_n940), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n903), .A3(new_n943), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n923), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n947), .A2(KEYINPUT108), .A3(new_n948), .A4(new_n923), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n953), .B(new_n921), .C1(new_n941), .C2(new_n944), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n946), .A2(new_n951), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n926), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n902), .A2(new_n945), .A3(new_n949), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n891), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT109), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n956), .A2(new_n963), .A3(new_n960), .A4(new_n957), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n902), .B1(new_n945), .B2(new_n949), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT43), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n956), .A2(KEYINPUT43), .A3(new_n960), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n959), .A2(new_n965), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(G397));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n490), .B1(new_n499), .B2(new_n501), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT110), .B(G1384), .Z(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n467), .A2(G40), .A3(new_n472), .A4(new_n475), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(G1996), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT112), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(new_n703), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n724), .B(G2067), .Z(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT113), .ZN(new_n987));
  INV_X1    g562(.A(new_n701), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n987), .B1(G1996), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(new_n982), .ZN(new_n990));
  INV_X1    g565(.A(new_n982), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n823), .B(new_n825), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n992), .B(KEYINPUT114), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n985), .B(new_n990), .C1(new_n991), .C2(new_n993), .ZN(new_n994));
  OR3_X1    g569(.A1(new_n808), .A2(KEYINPUT111), .A3(new_n811), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n808), .A2(new_n811), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT111), .B1(new_n808), .B2(new_n811), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n995), .B(new_n991), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n1001));
  NAND3_X1  g576(.A1(G286), .A2(new_n1001), .A3(G8), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT121), .B1(G168), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n975), .B1(new_n976), .B2(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT45), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1007), .B(new_n981), .C1(G164), .C2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1006), .B1(new_n1010), .B2(new_n782), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n981), .B1(G164), .B2(new_n1009), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT45), .B1(new_n881), .B2(new_n1008), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1006), .B(new_n782), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n976), .A2(G1384), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n980), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n713), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1005), .B1(new_n1011), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n1020), .B2(new_n1011), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1023), .A3(KEYINPUT51), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1022), .A2(new_n1025), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT122), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT62), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT122), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT62), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1015), .A2(new_n981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n585), .A2(new_n587), .A3(G1976), .A4(new_n588), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(G8), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1003), .B1(new_n1015), .B2(new_n981), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(KEYINPUT116), .A3(new_n1037), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1042), .A3(KEYINPUT52), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n1044));
  INV_X1    g619(.A(G1981), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n590), .A2(new_n1045), .A3(new_n594), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1045), .B1(new_n590), .B2(new_n594), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1048), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT49), .A3(new_n1046), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1051), .A3(new_n1041), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(new_n1041), .A3(new_n1037), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1043), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1043), .A2(KEYINPUT118), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT50), .B1(new_n976), .B2(G1384), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n981), .ZN(new_n1062));
  OR2_X1    g637(.A1(G164), .A2(G1384), .ZN(new_n1063));
  OAI22_X1  g638(.A1(new_n1062), .A2(KEYINPUT117), .B1(new_n1063), .B2(KEYINPUT50), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1062), .A2(KEYINPUT117), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1064), .A2(new_n1065), .A3(G2090), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n975), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n976), .A2(new_n977), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n980), .B1(new_n1068), .B2(KEYINPUT45), .ZN(new_n1069));
  AOI21_X1  g644(.A(G1971), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G303), .A2(G8), .ZN(new_n1072));
  NOR2_X1   g647(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(G2090), .ZN(new_n1079));
  OAI21_X1  g654(.A(G8), .B1(new_n1079), .B2(new_n1070), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(new_n1076), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1060), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1010), .A2(new_n1083), .A3(G2078), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1961), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1086));
  OR3_X1    g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1083), .B1(new_n1090), .B2(G2078), .ZN(new_n1091));
  AOI21_X1  g666(.A(G301), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1082), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1030), .A2(new_n1035), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1041), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G288), .A2(G1976), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1047), .B1(new_n1052), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1081), .A2(new_n1056), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(G8), .B(G168), .C1(new_n1020), .C2(new_n1011), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1060), .A2(new_n1077), .A3(new_n1081), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1056), .B1(new_n1080), .B2(new_n1076), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1104), .A2(KEYINPUT63), .A3(new_n1081), .A4(new_n1100), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1098), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n572), .B2(new_n573), .ZN(new_n1107));
  AOI22_X1  g682(.A1(G299), .A2(KEYINPUT57), .B1(new_n569), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1067), .A2(new_n1069), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1108), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1036), .A2(G2067), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1078), .B2(new_n788), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n615), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1113), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n615), .ZN(new_n1119));
  AOI211_X1 g694(.A(new_n1119), .B(new_n1115), .C1(new_n1078), .C2(new_n788), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT60), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1116), .A2(new_n1122), .A3(new_n1119), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1036), .A2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT120), .B(G1996), .Z(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1090), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n558), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1127), .B2(new_n558), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1121), .B(new_n1123), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1114), .A2(KEYINPUT61), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(new_n1113), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1118), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1069), .A2(KEYINPUT53), .A3(new_n741), .A4(new_n978), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT124), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1086), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1091), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(G171), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1136), .B1(new_n1092), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1114), .A2(KEYINPUT61), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1136), .B1(new_n1140), .B2(G171), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1089), .A2(G301), .A3(new_n1091), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(new_n1146), .A3(new_n1082), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1106), .B1(new_n1135), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1000), .B1(new_n1094), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n997), .A2(new_n991), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT126), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n994), .ZN(new_n1154));
  INV_X1    g729(.A(new_n823), .ZN(new_n1155));
  NOR4_X1   g730(.A1(new_n990), .A2(new_n985), .A3(new_n825), .A4(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n724), .A2(G2067), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n991), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n991), .B1(new_n987), .B2(new_n988), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT47), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1154), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1149), .A2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g740(.A(G227), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1167), .A2(G319), .ZN(new_n1168));
  XNOR2_X1  g742(.A(new_n1168), .B(KEYINPUT127), .ZN(new_n1169));
  NOR3_X1   g743(.A1(G229), .A2(G401), .A3(new_n1169), .ZN(new_n1170));
  AND3_X1   g744(.A1(new_n967), .A2(new_n892), .A3(new_n1170), .ZN(G308));
  NAND3_X1  g745(.A1(new_n967), .A2(new_n892), .A3(new_n1170), .ZN(G225));
endmodule


