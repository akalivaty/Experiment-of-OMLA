//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n206), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n216), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT66), .B(G244), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G77), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G97), .A2(G257), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n210), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n225), .B1(KEYINPUT1), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  INV_X1    g0050(.A(G50), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n201), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n249), .B(new_n253), .ZN(G351));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G222), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n255), .B(new_n257), .C1(new_n258), .C2(new_n256), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n259), .B(new_n262), .C1(G77), .C2(new_n255), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  AND2_X1   g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  OAI21_X1  g0065(.A(G274), .B1(new_n265), .B2(new_n219), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n264), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n268), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n270), .A2(new_n261), .A3(KEYINPUT69), .A4(G274), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n261), .A2(new_n268), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n275), .A2(G226), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(G226), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n263), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G190), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(G200), .B2(new_n279), .ZN(new_n282));
  OAI21_X1  g0082(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT71), .A2(G58), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT8), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n220), .A3(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n283), .B(new_n286), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n219), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT72), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT72), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n295), .A2(new_n267), .A3(G13), .A4(G20), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n290), .A2(new_n292), .B1(new_n251), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n292), .B1(new_n294), .B2(new_n296), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n267), .A2(G20), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(KEYINPUT9), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n298), .B2(new_n302), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n282), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT10), .B1(new_n282), .B2(KEYINPUT74), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n282), .B1(KEYINPUT74), .B2(KEYINPUT10), .C1(new_n304), .C2(new_n306), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n279), .A2(G179), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n279), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n303), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n309), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT76), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n317));
  INV_X1    g0117(.A(G77), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n220), .A2(G33), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT11), .A3(new_n292), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT11), .B1(new_n320), .B2(new_n292), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n316), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n292), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT11), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(KEYINPUT76), .A3(new_n321), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT12), .ZN(new_n329));
  OAI21_X1  g0129(.A(G68), .B1(new_n301), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n294), .A2(new_n296), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n331), .A2(new_n329), .A3(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n329), .B2(new_n331), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n324), .A2(new_n328), .A3(new_n330), .A4(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT77), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n272), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n269), .A2(KEYINPUT75), .A3(new_n271), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G97), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n240), .A2(G1698), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G226), .B2(G1698), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n339), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(new_n262), .B1(new_n274), .B2(G238), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n337), .A2(new_n338), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT13), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT13), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n337), .A2(new_n346), .A3(new_n349), .A4(new_n338), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT14), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(G169), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(G179), .A3(new_n350), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n352), .B1(new_n351), .B2(G169), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n335), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n334), .B1(new_n351), .B2(G200), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n348), .A2(G190), .A3(new_n350), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G238), .A2(G1698), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n255), .B(new_n361), .C1(new_n240), .C2(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n262), .C1(G107), .C2(new_n255), .ZN(new_n363));
  INV_X1    g0163(.A(new_n226), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n273), .ZN(new_n365));
  INV_X1    g0165(.A(new_n272), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g0169(.A(KEYINPUT8), .B(G58), .Z(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n372), .B(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n371), .B1(new_n374), .B2(new_n319), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n292), .B1(new_n318), .B2(new_n297), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n301), .A2(G77), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n312), .B1(new_n365), .B2(new_n366), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n369), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n367), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(G190), .B2(new_n367), .ZN(new_n384));
  INV_X1    g0184(.A(new_n378), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n315), .A2(new_n357), .A3(new_n360), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT82), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT81), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n258), .A2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(KEYINPUT79), .C1(new_n343), .C2(new_n342), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT79), .B1(new_n255), .B2(new_n390), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(G226), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n261), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT80), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n273), .B2(new_n240), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n261), .A2(new_n268), .A3(KEYINPUT80), .A4(G232), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n272), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n389), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n390), .B1(new_n342), .B2(new_n343), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT79), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(new_n396), .A3(new_n395), .A4(new_n391), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n262), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n400), .A2(new_n401), .B1(new_n269), .B2(new_n271), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT81), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n404), .A2(new_n382), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(G190), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G58), .A2(G68), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n203), .A2(new_n205), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n288), .A2(G159), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT7), .B1(new_n344), .B2(new_n220), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT7), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n342), .A2(new_n343), .A3(new_n424), .A4(G20), .ZN(new_n425));
  OAI21_X1  g0225(.A(G68), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT78), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n419), .A2(new_n427), .A3(new_n420), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n422), .A2(KEYINPUT16), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT16), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n424), .B1(new_n255), .B2(G20), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n344), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n202), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n430), .B1(new_n433), .B2(new_n421), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n434), .A3(new_n292), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n331), .A2(new_n285), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n301), .B2(new_n285), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n416), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n416), .B2(new_n438), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n388), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT81), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT81), .B1(new_n409), .B2(new_n410), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n414), .B1(new_n445), .B2(new_n382), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n435), .A2(new_n437), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT17), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n416), .A2(new_n438), .A3(new_n439), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(KEYINPUT82), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT18), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n413), .A2(G179), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n445), .B2(new_n312), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n453), .B2(new_n447), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n404), .A2(new_n312), .A3(new_n411), .ZN(new_n455));
  INV_X1    g0255(.A(new_n452), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n451), .A2(new_n447), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n442), .A2(new_n450), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n387), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G303), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n344), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G264), .A2(G1698), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n213), .B2(G1698), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n462), .B(new_n262), .C1(new_n344), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G41), .ZN(new_n467));
  INV_X1    g0267(.A(G41), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n267), .B(G45), .C1(new_n468), .C2(KEYINPUT5), .ZN(new_n469));
  OR3_X1    g0269(.A1(new_n266), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G270), .B(new_n261), .C1(new_n469), .C2(new_n467), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n465), .A2(new_n470), .A3(G179), .A4(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n291), .A2(new_n219), .B1(G20), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n220), .C1(G33), .C2(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n474), .A2(KEYINPUT20), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT20), .B1(new_n474), .B2(new_n477), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n478), .A2(new_n479), .B1(G116), .B2(new_n331), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n267), .A2(G33), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n299), .A2(G116), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT87), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n473), .A2(G20), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n477), .A2(new_n292), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT20), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n474), .A2(KEYINPUT20), .A3(new_n477), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n487), .A2(new_n488), .B1(new_n297), .B2(new_n473), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT87), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n299), .A2(G116), .A3(new_n481), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n472), .B1(new_n483), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n465), .A2(new_n470), .A3(new_n471), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G169), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n480), .A2(new_n482), .A3(KEYINPUT87), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n490), .B1(new_n489), .B2(new_n491), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT21), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n493), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n495), .B1(new_n483), .B2(new_n492), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT21), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n465), .A2(new_n471), .A3(new_n470), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G190), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n494), .A2(G200), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n483), .A3(new_n492), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n501), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  OAI211_X1 g0310(.A(G257), .B(new_n261), .C1(new_n469), .C2(new_n467), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n470), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(G250), .B1(new_n342), .B2(new_n343), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G1698), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  INV_X1    g0316(.A(G244), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n344), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n516), .A2(G1698), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(G244), .C1(new_n343), .C2(new_n342), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n515), .A2(new_n475), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n512), .B1(new_n521), .B2(new_n262), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n510), .B1(new_n522), .B2(new_n382), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT84), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n476), .B1(new_n299), .B2(new_n481), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n331), .A2(new_n476), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n292), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n331), .A2(new_n529), .A3(new_n481), .ZN(new_n530));
  OAI211_X1 g0330(.A(KEYINPUT84), .B(new_n526), .C1(new_n530), .C2(new_n476), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT83), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n289), .A2(new_n318), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g0334(.A(G97), .B(G107), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT6), .ZN(new_n536));
  INV_X1    g0336(.A(G107), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n476), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n532), .B(new_n534), .C1(new_n539), .C2(new_n220), .ZN(new_n540));
  AND2_X1   g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n220), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT83), .B1(new_n545), .B2(new_n533), .ZN(new_n546));
  OAI21_X1  g0346(.A(G107), .B1(new_n423), .B2(new_n425), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n528), .A2(new_n531), .B1(new_n548), .B2(new_n292), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n518), .A2(new_n475), .A3(new_n520), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n256), .B1(new_n513), .B2(KEYINPUT4), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n262), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n470), .A2(new_n511), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(G190), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(KEYINPUT85), .A3(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n523), .A2(new_n549), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G257), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G294), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n513), .C2(G1698), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n262), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n261), .B1(new_n469), .B2(new_n467), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G264), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n470), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n382), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(G190), .B2(new_n565), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n220), .B2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n537), .A2(KEYINPUT23), .A3(G20), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n220), .A2(G33), .A3(G116), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G87), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n574), .A2(G20), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n342), .B2(new_n343), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT22), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT89), .B1(new_n577), .B2(KEYINPUT88), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT88), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT89), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT22), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n255), .A2(new_n575), .B1(new_n578), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n573), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT90), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n573), .B(KEYINPUT90), .C1(new_n583), .C2(new_n584), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n576), .A2(new_n582), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n255), .A2(new_n578), .A3(new_n581), .A4(new_n575), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT90), .B1(new_n593), .B2(new_n573), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n292), .B(new_n588), .C1(new_n590), .C2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n331), .A2(G107), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n596), .A2(KEYINPUT25), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(KEYINPUT25), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n530), .B2(G107), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n567), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n531), .A2(new_n528), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n548), .A2(new_n292), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(G169), .B1(new_n552), .B2(new_n553), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n522), .A2(new_n368), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G45), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n209), .B1(new_n608), .B2(G1), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n267), .A2(G45), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n261), .B(new_n609), .C1(G274), .C2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n610), .A2(G274), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n614), .A2(KEYINPUT86), .A3(new_n261), .A4(new_n609), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n517), .A2(G1698), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(G238), .B2(G1698), .ZN(new_n618));
  INV_X1    g0418(.A(G33), .ZN(new_n619));
  OAI22_X1  g0419(.A1(new_n618), .A2(new_n344), .B1(new_n619), .B2(new_n473), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n262), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n616), .A2(new_n368), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(G169), .B1(new_n616), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n372), .A2(new_n373), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n372), .A2(new_n373), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n297), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT19), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n220), .B1(new_n339), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n574), .A2(new_n476), .A3(new_n537), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n220), .B(G68), .C1(new_n342), .C2(new_n343), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n628), .B1(new_n319), .B2(new_n476), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n292), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n299), .A2(new_n481), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n627), .B(new_n635), .C1(new_n636), .C2(new_n374), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n382), .B1(new_n616), .B2(new_n621), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n299), .A2(G87), .A3(new_n481), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n627), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n613), .A2(new_n615), .B1(new_n620), .B2(new_n262), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G190), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n624), .A2(new_n637), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n557), .A2(new_n600), .A3(new_n607), .A4(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n595), .A2(new_n599), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT91), .B1(new_n565), .B2(new_n368), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n560), .A2(new_n262), .B1(new_n563), .B2(G264), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(G179), .A4(new_n470), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n565), .A2(G169), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n460), .A2(new_n509), .A3(new_n646), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT92), .ZN(G372));
  INV_X1    g0456(.A(new_n314), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n351), .A2(G169), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n354), .A3(new_n353), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n335), .B1(new_n360), .B2(new_n381), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT94), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n450), .B(new_n442), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n458), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n309), .A2(new_n310), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n657), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n501), .A2(new_n654), .A3(new_n503), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT93), .B1(new_n668), .B2(new_n645), .ZN(new_n669));
  INV_X1    g0469(.A(new_n638), .ZN(new_n670));
  INV_X1    g0470(.A(new_n640), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n643), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n642), .A2(new_n368), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n637), .C1(G169), .C2(new_n642), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n607), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n604), .B1(new_n368), .B2(new_n522), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n644), .A2(new_n677), .A3(new_n603), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n679), .A3(new_n674), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n501), .A2(new_n654), .A3(new_n503), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT85), .B1(new_n555), .B2(G200), .ZN(new_n683));
  AOI211_X1 g0483(.A(new_n510), .B(new_n382), .C1(new_n552), .C2(new_n553), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n601), .A2(new_n602), .A3(new_n554), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n678), .B2(new_n603), .ZN(new_n687));
  INV_X1    g0487(.A(new_n647), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n675), .B1(new_n688), .B2(new_n567), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n682), .A2(new_n687), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n669), .A2(new_n681), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n460), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n667), .A2(new_n693), .ZN(G369));
  NAND2_X1  g0494(.A1(new_n501), .A2(new_n503), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n267), .A2(new_n220), .A3(G13), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G213), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n497), .B2(new_n498), .ZN(new_n702));
  MUX2_X1   g0502(.A(new_n695), .B(new_n509), .S(new_n702), .Z(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n701), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n654), .B(new_n600), .C1(new_n688), .C2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n654), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n701), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n704), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n695), .A2(new_n705), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n706), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n654), .A2(new_n701), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(G399));
  NOR2_X1   g0515(.A1(new_n212), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n630), .A2(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n217), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n646), .A2(new_n509), .A3(new_n654), .A4(new_n705), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  INV_X1    g0524(.A(new_n472), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n642), .A3(new_n649), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n724), .B1(new_n726), .B2(new_n555), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n504), .A2(G179), .A3(new_n642), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n555), .A3(new_n565), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n649), .A2(new_n642), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n522), .A3(KEYINPUT30), .A4(new_n725), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT31), .B1(new_n732), .B2(new_n701), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n722), .B1(new_n723), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n692), .A2(new_n705), .ZN(new_n737));
  XNOR2_X1  g0537(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n682), .A2(new_n687), .A3(new_n672), .A4(new_n600), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n701), .B1(new_n681), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n736), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n721), .B1(new_n743), .B2(G1), .ZN(G364));
  AND2_X1   g0544(.A1(new_n220), .A2(G13), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G45), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n717), .A2(G1), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n368), .A2(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n220), .A2(G190), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n382), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G77), .A2(new_n752), .B1(new_n755), .B2(G107), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n220), .A2(new_n280), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n749), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n756), .B1(new_n201), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n220), .B1(new_n760), .B2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n476), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n757), .A2(new_n753), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n255), .B1(new_n763), .B2(new_n574), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n759), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n750), .A2(new_n760), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G159), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NAND3_X1  g0569(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n280), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n772), .A2(new_n202), .B1(new_n774), .B2(new_n251), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n763), .A2(new_n461), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n754), .B1(new_n751), .B2(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n777), .B(new_n780), .C1(G329), .C2(new_n767), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n344), .B1(new_n758), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  INV_X1    g0584(.A(G294), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n772), .A2(new_n784), .B1(new_n785), .B2(new_n761), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n783), .B(new_n786), .C1(G326), .C2(new_n773), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n765), .A2(new_n776), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n219), .B1(G20), .B2(new_n312), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n748), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n253), .A2(G45), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT97), .Z(new_n793));
  NOR2_X1   g0593(.A1(new_n212), .A2(new_n255), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(G45), .C2(new_n217), .ZN(new_n795));
  INV_X1    g0595(.A(G355), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n255), .A2(new_n211), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT96), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n795), .B1(G116), .B2(new_n211), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n789), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n791), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n802), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n703), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n748), .B1(new_n703), .B2(G330), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(G330), .B2(new_n703), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NOR2_X1   g0610(.A1(new_n380), .A2(new_n701), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n385), .A2(new_n705), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n384), .B2(new_n385), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n814), .B2(new_n381), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n737), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n367), .A2(G190), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n385), .B(new_n817), .C1(new_n382), .C2(new_n367), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n385), .B2(new_n705), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n811), .B1(new_n819), .B2(new_n380), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n692), .A2(new_n705), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n736), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n748), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  INV_X1    g0625(.A(new_n758), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G143), .A2(new_n826), .B1(new_n752), .B2(G159), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n774), .B2(new_n828), .C1(new_n287), .C2(new_n772), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT34), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n255), .B1(new_n754), .B2(new_n202), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n763), .A2(new_n251), .B1(new_n766), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n761), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n832), .B(new_n834), .C1(G58), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n830), .B2(new_n829), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n754), .A2(new_n574), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n758), .A2(new_n785), .B1(new_n751), .B2(new_n473), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n839), .B(new_n840), .C1(G311), .C2(new_n767), .ZN(new_n841));
  INV_X1    g0641(.A(new_n762), .ZN(new_n842));
  INV_X1    g0642(.A(new_n763), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n255), .B1(new_n843), .B2(G107), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n771), .A2(G283), .B1(new_n773), .B2(G303), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n841), .A2(new_n842), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT98), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n789), .B1(new_n838), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n789), .A2(new_n800), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n747), .B1(new_n318), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n848), .B(new_n850), .C1(new_n820), .C2(new_n801), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n825), .A2(new_n851), .ZN(G384));
  NOR2_X1   g0652(.A1(new_n745), .A2(new_n267), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n739), .A2(new_n460), .A3(new_n742), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n667), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT99), .ZN(new_n856));
  INV_X1    g0656(.A(new_n699), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n458), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n433), .B1(KEYINPUT78), .B2(new_n421), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT16), .B1(new_n861), .B2(new_n428), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n429), .A2(new_n292), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n437), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n453), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n416), .A2(new_n438), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n857), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n453), .A2(new_n447), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n447), .A2(new_n857), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n870), .A2(new_n866), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n867), .ZN(new_n874));
  AOI221_X4 g0674(.A(new_n860), .B1(new_n869), .B2(new_n873), .C1(new_n459), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n459), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n869), .A2(new_n873), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n821), .A2(new_n812), .ZN(new_n880));
  INV_X1    g0680(.A(new_n360), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n335), .B(new_n701), .C1(new_n660), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n335), .A2(new_n701), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n357), .A2(new_n360), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n859), .B1(new_n879), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n660), .A2(new_n335), .A3(new_n705), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n876), .A2(new_n877), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n860), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n870), .A2(new_n866), .A3(new_n872), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(new_n871), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n448), .A2(new_n449), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n872), .B1(new_n458), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n860), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n894), .A2(new_n900), .A3(new_n891), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n890), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n888), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n856), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n723), .A2(new_n735), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n885), .A2(new_n906), .A3(KEYINPUT40), .A4(new_n820), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n894), .B2(new_n900), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n815), .B1(new_n882), .B2(new_n884), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n906), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n875), .B2(new_n878), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n460), .A2(new_n906), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n722), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n914), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n853), .B1(new_n905), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n905), .B2(new_n917), .ZN(new_n919));
  INV_X1    g0719(.A(new_n539), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT35), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(KEYINPUT35), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(G116), .A4(new_n221), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT36), .Z(new_n924));
  NAND3_X1  g0724(.A1(new_n218), .A2(G77), .A3(new_n417), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n251), .A2(G68), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n267), .B(G13), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n919), .A2(new_n928), .ZN(G367));
  INV_X1    g0729(.A(new_n803), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n244), .B2(new_n794), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n211), .B2(new_n374), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n748), .ZN(new_n933));
  AOI22_X1  g0733(.A1(G77), .A2(new_n755), .B1(new_n767), .B2(G137), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n934), .B1(new_n251), .B2(new_n751), .C1(new_n201), .C2(new_n763), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n761), .A2(new_n202), .ZN(new_n936));
  INV_X1    g0736(.A(G159), .ZN(new_n937));
  INV_X1    g0737(.A(G143), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n772), .A2(new_n937), .B1(new_n774), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n255), .B1(new_n758), .B2(new_n287), .ZN(new_n940));
  NOR4_X1   g0740(.A1(new_n935), .A2(new_n936), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n763), .A2(new_n473), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n942), .A2(KEYINPUT46), .B1(G311), .B2(new_n773), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n943), .B1(KEYINPUT46), .B2(new_n942), .C1(new_n537), .C2(new_n761), .ZN(new_n944));
  AOI22_X1  g0744(.A1(G303), .A2(new_n826), .B1(new_n752), .B2(G283), .ZN(new_n945));
  INV_X1    g0745(.A(G317), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n946), .B2(new_n766), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n344), .B1(new_n754), .B2(new_n476), .C1(new_n772), .C2(new_n785), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  AOI21_X1  g0751(.A(new_n933), .B1(new_n951), .B2(new_n789), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n671), .A2(new_n705), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n624), .A3(new_n637), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n675), .B2(new_n953), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(new_n805), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n746), .A2(G1), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT103), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT45), .ZN(new_n960));
  INV_X1    g0760(.A(new_n714), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n678), .A2(new_n603), .A3(new_n701), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT100), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n687), .B1(new_n549), .B2(new_n705), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n960), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n714), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n714), .A2(KEYINPUT44), .A3(new_n965), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT44), .B1(new_n714), .B2(new_n965), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n709), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n710), .A2(new_n969), .A3(new_n972), .A4(new_n971), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n743), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT102), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n711), .A2(new_n706), .A3(new_n708), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n712), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n711), .A2(new_n706), .A3(new_n708), .A4(KEYINPUT102), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(new_n704), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n959), .B1(new_n976), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n974), .A2(new_n975), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n987), .A2(new_n984), .A3(KEYINPUT103), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n743), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n716), .B(KEYINPUT41), .Z(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n958), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n955), .B(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n965), .A2(new_n712), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT42), .Z(new_n995));
  OAI21_X1  g0795(.A(new_n607), .B1(new_n966), .B2(new_n654), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n705), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n993), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT101), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT101), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n995), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n710), .A2(new_n966), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n957), .B1(new_n992), .B2(new_n1006), .ZN(G387));
  OAI22_X1  g0807(.A1(new_n763), .A2(new_n785), .B1(new_n761), .B2(new_n778), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G317), .A2(new_n826), .B1(new_n752), .B2(G303), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n774), .B2(new_n782), .C1(new_n779), .C2(new_n772), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n255), .B1(new_n767), .B2(G326), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n473), .B2(new_n754), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT105), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1015), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n374), .A2(new_n761), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n773), .A2(G159), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n255), .B1(new_n754), .B2(new_n476), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n285), .B2(new_n771), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n763), .A2(new_n318), .B1(new_n751), .B2(new_n202), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n758), .A2(new_n251), .B1(new_n766), .B2(new_n287), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n790), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n798), .A2(new_n718), .B1(G107), .B2(new_n211), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n241), .A2(G45), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n370), .A2(new_n251), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(KEYINPUT104), .B(KEYINPUT50), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n718), .B(new_n608), .C1(new_n202), .C2(new_n318), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n212), .B(new_n255), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1030), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n748), .B1(new_n1038), .B2(new_n930), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1029), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n708), .A2(new_n706), .A3(new_n802), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n958), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n977), .A2(KEYINPUT106), .A3(new_n983), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n984), .A2(new_n716), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT106), .B1(new_n977), .B2(new_n983), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1042), .B1(new_n1043), .B2(new_n983), .C1(new_n1045), .C2(new_n1046), .ZN(G393));
  AOI21_X1  g0847(.A(new_n717), .B1(new_n987), .B2(new_n984), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n986), .B2(new_n988), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n803), .B1(new_n476), .B2(new_n211), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n248), .B2(new_n794), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n826), .A2(G159), .B1(G150), .B2(new_n773), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n763), .A2(new_n202), .B1(new_n766), .B2(new_n938), .ZN(new_n1054));
  OR4_X1    g0854(.A1(new_n344), .A2(new_n1053), .A3(new_n839), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n370), .A2(new_n752), .B1(new_n835), .B2(G77), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n251), .B2(new_n772), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT107), .Z(new_n1058));
  AOI22_X1  g0858(.A1(new_n835), .A2(G116), .B1(G303), .B2(new_n771), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1059), .A2(KEYINPUT108), .B1(G294), .B2(new_n752), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(KEYINPUT108), .B2(new_n1059), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT109), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n774), .A2(new_n946), .B1(new_n758), .B2(new_n779), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n255), .B1(new_n755), .B2(G107), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G283), .A2(new_n843), .B1(new_n767), .B2(G322), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1055), .A2(new_n1058), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n747), .B(new_n1051), .C1(new_n1068), .C2(new_n789), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n965), .B2(new_n805), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n987), .B2(new_n1043), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(KEYINPUT110), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT110), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1073), .B(new_n1070), .C1(new_n987), .C2(new_n1043), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1049), .A2(new_n1075), .ZN(G390));
  NOR4_X1   g0876(.A1(new_n645), .A2(new_n508), .A3(new_n707), .A4(new_n701), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n734), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(G330), .B(new_n820), .C1(new_n1077), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n885), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1081), .A2(new_n1082), .B1(new_n909), .B2(new_n736), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n682), .A2(new_n687), .A3(new_n689), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n680), .B1(new_n1084), .B2(KEYINPUT93), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n701), .B1(new_n1085), .B2(new_n691), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n811), .B1(new_n1086), .B2(new_n820), .ZN(new_n1087));
  OAI21_X1  g0887(.A(KEYINPUT111), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT111), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n909), .A2(new_n736), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n885), .B1(new_n736), .B2(new_n820), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n880), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n819), .A2(new_n380), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n811), .B1(new_n741), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1088), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n460), .A2(new_n736), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n667), .A2(new_n854), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n889), .B1(new_n1087), .B2(new_n1082), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT39), .B1(new_n875), .B2(new_n878), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n901), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n894), .A2(new_n900), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1104), .B(new_n889), .C1(new_n1082), .C2(new_n1094), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1090), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1090), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1103), .A2(new_n1108), .A3(new_n1105), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1100), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1099), .B(KEYINPUT112), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1103), .A2(new_n1108), .A3(new_n1105), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1108), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n716), .B(new_n1110), .C1(new_n1111), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n958), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1102), .A2(new_n800), .A3(new_n901), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n849), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n748), .B1(new_n285), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n774), .A2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n344), .B(new_n1121), .C1(G125), .C2(new_n767), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT54), .B(G143), .Z(new_n1123));
  AOI22_X1  g0923(.A1(new_n752), .A2(new_n1123), .B1(new_n755), .B2(G50), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(new_n833), .C2(new_n758), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n763), .A2(new_n287), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n828), .B2(new_n772), .C1(new_n937), .C2(new_n761), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n344), .B1(new_n763), .B2(new_n574), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT115), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n754), .A2(new_n202), .B1(new_n766), .B2(new_n785), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G116), .B2(new_n826), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n835), .A2(G77), .B1(G283), .B2(new_n773), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n772), .A2(new_n537), .B1(new_n751), .B2(new_n476), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT114), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1125), .A2(new_n1129), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1119), .B1(new_n1138), .B2(new_n789), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT116), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1117), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1115), .A2(new_n1116), .A3(new_n1141), .ZN(G378));
  INV_X1    g0942(.A(KEYINPUT121), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1104), .A2(KEYINPUT40), .A3(new_n911), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n910), .B1(new_n893), .B2(new_n894), .ZN(new_n1145));
  OAI211_X1 g0945(.A(G330), .B(new_n1144), .C1(new_n1145), .C2(KEYINPUT40), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n888), .A3(new_n903), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n889), .B1(new_n1102), .B2(new_n901), .ZN(new_n1148));
  OAI211_X1 g0948(.A(G330), .B(new_n914), .C1(new_n1148), .C2(new_n887), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n303), .A2(new_n857), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT55), .Z(new_n1151));
  XNOR2_X1  g0951(.A(new_n315), .B(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(KEYINPUT120), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1147), .A2(new_n1149), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1143), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1158), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1147), .A2(new_n1149), .A3(new_n1158), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1164), .A2(KEYINPUT121), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT122), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1112), .A2(new_n1113), .A3(new_n1099), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1098), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1110), .A2(KEYINPUT122), .A3(new_n1098), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT57), .B1(new_n1167), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT57), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1169), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT122), .B1(new_n1110), .B2(new_n1098), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n716), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1174), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n255), .A2(G41), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G50), .B(new_n1182), .C1(new_n619), .C2(new_n468), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n754), .A2(new_n201), .B1(new_n766), .B2(new_n778), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n318), .B2(new_n763), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT117), .B1(new_n758), .B2(new_n537), .ZN(new_n1186));
  OR3_X1    g0986(.A1(new_n758), .A2(KEYINPUT117), .A3(new_n537), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1184), .B(new_n1185), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n774), .A2(new_n473), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n936), .B(new_n1189), .C1(G97), .C2(new_n771), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(new_n374), .C2(new_n751), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1183), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n843), .A2(new_n1123), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT118), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n758), .A2(new_n1120), .B1(new_n751), .B2(new_n828), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G132), .B2(new_n771), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n835), .A2(G150), .B1(G125), .B2(new_n773), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n755), .A2(G159), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1193), .B1(new_n1192), .B2(new_n1191), .C1(new_n1200), .C2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n789), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n747), .B1(new_n251), .B2(new_n849), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n1157), .C2(new_n801), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1167), .B2(new_n958), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1181), .A2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n1082), .A2(new_n800), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n255), .B1(new_n754), .B2(new_n201), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT123), .Z(new_n1214));
  AOI22_X1  g1014(.A1(G150), .A2(new_n752), .B1(new_n767), .B2(G128), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G137), .A2(new_n826), .B1(new_n843), .B2(G159), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n774), .A2(new_n833), .B1(new_n761), .B2(new_n251), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n771), .B2(new_n1123), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n344), .B1(new_n754), .B2(new_n318), .C1(new_n774), .C2(new_n785), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G116), .B2(new_n771), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G107), .A2(new_n752), .B1(new_n767), .B2(G303), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G97), .A2(new_n843), .B1(new_n826), .B2(G283), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1221), .A2(new_n1021), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n790), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n747), .B(new_n1225), .C1(new_n202), .C2(new_n849), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1096), .A2(new_n958), .B1(new_n1212), .B2(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n991), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1227), .B1(new_n1111), .B2(new_n1229), .ZN(G381));
  NAND3_X1  g1030(.A1(new_n976), .A2(new_n959), .A3(new_n985), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT103), .B1(new_n987), .B2(new_n984), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n977), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1043), .B1(new_n1233), .B2(new_n990), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1005), .ZN(new_n1235));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n957), .A3(new_n1236), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1238));
  OR4_X1    g1038(.A1(G378), .A2(G375), .A3(new_n1237), .A4(new_n1238), .ZN(G407));
  INV_X1    g1039(.A(G378), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n700), .A2(G213), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT124), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G407), .B(G213), .C1(G375), .C2(new_n1243), .ZN(G409));
  XNOR2_X1  g1044(.A(G393), .B(new_n809), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1235), .A2(new_n957), .A3(new_n1236), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1236), .B1(new_n1235), .B2(new_n957), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G387), .A2(G390), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1245), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1237), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G378), .B(new_n1210), .C1(new_n1174), .C2(new_n1180), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1167), .A2(new_n991), .A3(new_n1173), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1209), .B1(new_n1255), .B2(new_n958), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1240), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1242), .B1(new_n1253), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1228), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1228), .A2(new_n1260), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1261), .A2(new_n716), .A3(new_n1099), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1227), .ZN(new_n1264));
  INV_X1    g1064(.A(G384), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(G384), .A3(new_n1227), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1259), .A2(KEYINPUT127), .A3(new_n1270), .ZN(new_n1271));
  XOR2_X1   g1071(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1272));
  INV_X1    g1072(.A(new_n1241), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1253), .B2(new_n1258), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1274), .B2(new_n1269), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT127), .B1(new_n1259), .B2(new_n1270), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1271), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1242), .A2(G2897), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1268), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(G2897), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1268), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1278), .B1(new_n1283), .B2(new_n1259), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1252), .B1(new_n1277), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1248), .A2(new_n1278), .A3(new_n1251), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1253), .A2(new_n1258), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1242), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1268), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1287), .B(new_n1292), .C1(new_n1274), .C2(new_n1283), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT63), .B1(new_n1274), .B2(new_n1269), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1286), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1248), .A2(new_n1278), .A3(new_n1251), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1288), .A2(new_n1241), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1282), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1290), .B1(new_n1297), .B2(new_n1268), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(KEYINPUT125), .A4(new_n1292), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1295), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1285), .A2(new_n1301), .ZN(G405));
  AOI21_X1  g1102(.A(G378), .B1(new_n1181), .B2(new_n1210), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1253), .ZN(new_n1304));
  OR3_X1    g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1269), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1269), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1252), .ZN(G402));
endmodule


