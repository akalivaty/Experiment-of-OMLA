//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT65), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n212), .B1(KEYINPUT1), .B2(new_n224), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n225), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(new_n206), .B2(G20), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G50), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n249), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G58), .ZN(new_n257));
  OR3_X1    g0057(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT8), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n207), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n253), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n251), .B1(G50), .B2(new_n252), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(KEYINPUT74), .A3(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n270), .A2(KEYINPUT74), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(KEYINPUT74), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n272), .B(new_n273), .C1(new_n267), .C2(new_n268), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(KEYINPUT67), .A3(new_n206), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT67), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  INV_X1    g0084(.A(new_n225), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G226), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n206), .A2(new_n278), .B1(new_n285), .B2(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT3), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n298), .A2(G223), .B1(G77), .B2(new_n296), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT3), .B(G33), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G222), .A3(new_n297), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n285), .A2(new_n286), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n288), .B1(new_n289), .B2(new_n291), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT75), .B1(new_n304), .B2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT75), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(G200), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n275), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n306), .B2(new_n304), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n271), .B2(new_n274), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G179), .B2(new_n304), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n269), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n256), .A2(new_n258), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n250), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n322), .B2(new_n252), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n325), .A2(new_n326), .A3(new_n292), .ZN(new_n327));
  INV_X1    g0127(.A(new_n293), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT7), .B1(new_n329), .B2(G20), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT81), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n294), .ZN(new_n332));
  NAND2_X1  g0132(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(G33), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(G20), .B1(new_n334), .B2(new_n293), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT7), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n213), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  INV_X1    g0139(.A(new_n263), .ZN(new_n340));
  INV_X1    g0140(.A(G159), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT65), .B(G68), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n228), .B1(new_n343), .B2(new_n257), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n339), .B(new_n342), .C1(new_n344), .C2(G20), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n253), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n336), .A2(G20), .ZN(new_n347));
  AOI21_X1  g0147(.A(G33), .B1(new_n332), .B2(new_n333), .ZN(new_n348));
  INV_X1    g0148(.A(new_n295), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n336), .B1(new_n300), .B2(G20), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n343), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n201), .B1(new_n217), .B2(G58), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n353), .A2(new_n207), .B1(new_n341), .B2(new_n340), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n339), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n324), .B1(new_n346), .B2(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n283), .A2(new_n287), .B1(new_n290), .B2(G232), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(G223), .A2(G1698), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n289), .B2(G1698), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n334), .A3(new_n293), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G87), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT82), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n303), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(G200), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n361), .A2(new_n363), .ZN(new_n366));
  OAI211_X1 g0166(.A(G190), .B(new_n357), .C1(new_n366), .C2(new_n303), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n356), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n356), .A2(KEYINPUT17), .A3(new_n368), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(G169), .B1(new_n358), .B2(new_n364), .ZN(new_n374));
  OAI211_X1 g0174(.A(G179), .B(new_n357), .C1(new_n366), .C2(new_n303), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT18), .B1(new_n356), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n335), .A2(new_n336), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n336), .B(new_n207), .C1(new_n327), .C2(new_n328), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n345), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(new_n355), .A3(new_n249), .ZN(new_n382));
  INV_X1    g0182(.A(new_n324), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT18), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n374), .A2(new_n375), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n377), .A2(KEYINPUT83), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT83), .B1(new_n377), .B2(new_n387), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n373), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n283), .A2(new_n287), .B1(new_n290), .B2(G238), .ZN(new_n391));
  INV_X1    g0191(.A(G232), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(G226), .B2(G1698), .ZN(new_n394));
  INV_X1    g0194(.A(G97), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n394), .A2(new_n296), .B1(new_n292), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(G33), .A2(G41), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n225), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT77), .B1(new_n400), .B2(KEYINPUT13), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n391), .A2(new_n402), .A3(new_n399), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT13), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(KEYINPUT76), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n405), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n391), .A2(new_n399), .A3(new_n402), .A4(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n401), .A2(new_n406), .A3(G190), .A4(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n400), .A2(KEYINPUT13), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n404), .B1(new_n391), .B2(new_n399), .ZN(new_n411));
  OAI21_X1  g0211(.A(G200), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT12), .B1(new_n217), .B2(new_n252), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT78), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT78), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(KEYINPUT12), .C1(new_n217), .C2(new_n252), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OR3_X1    g0217(.A1(new_n252), .A2(KEYINPUT12), .A3(G68), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(G68), .B2(new_n250), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n217), .A2(new_n207), .ZN(new_n420));
  INV_X1    g0220(.A(G77), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n340), .A2(new_n202), .B1(new_n260), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n249), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT11), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(new_n249), .C1(new_n420), .C2(new_n422), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n419), .A2(KEYINPUT79), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT79), .B1(new_n419), .B2(new_n427), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n409), .B(new_n412), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT80), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n419), .A2(new_n427), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT79), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n419), .A2(KEYINPUT79), .A3(new_n427), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT80), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n409), .A4(new_n412), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G169), .B1(new_n410), .B2(new_n411), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n401), .A2(new_n406), .A3(G179), .A4(new_n408), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(G169), .C1(new_n410), .C2(new_n411), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n436), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g0248(.A(KEYINPUT8), .B(G58), .Z(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT15), .B(G87), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT71), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n261), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT71), .B1(new_n451), .B2(new_n260), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n450), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n249), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n252), .A2(G77), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n250), .B2(G77), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT72), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n300), .A2(G232), .A3(new_n297), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT70), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT70), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n300), .A2(new_n465), .A3(G232), .A4(new_n297), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n298), .A2(G238), .B1(G107), .B2(new_n296), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n303), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G244), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n288), .B1(new_n470), .B2(new_n291), .ZN(new_n471));
  OAI21_X1  g0271(.A(G200), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n457), .A2(KEYINPUT72), .A3(new_n459), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n462), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT73), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT73), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n462), .A2(new_n472), .A3(new_n476), .A4(new_n473), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n469), .A2(new_n471), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G190), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n462), .A2(new_n473), .ZN(new_n481));
  INV_X1    g0281(.A(G179), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n316), .B1(new_n469), .B2(new_n471), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NOR4_X1   g0286(.A1(new_n321), .A2(new_n390), .A3(new_n448), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n206), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n253), .A2(KEYINPUT84), .A3(new_n252), .A4(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT84), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n252), .A2(new_n488), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n249), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n492), .A3(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT92), .A2(KEYINPUT25), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n206), .A2(new_n496), .A3(G13), .A4(G20), .ZN(new_n497));
  MUX2_X1   g0297(.A(new_n494), .B(new_n495), .S(new_n497), .Z(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT93), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n493), .A2(KEYINPUT93), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT91), .B1(new_n496), .B2(G20), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI211_X1 g0306(.A(KEYINPUT91), .B(KEYINPUT23), .C1(new_n496), .C2(G20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n506), .A2(new_n507), .B1(G20), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G87), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n510), .A2(KEYINPUT22), .A3(G20), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n300), .A2(KEYINPUT90), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT90), .B1(new_n300), .B2(new_n511), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n334), .A2(new_n207), .A3(G87), .A4(new_n293), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n509), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n249), .B1(new_n517), .B2(KEYINPUT24), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT24), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n519), .B(new_n509), .C1(new_n514), .C2(new_n516), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n503), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G250), .A2(G1698), .ZN(new_n522));
  INV_X1    g0322(.A(G257), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(G1698), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n524), .A2(new_n334), .A3(new_n293), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT94), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(KEYINPUT94), .A3(new_n526), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n398), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(KEYINPUT5), .A2(G41), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(KEYINPUT5), .A2(G41), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n206), .B(G45), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(G274), .B1(new_n397), .B2(new_n225), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT85), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n206), .A2(G45), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT5), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n276), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n538), .B1(new_n540), .B2(new_n532), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT85), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n287), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n535), .A2(new_n303), .ZN(new_n545));
  INV_X1    g0345(.A(G264), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n531), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n316), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n303), .B1(new_n527), .B2(new_n528), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n547), .B1(new_n551), .B2(new_n530), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(new_n482), .A3(new_n544), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n521), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G283), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n555), .B(new_n207), .C1(G33), .C2(new_n395), .ZN(new_n556));
  INV_X1    g0356(.A(G116), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n249), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n556), .A2(KEYINPUT20), .A3(new_n249), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n252), .A2(G116), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n491), .A2(new_n249), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(G116), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n316), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n546), .A2(new_n297), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n334), .A2(new_n293), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT89), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n334), .A2(KEYINPUT89), .A3(new_n293), .A4(new_n568), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n334), .A2(G257), .A3(new_n297), .A4(new_n293), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n296), .A2(G303), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n303), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n541), .A2(new_n398), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n537), .A2(new_n543), .B1(new_n578), .B2(G270), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n567), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n567), .B(KEYINPUT21), .C1(new_n577), .C2(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n573), .A2(new_n576), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n398), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n563), .A2(new_n566), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(G179), .A3(new_n579), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n554), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n252), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n395), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n489), .A2(new_n492), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n395), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n496), .B1(new_n350), .B2(new_n351), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n596), .A2(new_n395), .A3(G107), .ZN(new_n597));
  XNOR2_X1  g0397(.A(G97), .B(G107), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI22_X1  g0399(.A1(new_n599), .A2(new_n207), .B1(new_n421), .B2(new_n340), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n594), .B1(new_n601), .B2(new_n249), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n334), .A2(G244), .A3(new_n297), .A4(new_n293), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT4), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(KEYINPUT4), .A2(G244), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n293), .A2(new_n295), .A3(new_n606), .A4(new_n297), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n293), .A2(new_n295), .A3(G250), .A4(G1698), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n607), .A2(new_n608), .A3(new_n555), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n303), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT85), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n542), .B1(new_n541), .B2(new_n287), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n611), .A2(new_n612), .B1(new_n523), .B2(new_n545), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G190), .ZN(new_n615));
  OAI21_X1  g0415(.A(G200), .B1(new_n610), .B2(new_n613), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n602), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(G169), .B1(new_n610), .B2(new_n613), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n537), .A2(new_n543), .B1(new_n578), .B2(G257), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n607), .A2(new_n608), .A3(new_n555), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n604), .B2(new_n603), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n619), .B(G179), .C1(new_n621), .C2(new_n303), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n249), .B1(new_n595), .B2(new_n600), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n592), .C1(new_n395), .C2(new_n593), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT86), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT86), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n623), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n617), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(G200), .B1(new_n577), .B2(new_n580), .ZN(new_n631));
  INV_X1    g0431(.A(new_n587), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n574), .A2(new_n575), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n571), .B2(new_n572), .ZN(new_n634));
  OAI211_X1 g0434(.A(G190), .B(new_n579), .C1(new_n634), .C2(new_n303), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n549), .A2(new_n306), .ZN(new_n637));
  INV_X1    g0437(.A(G200), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n552), .B2(new_n544), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n521), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n636), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n334), .A2(new_n207), .A3(G68), .A4(new_n293), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n260), .A2(new_n395), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(KEYINPUT19), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n207), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n510), .A2(new_n395), .A3(new_n496), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT87), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT87), .B1(new_n647), .B2(new_n648), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n249), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n451), .A2(new_n591), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n489), .A2(new_n492), .A3(new_n452), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(G238), .A2(G1698), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n470), .B2(G1698), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n334), .A3(new_n293), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n303), .B1(new_n658), .B2(new_n508), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n303), .A2(G250), .A3(new_n538), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n536), .B2(new_n538), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n482), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n316), .B1(new_n659), .B2(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n655), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(G200), .B1(new_n659), .B2(new_n661), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n489), .A2(new_n492), .A3(G87), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n652), .A3(new_n653), .A4(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n669), .A2(KEYINPUT88), .B1(G190), .B2(new_n662), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n652), .A2(new_n653), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(new_n667), .A4(new_n668), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n666), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n590), .A2(new_n630), .A3(new_n642), .A4(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n487), .A2(new_n676), .ZN(G372));
  OAI21_X1  g0477(.A(KEYINPUT96), .B1(new_n356), .B2(new_n376), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT96), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n384), .A2(new_n679), .A3(new_n386), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n385), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(new_n680), .A3(KEYINPUT18), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n485), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n439), .A2(new_n685), .B1(new_n446), .B2(new_n445), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n371), .A2(new_n372), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n319), .B1(new_n688), .B2(new_n315), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n623), .A2(new_n625), .A3(new_n628), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n628), .B1(new_n623), .B2(new_n625), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(KEYINPUT26), .A3(new_n674), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n655), .A2(new_n665), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n659), .A2(new_n661), .A3(new_n306), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n669), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n623), .A2(KEYINPUT95), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT95), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n618), .A2(new_n622), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n702), .A3(new_n625), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n695), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n694), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n588), .A2(new_n584), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n579), .B1(new_n634), .B2(new_n303), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT21), .B1(new_n707), .B2(new_n567), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n521), .A2(new_n550), .A3(new_n553), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n514), .A2(new_n516), .ZN(new_n712));
  INV_X1    g0512(.A(new_n509), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n519), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n517), .A2(KEYINPUT24), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n249), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n549), .A2(G200), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n552), .A2(G190), .A3(new_n544), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n503), .A4(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n630), .A2(new_n711), .A3(new_n720), .A4(new_n698), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n705), .A2(new_n721), .A3(new_n696), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n690), .B1(new_n487), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT97), .ZN(G369));
  NAND3_X1  g0524(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(KEYINPUT27), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT98), .Z(new_n727));
  INV_X1    g0527(.A(G213), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n725), .B2(KEYINPUT27), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n727), .A2(G343), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n587), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n589), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(new_n731), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n732), .B1(new_n734), .B2(new_n589), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT99), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n730), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n720), .B1(new_n641), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n710), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n554), .A2(new_n739), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n589), .A2(new_n739), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n741), .A2(new_n747), .B1(new_n554), .B2(new_n739), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n745), .A2(new_n748), .ZN(G399));
  NAND2_X1  g0549(.A1(new_n210), .A2(new_n276), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n648), .A2(G116), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(G1), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n229), .B2(new_n750), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n693), .A2(new_n695), .A3(new_n674), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT26), .B1(new_n699), .B2(new_n703), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n721), .A2(new_n696), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n739), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT29), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n722), .A2(new_n739), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(KEYINPUT29), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT31), .B1(new_n675), .B2(new_n730), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n707), .A2(new_n482), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n763), .A2(new_n614), .A3(new_n662), .A4(new_n552), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT30), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n614), .A2(G179), .A3(new_n662), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(new_n707), .A3(new_n549), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n730), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n730), .A2(KEYINPUT31), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n770), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT100), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n766), .B1(new_n775), .B2(KEYINPUT100), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n761), .B1(G330), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n754), .B1(new_n780), .B2(G1), .ZN(G364));
  INV_X1    g0581(.A(new_n750), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n207), .A2(G13), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n206), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n738), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G330), .B2(new_n736), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n210), .A2(new_n300), .ZN(new_n789));
  INV_X1    g0589(.A(G355), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(G116), .B2(new_n210), .ZN(new_n791));
  INV_X1    g0591(.A(new_n329), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n210), .ZN(new_n793));
  INV_X1    g0593(.A(new_n229), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(new_n277), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n243), .A2(new_n277), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n225), .B1(G20), .B2(new_n316), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n786), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n482), .A2(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n207), .A2(G190), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n300), .B1(new_n807), .B2(new_n421), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n207), .A2(new_n306), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n482), .A2(new_n638), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n805), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n811), .A2(new_n202), .B1(new_n812), .B2(new_n257), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n482), .A2(G200), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT101), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n806), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n808), .B(new_n813), .C1(new_n819), .C2(G107), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n810), .A2(new_n806), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT102), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n821), .A2(new_n822), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n817), .A2(new_n809), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n827), .A2(G68), .B1(new_n829), .B2(G87), .ZN(new_n830));
  NOR2_X1   g0630(.A1(G179), .A2(G200), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n806), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G159), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT32), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n831), .A2(G190), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G20), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n834), .A2(KEYINPUT32), .B1(G97), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n820), .A2(new_n830), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT33), .B(G317), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n827), .A2(new_n840), .B1(new_n819), .B2(G283), .ZN(new_n841));
  INV_X1    g0641(.A(G326), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n296), .B1(new_n811), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G322), .ZN(new_n844));
  INV_X1    g0644(.A(G311), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n812), .A2(new_n844), .B1(new_n807), .B2(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n843), .B(new_n846), .C1(G294), .C2(new_n837), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n833), .A2(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n833), .A2(KEYINPUT103), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G329), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n829), .A2(G303), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n841), .A2(new_n847), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n839), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n804), .B1(new_n801), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n800), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n736), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n788), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G396));
  INV_X1    g0660(.A(new_n786), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n779), .A2(G330), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n481), .A2(new_n730), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n685), .B1(new_n480), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n485), .A2(new_n730), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n760), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n722), .A2(new_n739), .A3(new_n866), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n861), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n862), .A2(new_n870), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(KEYINPUT106), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(KEYINPUT106), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n801), .A2(new_n798), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n861), .B1(new_n421), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n801), .ZN(new_n877));
  INV_X1    g0677(.A(new_n811), .ZN(new_n878));
  INV_X1    g0678(.A(new_n807), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n878), .A2(G137), .B1(new_n879), .B2(G159), .ZN(new_n880));
  INV_X1    g0680(.A(G143), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(new_n812), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G150), .B2(new_n827), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(KEYINPUT34), .ZN(new_n884));
  INV_X1    g0684(.A(new_n837), .ZN(new_n885));
  INV_X1    g0685(.A(G132), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n329), .B1(new_n257), .B2(new_n885), .C1(new_n850), .C2(new_n886), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n202), .A2(new_n828), .B1(new_n818), .B2(new_n213), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n883), .A2(KEYINPUT34), .ZN(new_n890));
  INV_X1    g0690(.A(new_n812), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n891), .A2(G294), .B1(new_n837), .B2(G97), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT105), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n510), .A2(new_n818), .B1(new_n828), .B2(new_n496), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n296), .B1(new_n850), .B2(new_n845), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G303), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n811), .A2(new_n897), .B1(new_n807), .B2(new_n557), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n827), .B2(G283), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT104), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n889), .A2(new_n890), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n876), .B1(new_n877), .B2(new_n901), .C1(new_n866), .C2(new_n799), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n874), .A2(new_n902), .ZN(G384));
  NAND2_X1  g0703(.A1(new_n598), .A2(new_n596), .ZN(new_n904));
  INV_X1    g0704(.A(new_n597), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n906), .A2(KEYINPUT35), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(KEYINPUT35), .ZN(new_n908));
  NOR4_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(new_n227), .A4(new_n557), .ZN(new_n909));
  XOR2_X1   g0709(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n794), .B(G77), .C1(new_n257), .C2(new_n343), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n202), .A2(G68), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n206), .B(G13), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT112), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n381), .A2(new_n249), .ZN(new_n917));
  INV_X1    g0717(.A(new_n354), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT16), .B1(new_n338), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n383), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n386), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n727), .A2(new_n729), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n921), .A2(new_n924), .A3(new_n369), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT37), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT37), .B1(new_n356), .B2(new_n368), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n384), .B1(new_n386), .B2(new_n923), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT83), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n356), .A2(new_n376), .A3(KEYINPUT18), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n377), .A2(new_n387), .A3(KEYINPUT83), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n687), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n930), .B1(new_n936), .B2(new_n924), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(KEYINPUT38), .B(new_n930), .C1(new_n936), .C2(new_n924), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(KEYINPUT108), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT108), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n942), .A3(new_n938), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(KEYINPUT39), .A3(new_n943), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n925), .A2(KEYINPUT37), .B1(new_n927), .B2(new_n928), .ZN(new_n945));
  INV_X1    g0745(.A(new_n924), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n945), .B1(new_n390), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT39), .B1(new_n947), .B2(KEYINPUT38), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n384), .A2(new_n923), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n684), .B2(new_n373), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n356), .A2(new_n376), .A3(KEYINPUT96), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n679), .B1(new_n384), .B2(new_n386), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n369), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT109), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n678), .A2(new_n680), .B1(new_n356), .B2(new_n368), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(KEYINPUT109), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT37), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n929), .B(KEYINPUT110), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n950), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n948), .B(KEYINPUT111), .C1(new_n960), .C2(KEYINPUT38), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n944), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n929), .B(KEYINPUT110), .Z(new_n963));
  NAND2_X1  g0763(.A1(new_n953), .A2(new_n954), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n956), .A2(KEYINPUT109), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n964), .A2(new_n965), .A3(new_n949), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n966), .B2(KEYINPUT37), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n938), .B1(new_n967), .B2(new_n950), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT111), .B1(new_n968), .B2(new_n948), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n916), .B1(new_n962), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n948), .B1(new_n960), .B2(KEYINPUT38), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT111), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n973), .A2(KEYINPUT112), .A3(new_n944), .A4(new_n961), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n447), .A2(new_n730), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n941), .A2(new_n943), .ZN(new_n978));
  INV_X1    g0778(.A(new_n865), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n869), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n446), .A2(new_n730), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n439), .A2(new_n447), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n981), .B1(new_n439), .B2(new_n447), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n978), .A2(new_n986), .B1(new_n684), .B2(new_n923), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n977), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n487), .A2(new_n761), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n689), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n989), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n866), .B1(new_n982), .B2(new_n983), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n709), .A2(new_n710), .A3(new_n720), .A4(new_n733), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n602), .A2(new_n615), .A3(new_n616), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n691), .B2(new_n692), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n670), .A2(new_n673), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n696), .ZN(new_n998));
  NOR4_X1   g0798(.A1(new_n994), .A2(new_n996), .A3(new_n998), .A4(new_n730), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT31), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n772), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n775), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n774), .B1(new_n1002), .B2(new_n767), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n993), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n941), .A2(new_n1005), .A3(new_n943), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT40), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n940), .B1(new_n960), .B2(KEYINPUT38), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1003), .B1(new_n762), .B2(new_n772), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1009), .A2(new_n1007), .A3(new_n993), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1006), .A2(new_n1007), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(new_n487), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(G330), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1011), .B1(new_n487), .B2(new_n1012), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n992), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n206), .B2(new_n783), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n992), .A2(new_n1016), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n915), .B1(new_n1018), .B2(new_n1019), .ZN(G367));
  OAI221_X1 g0820(.A(new_n802), .B1(new_n210), .B2(new_n451), .C1(new_n793), .C2(new_n239), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(new_n786), .ZN(new_n1022));
  INV_X1    g0822(.A(G150), .ZN(new_n1023));
  INV_X1    g0823(.A(G137), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n812), .A2(new_n1023), .B1(new_n832), .B2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n300), .B1(new_n811), .B2(new_n881), .C1(new_n885), .C2(new_n213), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(G50), .C2(new_n879), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n827), .A2(G159), .B1(new_n819), .B2(G77), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n257), .C2(new_n828), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n827), .A2(G294), .B1(new_n819), .B2(G97), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G311), .A2(new_n878), .B1(new_n891), .B2(G303), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT117), .B(G317), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n833), .A2(new_n1033), .B1(new_n879), .B2(G283), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n329), .B1(G107), .B2(new_n837), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n828), .A2(new_n557), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT46), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1029), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT47), .Z(new_n1040));
  AOI21_X1  g0840(.A(new_n739), .B1(new_n671), .B2(new_n668), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT113), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(new_n696), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n696), .A3(new_n698), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1022), .B1(new_n1040), .B2(new_n877), .C1(new_n1045), .C2(new_n857), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n743), .B(new_n747), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(new_n737), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n780), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n630), .B1(new_n602), .B2(new_n739), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n703), .A2(new_n739), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n748), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT45), .Z(new_n1055));
  NOR2_X1   g0855(.A1(new_n748), .A2(new_n1053), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT44), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n745), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(KEYINPUT116), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT116), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1055), .B(new_n1057), .C1(new_n1061), .C2(new_n745), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1050), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n780), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n750), .B(KEYINPUT41), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n785), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n743), .A2(new_n746), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1053), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT42), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1068), .A2(new_n710), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n739), .B1(new_n1071), .B2(new_n693), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1045), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT43), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1045), .A2(KEYINPUT43), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1070), .A2(new_n1075), .A3(new_n1074), .A4(new_n1072), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT114), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1059), .A2(new_n1080), .A3(new_n1053), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT114), .B1(new_n745), .B2(new_n1068), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT115), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1078), .B(new_n1079), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1078), .A2(new_n1083), .A3(new_n1084), .A4(new_n1079), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1046), .B1(new_n1066), .B2(new_n1089), .ZN(G387));
  OAI22_X1  g0890(.A1(new_n789), .A2(new_n751), .B1(G107), .B2(new_n210), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n236), .A2(new_n277), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n751), .ZN(new_n1093));
  AOI211_X1 g0893(.A(G45), .B(new_n1093), .C1(G68), .C2(G77), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n254), .A2(G50), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT50), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n793), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1091), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n792), .B1(new_n842), .B2(new_n832), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n891), .A2(new_n1033), .B1(new_n878), .B2(G322), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n897), .B2(new_n807), .C1(new_n826), .C2(new_n845), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT48), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n829), .A2(G294), .B1(G283), .B2(new_n837), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT49), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1099), .B(new_n1108), .C1(G116), .C2(new_n819), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n829), .A2(G77), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT119), .B(G150), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n792), .B1(new_n833), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(new_n395), .C2(new_n818), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT120), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n878), .A2(G159), .B1(new_n879), .B2(G68), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n202), .B2(new_n812), .C1(new_n451), .C2(new_n885), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n259), .B2(new_n827), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1109), .A2(new_n1110), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n786), .B1(new_n803), .B2(new_n1098), .C1(new_n1119), .C2(new_n877), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n743), .B2(new_n800), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1048), .A2(new_n785), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1122), .A2(KEYINPUT118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(KEYINPUT118), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n780), .A2(new_n1048), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1049), .A2(new_n782), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(G393));
  XNOR2_X1  g0928(.A(new_n1058), .B(new_n745), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n785), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n802), .B1(new_n395), .B2(new_n210), .C1(new_n793), .C2(new_n246), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n786), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G107), .A2(new_n819), .B1(new_n829), .B2(G283), .ZN(new_n1133));
  INV_X1    g0933(.A(G317), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n811), .A2(new_n1134), .B1(new_n812), .B2(new_n845), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT52), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n827), .A2(G303), .B1(new_n1136), .B2(new_n1135), .ZN(new_n1138));
  INV_X1    g0938(.A(G294), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n296), .B1(new_n832), .B2(new_n844), .C1(new_n1139), .C2(new_n807), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(G116), .B2(new_n837), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1133), .A2(new_n1137), .A3(new_n1138), .A4(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n811), .A2(new_n1023), .B1(new_n812), .B2(new_n341), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT51), .Z(new_n1144));
  OAI22_X1  g0944(.A1(new_n510), .A2(new_n818), .B1(new_n828), .B2(new_n343), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n329), .B1(new_n881), .B2(new_n832), .C1(new_n421), .C2(new_n885), .ZN(new_n1146));
  OR3_X1    g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n826), .A2(new_n202), .B1(new_n254), .B2(new_n807), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT121), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1142), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1132), .B1(new_n1150), .B2(new_n801), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1053), .B2(new_n857), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1063), .A2(new_n782), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1129), .A2(new_n1050), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1130), .B(new_n1152), .C1(new_n1153), .C2(new_n1154), .ZN(G390));
  INV_X1    g0955(.A(new_n976), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT122), .B1(new_n986), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT122), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1158), .B(new_n976), .C1(new_n980), .C2(new_n985), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n970), .A2(new_n974), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n758), .A2(new_n864), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n865), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1156), .B(new_n1008), .C1(new_n1163), .C2(new_n984), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G330), .B(new_n866), .C1(new_n773), .C2(new_n778), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(new_n984), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1161), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1012), .A2(G330), .A3(new_n866), .A4(new_n985), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n970), .A2(new_n798), .A3(new_n974), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n875), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n786), .B1(new_n259), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G116), .A2(new_n891), .B1(new_n879), .B2(G97), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n300), .B1(new_n878), .B2(G283), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n421), .C2(new_n885), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G68), .A2(new_n819), .B1(new_n829), .B2(G87), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n496), .B2(new_n826), .C1(new_n1139), .C2(new_n850), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n829), .A2(new_n1112), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT53), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT53), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n837), .A2(G159), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT54), .B(G143), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n812), .A2(new_n886), .B1(new_n807), .B2(new_n1183), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n296), .B(new_n1184), .C1(G128), .C2(new_n878), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n851), .A2(G125), .B1(new_n819), .B2(G50), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1024), .B2(new_n826), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1176), .A2(new_n1178), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1173), .B1(new_n1189), .B2(new_n801), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1170), .A2(new_n785), .B1(new_n1171), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n984), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1168), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n980), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1012), .A2(G330), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n985), .B1(new_n1195), .B2(new_n866), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1163), .B1(new_n1165), .B2(new_n984), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n487), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n990), .A3(new_n689), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1168), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1161), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1192), .A2(new_n1168), .B1(new_n979), .B2(new_n869), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(new_n1200), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1206), .A2(new_n1207), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1203), .A2(new_n1212), .A3(new_n782), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1191), .A2(new_n1213), .ZN(G378));
  NAND2_X1  g1014(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n269), .A2(new_n922), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n315), .A2(new_n320), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n315), .B2(new_n320), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1217), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n321), .A2(new_n1218), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n315), .A2(new_n320), .A3(new_n1219), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(new_n1224), .A3(new_n1216), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1010), .A2(new_n1008), .ZN(new_n1227));
  AND4_X1   g1027(.A1(G330), .A2(new_n1215), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1226), .B1(new_n1011), .B2(G330), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n977), .A3(new_n988), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1156), .B1(new_n970), .B2(new_n974), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1232), .A2(new_n987), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1222), .A2(new_n1225), .A3(new_n798), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n786), .B1(G50), .B2(new_n1172), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G41), .B1(new_n879), .B2(new_n452), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(new_n496), .B2(new_n812), .C1(new_n557), .C2(new_n811), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n329), .B(new_n1238), .C1(G68), .C2(new_n837), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n818), .A2(new_n257), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n851), .A2(G283), .B1(new_n827), .B2(G97), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1239), .A2(new_n1111), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT58), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n292), .B1(new_n332), .B2(new_n333), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n202), .B1(new_n1245), .B2(G41), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1183), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n827), .A2(G132), .B1(new_n829), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n837), .A2(G150), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n879), .A2(G137), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G125), .A2(new_n878), .B1(new_n891), .B2(G128), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n819), .A2(G159), .ZN(new_n1255));
  AOI211_X1 g1055(.A(G33), .B(G41), .C1(new_n833), .C2(G124), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1244), .B(new_n1246), .C1(new_n1253), .C2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT123), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n877), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1236), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1234), .A2(new_n785), .B1(new_n1235), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT57), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1167), .A2(new_n1169), .A3(new_n1202), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(new_n1200), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n782), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1212), .A2(new_n1201), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT57), .B1(new_n1269), .B2(new_n1234), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1263), .B1(new_n1268), .B2(new_n1270), .ZN(G375));
  AOI21_X1  g1071(.A(new_n861), .B1(new_n213), .B2(new_n875), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n811), .A2(new_n886), .B1(new_n812), .B2(new_n1024), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n329), .B1(new_n202), .B2(new_n885), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(G150), .C2(new_n879), .ZN(new_n1275));
  INV_X1    g1075(.A(G128), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n850), .A2(new_n1276), .B1(new_n828), .B2(new_n341), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1240), .B(new_n1277), .C1(new_n827), .C2(new_n1247), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n300), .B1(new_n891), .B2(G283), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1279), .B1(new_n1139), .B2(new_n811), .C1(new_n451), .C2(new_n885), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n421), .A2(new_n818), .B1(new_n828), .B2(new_n395), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(G303), .C2(new_n851), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n826), .A2(new_n557), .B1(new_n496), .B2(new_n807), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(KEYINPUT124), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1275), .A2(new_n1278), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  OAI221_X1 g1085(.A(new_n1272), .B1(new_n877), .B2(new_n1285), .C1(new_n985), .C2(new_n799), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1210), .B2(new_n784), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1202), .A2(new_n1065), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(G381));
  NOR4_X1   g1091(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1292), .B(new_n1046), .C1(new_n1066), .C2(new_n1089), .ZN(new_n1293));
  OR4_X1    g1093(.A1(G378), .A2(G375), .A3(new_n1293), .A4(G381), .ZN(G407));
  INV_X1    g1094(.A(G375), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1191), .A2(new_n1213), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n728), .A2(G343), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(G407), .A2(G213), .A3(new_n1298), .ZN(G409));
  INV_X1    g1099(.A(G390), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G387), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G390), .B(new_n1046), .C1(new_n1066), .C2(new_n1089), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(new_n859), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1301), .A2(new_n1304), .A3(new_n1302), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1309), .B(new_n1310), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G378), .B(new_n1263), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1269), .A2(new_n1065), .A3(new_n1234), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1263), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1296), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1297), .B1(new_n1312), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n874), .A2(new_n1318), .A3(new_n902), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT60), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(new_n1290), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1210), .A2(KEYINPUT60), .A3(new_n1200), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n782), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1288), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1320), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1288), .B(new_n1319), .C1(new_n1323), .C2(new_n1325), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1316), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1297), .A2(G2897), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1327), .A2(new_n1328), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1334), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  OR2_X1    g1138(.A1(new_n1316), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1316), .A2(KEYINPUT63), .A3(new_n1330), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1311), .A2(new_n1333), .A3(new_n1339), .A4(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1316), .A2(new_n1342), .A3(new_n1330), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1344), .B1(new_n1316), .B2(new_n1338), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1342), .B1(new_n1316), .B2(new_n1330), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1343), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1341), .B1(new_n1347), .B2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(G375), .A2(new_n1296), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1312), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1330), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1351), .A2(new_n1312), .A3(new_n1329), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1355), .B(new_n1348), .ZN(G402));
endmodule


