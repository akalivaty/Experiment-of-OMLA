//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n461), .A2(new_n462), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n461), .B1(G2104), .B2(new_n462), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI22_X1  g044(.A1(new_n465), .A2(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n462), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n470), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(new_n468), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  XOR2_X1   g050(.A(KEYINPUT3), .B(G2104), .Z(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n462), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n462), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n475), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT68), .ZN(G162));
  OAI21_X1  g057(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n462), .A2(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n476), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n467), .A2(G138), .A3(new_n462), .A4(new_n486), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n467), .A2(G126), .A3(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n467), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT5), .B(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT71), .B1(new_n502), .B2(KEYINPUT6), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n499), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n500), .B2(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n502), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n511), .A2(KEYINPUT72), .A3(new_n499), .A4(new_n501), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n511), .A2(G543), .A3(new_n501), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n516), .A2(G50), .B1(new_n522), .B2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n515), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n499), .A2(KEYINPUT73), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n518), .A2(new_n527), .A3(new_n519), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(G51), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n514), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n514), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n529), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n543), .A2(G651), .B1(G52), .B2(new_n516), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n529), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n551), .B(new_n547), .C1(new_n529), .C2(new_n548), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n550), .A2(G651), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n507), .A2(G81), .A3(new_n512), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n516), .A2(G43), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n554), .A2(KEYINPUT76), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT76), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n553), .B(KEYINPUT77), .C1(new_n556), .C2(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  AND2_X1   g143(.A1(new_n499), .A2(G65), .ZN(new_n569));
  AND2_X1   g144(.A1(G78), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n516), .A2(new_n573), .A3(G53), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(new_n516), .B2(G53), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n571), .B1(new_n513), .B2(new_n572), .C1(new_n574), .C2(new_n575), .ZN(G299));
  NAND4_X1  g151(.A1(new_n511), .A2(G49), .A3(G543), .A4(new_n501), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n507), .A2(G87), .A3(new_n512), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n520), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n516), .A2(G48), .B1(new_n585), .B2(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n507), .A2(G86), .A3(new_n512), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n529), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n502), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(new_n591), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n514), .A2(G85), .B1(G47), .B2(new_n516), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n520), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n516), .A2(G54), .B1(new_n600), .B2(G651), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n514), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT10), .B1(new_n514), .B2(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n597), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n562), .A2(new_n608), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n604), .A2(G559), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT80), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n474), .A2(G135), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT82), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n477), .A2(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n462), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NOR2_X1   g200(.A1(new_n465), .A2(new_n476), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(G2100), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n625), .A2(new_n630), .A3(new_n631), .ZN(G156));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(KEYINPUT14), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G14), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n643), .A2(new_n646), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT85), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT17), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT87), .Z(new_n658));
  INV_X1    g233(.A(new_n656), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n652), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n653), .A2(new_n655), .ZN(new_n663));
  INV_X1    g238(.A(new_n652), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n664), .B2(new_n654), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n658), .B(new_n662), .C1(new_n663), .C2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n670), .A2(new_n675), .A3(new_n673), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n678));
  AOI211_X1 g253(.A(new_n674), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n677), .B2(new_n678), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  NAND3_X1  g261(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT25), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n474), .A2(G139), .ZN(new_n690));
  AOI22_X1  g265(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n689), .B(new_n690), .C1(new_n462), .C2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G33), .B(new_n692), .S(G29), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G2072), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT95), .Z(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G26), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n474), .A2(G140), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n477), .A2(G128), .ZN(new_n700));
  OR2_X1    g275(.A1(G104), .A2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n698), .B1(new_n704), .B2(new_n696), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G2067), .ZN(new_n706));
  INV_X1    g281(.A(G2078), .ZN(new_n707));
  NOR2_X1   g282(.A1(G164), .A2(new_n696), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G27), .B2(new_n696), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n706), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n695), .B(new_n710), .C1(new_n707), .C2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n693), .A2(G2072), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT93), .Z(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NOR2_X1   g289(.A1(G171), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G5), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G1961), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n713), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT30), .B(G28), .ZN(new_n721));
  OR2_X1    g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  NAND2_X1  g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n721), .A2(new_n696), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n624), .B2(new_n696), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n696), .A2(G32), .ZN(new_n726));
  INV_X1    g301(.A(new_n465), .ZN(new_n727));
  AOI22_X1  g302(.A1(G105), .A2(new_n727), .B1(new_n474), .B2(G141), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT26), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n477), .B2(G129), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n726), .B1(new_n732), .B2(G29), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n725), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n696), .B1(new_n738), .B2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G160), .B2(G29), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(G2084), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT98), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(G2084), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT94), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n737), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n711), .A2(new_n720), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G21), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT96), .B1(new_n714), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G168), .A2(G16), .ZN(new_n750));
  MUX2_X1   g325(.A(KEYINPUT96), .B(new_n749), .S(new_n750), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G1966), .ZN(new_n752));
  NOR2_X1   g327(.A1(G29), .A2(G35), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G162), .B2(G29), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT29), .Z(new_n755));
  INV_X1    g330(.A(G2090), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n756), .B2(new_n755), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n604), .A2(new_n714), .ZN(new_n759));
  NOR2_X1   g334(.A1(G4), .A2(G16), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G1348), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n714), .A2(G20), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT23), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G299), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G1348), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n759), .A2(new_n768), .A3(new_n760), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n762), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n751), .A2(G1966), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n747), .A2(new_n758), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n714), .A2(G19), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n563), .B2(new_n714), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1341), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n714), .A2(G22), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G166), .B2(new_n714), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT90), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G1971), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n714), .A2(G23), .ZN(new_n783));
  INV_X1    g358(.A(G288), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n714), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT33), .B(G1976), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G6), .B(G305), .S(G16), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  INV_X1    g365(.A(G1981), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n781), .A2(G1971), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n788), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT34), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n788), .A2(new_n796), .A3(new_n792), .A4(new_n793), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n798));
  NOR2_X1   g373(.A1(G25), .A2(G29), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n477), .A2(G119), .ZN(new_n800));
  OR2_X1    g375(.A1(G95), .A2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n801), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G131), .B2(new_n474), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n799), .B1(new_n804), .B2(G29), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT89), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G1991), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  MUX2_X1   g383(.A(G24), .B(G290), .S(G16), .Z(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(G1986), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(G1986), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n797), .A2(new_n798), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n798), .B1(new_n797), .B2(new_n812), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n795), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT36), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n797), .A2(new_n812), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT91), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n813), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n820), .A2(new_n821), .A3(new_n795), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n778), .B1(new_n817), .B2(new_n822), .ZN(G311));
  AOI21_X1  g398(.A(new_n821), .B1(new_n820), .B2(new_n795), .ZN(new_n824));
  INV_X1    g399(.A(new_n795), .ZN(new_n825));
  AOI211_X1 g400(.A(KEYINPUT36), .B(new_n825), .C1(new_n819), .C2(new_n813), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n777), .B1(new_n824), .B2(new_n826), .ZN(G150));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n529), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G651), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n507), .A2(G93), .A3(new_n512), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n516), .A2(G55), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G860), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n604), .A2(new_n612), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n834), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n562), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n834), .B(new_n553), .C1(new_n556), .C2(new_n557), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n835), .B1(new_n846), .B2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n837), .B1(new_n847), .B2(new_n848), .ZN(G145));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n491), .A2(new_n850), .A3(new_n496), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n491), .B2(new_n496), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n704), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n732), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n692), .A2(KEYINPUT102), .ZN(new_n857));
  OR3_X1    g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n692), .A2(new_n856), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n855), .B(new_n859), .C1(new_n856), .C2(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n477), .A2(G130), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n462), .A2(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(G142), .B2(new_n474), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n804), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(new_n628), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n858), .A2(new_n870), .A3(new_n860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G162), .B(G160), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n624), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n874), .A3(new_n871), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(G395));
  XNOR2_X1  g455(.A(new_n616), .B(new_n844), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n604), .A2(G299), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n604), .A2(G299), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT41), .B1(new_n883), .B2(new_n884), .ZN(new_n888));
  INV_X1    g463(.A(new_n884), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n882), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G290), .B(G303), .ZN(new_n894));
  XOR2_X1   g469(.A(G288), .B(G305), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(KEYINPUT42), .Z(new_n897));
  AND3_X1   g472(.A1(new_n887), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n887), .B2(new_n893), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g476(.A(new_n900), .B1(G868), .B2(new_n834), .ZN(G331));
  INV_X1    g477(.A(new_n896), .ZN(new_n903));
  NAND2_X1  g478(.A1(G286), .A2(G301), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n536), .A2(new_n537), .A3(new_n540), .A4(new_n544), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n842), .A2(new_n843), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n843), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n562), .B2(new_n841), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(new_n907), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n892), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n911), .B2(new_n907), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n834), .B1(new_n560), .B2(new_n561), .ZN(new_n916));
  OAI211_X1 g491(.A(KEYINPUT104), .B(new_n906), .C1(new_n916), .C2(new_n910), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT105), .B1(new_n911), .B2(new_n907), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  NOR4_X1   g494(.A1(new_n916), .A2(new_n919), .A3(new_n906), .A4(new_n910), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n915), .B(new_n917), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n903), .B(new_n913), .C1(new_n921), .C2(new_n886), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT106), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n908), .A2(new_n919), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n911), .A2(KEYINPUT105), .A3(new_n907), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n926), .A2(new_n885), .A3(new_n915), .A4(new_n917), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n903), .A4(new_n913), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n885), .A2(KEYINPUT107), .A3(new_n890), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n891), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n933), .A3(new_n888), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n921), .A2(new_n934), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n909), .A2(new_n912), .A3(new_n886), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n937), .B2(new_n896), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n930), .A2(KEYINPUT43), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n927), .A2(new_n913), .ZN(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n940), .B2(new_n896), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT43), .B1(new_n930), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n930), .A2(new_n945), .A3(new_n938), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n930), .B2(new_n941), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(G397));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n853), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G40), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n470), .A2(new_n472), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT108), .Z(new_n959));
  INV_X1    g534(.A(G1996), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n732), .B(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n804), .A2(new_n807), .ZN(new_n962));
  INV_X1    g537(.A(G2067), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n703), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n804), .A2(new_n807), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n961), .A2(new_n962), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(G290), .A2(G1986), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n957), .B1(new_n959), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n497), .A2(KEYINPUT100), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n491), .A2(new_n850), .A3(new_n496), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n952), .A2(G1384), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT109), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n970), .A2(new_n975), .A3(new_n971), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n491), .B2(new_n496), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n955), .B1(new_n978), .B2(KEYINPUT45), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(G2072), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n977), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n955), .B1(new_n978), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n497), .A2(new_n984), .A3(new_n950), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n987), .A2(KEYINPUT114), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(KEYINPUT114), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n766), .ZN(new_n991));
  XOR2_X1   g566(.A(G299), .B(KEYINPUT57), .Z(new_n992));
  NAND3_X1  g567(.A1(new_n983), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n983), .B2(new_n991), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(KEYINPUT121), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n979), .B1(new_n974), .B2(new_n976), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n996), .A2(new_n982), .B1(new_n990), .B2(new_n766), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n992), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(KEYINPUT61), .A3(new_n999), .ZN(new_n1000));
  AOI211_X1 g575(.A(KEYINPUT50), .B(G1384), .C1(new_n491), .C2(new_n496), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n768), .B1(new_n985), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n497), .A2(new_n950), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n956), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n963), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1002), .A2(new_n1005), .A3(new_n604), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n604), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT60), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT60), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n605), .A2(new_n1009), .A3(new_n1005), .A4(new_n1002), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT59), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n975), .B1(new_n853), .B2(new_n972), .ZN(new_n1014));
  INV_X1    g589(.A(new_n976), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n980), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(G1996), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(G1341), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1004), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n563), .B(new_n1013), .C1(new_n1017), .C2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n996), .B2(new_n960), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1012), .B(KEYINPUT59), .C1(new_n1022), .C2(new_n562), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1011), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n993), .A2(KEYINPUT118), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n997), .A2(new_n1026), .A3(new_n992), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n994), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1000), .B(new_n1024), .C1(KEYINPUT61), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1007), .B2(new_n994), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n986), .A2(new_n987), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT123), .B(G1961), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI211_X1 g613(.A(G2078), .B(new_n979), .C1(new_n974), .C2(new_n976), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT125), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n707), .B(new_n980), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT125), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n1040), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1038), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT126), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n707), .A2(KEYINPUT53), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n977), .A2(new_n953), .A3(new_n955), .A4(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1046), .A2(new_n1047), .A3(G301), .A4(new_n1049), .ZN(new_n1050));
  AOI211_X1 g625(.A(KEYINPUT125), .B(new_n1041), .C1(new_n996), .C2(new_n707), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1044), .B1(new_n1043), .B2(new_n1040), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1037), .B(new_n1049), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT126), .B1(new_n1053), .B2(G171), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n497), .A2(new_n972), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n979), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1048), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1046), .B2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1034), .B(new_n1050), .C1(new_n1054), .C2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G303), .A2(G8), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT55), .ZN(new_n1061));
  INV_X1    g636(.A(new_n990), .ZN(new_n1062));
  INV_X1    g637(.A(G1971), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1062), .A2(new_n756), .B1(new_n1016), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1966), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n979), .B2(new_n1055), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1069));
  INV_X1    g644(.A(G2084), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n955), .A4(new_n987), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1071), .A3(G168), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G8), .ZN(new_n1073));
  AOI21_X1  g648(.A(G168), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT51), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(G8), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1065), .B1(new_n978), .B2(new_n955), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n579), .A2(new_n581), .A3(G1976), .A4(new_n580), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1079), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1084), .A2(new_n1086), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT111), .B(G1981), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n586), .A2(new_n587), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n791), .B1(new_n586), .B2(new_n587), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT49), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1092), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1094), .B(new_n1095), .C1(KEYINPUT112), .C2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1096), .A2(KEYINPUT112), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT49), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1100), .A3(new_n1080), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1089), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1061), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n996), .A2(G1971), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1035), .A2(G2090), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1103), .B(G8), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1066), .A2(new_n1078), .A3(new_n1102), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1034), .B1(new_n1053), .B2(G171), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1046), .A2(G301), .A3(new_n1057), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1059), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1030), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1033), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(G8), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1061), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1089), .A2(new_n1101), .A3(KEYINPUT113), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT113), .B1(new_n1089), .B2(new_n1101), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(KEYINPUT116), .B(new_n1115), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1122), .A2(new_n1065), .A3(G286), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1106), .A2(KEYINPUT63), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1066), .A2(new_n1102), .A3(new_n1106), .A4(new_n1123), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(KEYINPUT115), .A3(new_n1127), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1125), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1066), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1078), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1075), .A2(new_n1077), .A3(KEYINPUT62), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1133), .A2(new_n1137), .A3(new_n1138), .A4(new_n1058), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1101), .A2(new_n1087), .A3(new_n784), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1080), .B1(new_n1140), .B2(new_n1091), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n1106), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1133), .A2(new_n1137), .A3(new_n1058), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(KEYINPUT127), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1132), .A2(new_n1139), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n969), .B1(new_n1113), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT48), .B1(new_n959), .B2(new_n957), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n959), .A2(KEYINPUT48), .A3(new_n957), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n1148), .B(new_n1149), .C1(new_n957), .C2(new_n966), .ZN(new_n1150));
  INV_X1    g725(.A(new_n964), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n957), .B1(new_n732), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n957), .A2(new_n960), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1153), .A2(KEYINPUT46), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(KEYINPUT46), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT47), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n961), .A2(new_n964), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1158), .A2(new_n965), .B1(G2067), .B2(new_n703), .ZN(new_n1159));
  AOI211_X1 g734(.A(new_n1150), .B(new_n1157), .C1(new_n957), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1147), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g736(.A(G319), .B1(new_n648), .B2(new_n649), .ZN(new_n1163));
  NOR3_X1   g737(.A1(G229), .A2(G227), .A3(new_n1163), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n878), .B(new_n1164), .C1(new_n946), .C2(new_n947), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


