//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G107), .A2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(new_n211), .A2(KEYINPUT66), .B1(G68), .B2(G238), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT65), .Z(new_n214));
  OAI211_X1 g0014(.A(new_n212), .B(new_n214), .C1(KEYINPUT66), .C2(new_n211), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT1), .Z(new_n220));
  OR2_X1    g0020(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n221), .A2(G50), .A3(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n206), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(G257), .A2(G264), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n210), .A3(new_n230), .ZN(new_n231));
  AOI22_X1  g0031(.A1(new_n224), .A2(new_n227), .B1(KEYINPUT0), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n220), .B(new_n232), .C1(KEYINPUT0), .C2(new_n231), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G223), .A2(G1698), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G222), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n256), .B(new_n260), .C1(G77), .C2(new_n252), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT70), .B(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n262), .B(G274), .C1(new_n263), .C2(G45), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n261), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G200), .ZN(new_n269));
  INV_X1    g0069(.A(G190), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n272));
  INV_X1    g0072(.A(G150), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(KEYINPUT8), .A2(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT8), .A2(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n226), .A2(G33), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n272), .B1(new_n273), .B2(new_n275), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n225), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(G50), .B1(new_n226), .B2(G1), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT71), .ZN(new_n285));
  INV_X1    g0085(.A(new_n282), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n283), .B(new_n288), .C1(G50), .C2(new_n287), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n269), .B(new_n271), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT73), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n269), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n289), .B(KEYINPUT9), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(new_n295), .A3(new_n269), .A4(new_n271), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n268), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n268), .A2(G179), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n289), .B(new_n302), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G238), .A2(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(G232), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n252), .B(new_n308), .C1(new_n309), .C2(G1698), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G107), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n310), .A2(new_n260), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n266), .A2(G244), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n264), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n301), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT15), .B(G87), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n278), .A2(new_n275), .B1(new_n321), .B2(new_n279), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n226), .A2(new_n216), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n282), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n226), .A2(G1), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n282), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G77), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n324), .B(new_n327), .C1(G77), .C2(new_n287), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n317), .A2(new_n329), .A3(new_n264), .A4(new_n318), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n320), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n307), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  INV_X1    g0134(.A(G238), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n259), .A2(new_n265), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G226), .A2(G1698), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n309), .B2(G1698), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n338), .A2(new_n252), .B1(G33), .B2(G97), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n264), .B1(new_n335), .B2(new_n336), .C1(new_n339), .C2(new_n259), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n334), .B1(new_n343), .B2(G169), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI211_X1 g0145(.A(KEYINPUT14), .B(new_n301), .C1(new_n341), .C2(new_n342), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n343), .A2(new_n329), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G50), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n275), .A2(new_n351), .B1(new_n279), .B2(new_n216), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n226), .A2(G68), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n282), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  INV_X1    g0155(.A(new_n326), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n354), .A2(new_n355), .B1(new_n202), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n354), .A2(new_n355), .ZN(new_n358));
  INV_X1    g0158(.A(G13), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G1), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n353), .ZN(new_n361));
  XOR2_X1   g0161(.A(new_n361), .B(KEYINPUT12), .Z(new_n362));
  NOR3_X1   g0162(.A1(new_n357), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n350), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n343), .B2(new_n270), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n341), .B2(new_n342), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n333), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n264), .B1(new_n309), .B2(new_n336), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n311), .A2(new_n313), .A3(G223), .A4(new_n254), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT75), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n252), .A2(KEYINPUT75), .A3(G223), .A4(new_n254), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n252), .A2(G226), .A3(G1698), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n372), .B1(new_n260), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(G169), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n329), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n201), .A2(new_n202), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n274), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n252), .B2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n314), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n282), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n314), .B2(new_n226), .ZN(new_n395));
  AOI211_X1 g0195(.A(new_n389), .B(G20), .C1(new_n311), .C2(new_n313), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n388), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT74), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT74), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n393), .A2(new_n402), .A3(KEYINPUT16), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n394), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n287), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n278), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n356), .B2(new_n278), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n382), .B(new_n383), .C1(new_n404), .C2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n286), .B1(new_n399), .B2(new_n400), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n402), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n202), .B1(new_n390), .B2(new_n391), .ZN(new_n413));
  NOR4_X1   g0213(.A1(new_n413), .A2(new_n388), .A3(KEYINPUT74), .A4(new_n400), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n407), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n381), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .A3(new_n383), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n379), .A2(new_n260), .ZN(new_n419));
  INV_X1    g0219(.A(new_n372), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n270), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(G200), .B2(new_n380), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n415), .A2(new_n422), .A3(new_n416), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(new_n416), .A3(new_n422), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT76), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(KEYINPUT17), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n410), .A2(new_n418), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n319), .A2(G200), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n319), .A2(new_n270), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n432), .A2(new_n433), .A3(new_n328), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n371), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n258), .A2(KEYINPUT70), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT70), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G41), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT5), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(G270), .A3(new_n259), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n443), .A2(G274), .A3(new_n444), .A4(new_n446), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n311), .A2(new_n313), .A3(G264), .A4(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT79), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n252), .A2(new_n453), .A3(G264), .A4(G1698), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n252), .A2(G257), .A3(new_n254), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n314), .A2(G303), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n452), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n450), .B1(new_n260), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n262), .A2(G33), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n287), .A2(new_n459), .A3(new_n225), .A4(new_n281), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G116), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n405), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n281), .A2(new_n225), .B1(G20), .B2(new_n463), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  INV_X1    g0266(.A(G97), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n226), .C1(G33), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT20), .B1(new_n465), .B2(new_n468), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n462), .B(new_n464), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n458), .A2(G179), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n450), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n457), .A2(new_n260), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(G190), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n472), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n477), .C1(new_n458), .C2(new_n367), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n458), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n474), .A2(new_n475), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n465), .A2(new_n468), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT20), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(new_n469), .B1(G116), .B2(new_n461), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n301), .B1(new_n486), .B2(new_n464), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(new_n487), .A3(KEYINPUT21), .ZN(new_n488));
  AND4_X1   g0288(.A1(new_n473), .A2(new_n478), .A3(new_n481), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n311), .A2(new_n313), .A3(G244), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(G1698), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n493), .A2(new_n311), .A3(new_n313), .A4(G244), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n492), .A2(new_n466), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n252), .A2(G250), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G1698), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n259), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n447), .A2(G257), .A3(new_n259), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n449), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n301), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n286), .A2(KEYINPUT78), .A3(new_n287), .A4(new_n459), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT78), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n460), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n505), .A3(G97), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n287), .A2(G97), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT77), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n507), .B(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n315), .B1(new_n390), .B2(new_n391), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT6), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n467), .A2(new_n315), .ZN(new_n513));
  NOR2_X1   g0313(.A1(G97), .A2(G107), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n315), .A2(KEYINPUT6), .A3(G97), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n226), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n275), .A2(new_n216), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n511), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n510), .B1(new_n519), .B2(new_n286), .ZN(new_n520));
  INV_X1    g0320(.A(new_n501), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n492), .A2(new_n466), .A3(new_n494), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n254), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n260), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(new_n329), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n502), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n262), .A2(G45), .ZN(new_n527));
  AND2_X1   g0327(.A1(G33), .A2(G41), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(G250), .C1(new_n528), .C2(new_n225), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n446), .A2(G274), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n335), .A2(new_n254), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n217), .A2(G1698), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n252), .B1(G33), .B2(G116), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n532), .B(G190), .C1(new_n536), .C2(new_n259), .ZN(new_n537));
  XOR2_X1   g0337(.A(KEYINPUT15), .B(G87), .Z(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n287), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n209), .A2(new_n467), .A3(new_n315), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G97), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n226), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n542), .A3(KEYINPUT19), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n311), .A2(new_n313), .A3(new_n226), .A4(G68), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n279), .B2(new_n467), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n539), .B1(new_n547), .B2(new_n282), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n503), .A2(new_n505), .A3(G87), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n537), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G116), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n533), .A2(new_n534), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n314), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n531), .B1(new_n553), .B2(new_n260), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n503), .A2(new_n505), .A3(new_n538), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n548), .B1(new_n554), .B2(new_n329), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(new_n301), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n550), .A2(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(G200), .B1(new_n499), .B2(new_n501), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n506), .A2(new_n509), .ZN(new_n562));
  OAI21_X1  g0362(.A(G107), .B1(new_n395), .B2(new_n396), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n515), .A2(new_n516), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G20), .ZN(new_n565));
  INV_X1    g0365(.A(new_n518), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n562), .B1(new_n567), .B2(new_n282), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n521), .A2(G190), .A3(new_n524), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n561), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n526), .A2(new_n560), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n311), .A2(new_n313), .A3(G257), .A4(G1698), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n311), .A2(new_n313), .A3(G250), .A4(new_n254), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G294), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n260), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n447), .A2(G264), .A3(new_n259), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT82), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT82), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n579), .A2(G179), .A3(new_n449), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n576), .A2(new_n577), .A3(new_n449), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G169), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n311), .A2(new_n313), .A3(new_n226), .A4(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT22), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT22), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n252), .A2(new_n588), .A3(new_n226), .A4(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OR3_X1    g0390(.A1(new_n551), .A2(KEYINPUT80), .A3(G20), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT80), .B1(new_n551), .B2(G20), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n226), .B2(G107), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n315), .A2(KEYINPUT23), .A3(G20), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n591), .A2(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n590), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n599), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n590), .A2(new_n596), .A3(new_n597), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n282), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n360), .A2(G20), .A3(new_n315), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n604), .A2(KEYINPUT25), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n503), .A2(new_n505), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G107), .B1(KEYINPUT25), .B2(new_n604), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n585), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n580), .B1(new_n576), .B2(new_n577), .ZN(new_n611));
  INV_X1    g0411(.A(new_n449), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n613), .A2(G200), .B1(G190), .B2(new_n583), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n489), .A2(new_n571), .A3(new_n609), .A4(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n438), .A2(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n306), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n364), .A2(new_n350), .B1(new_n370), .B2(new_n332), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n430), .A2(new_n425), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT18), .B1(new_n417), .B2(new_n383), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n408), .A2(new_n409), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n620), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n625), .B2(new_n300), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n502), .A2(new_n520), .A3(new_n525), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT83), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n529), .A2(new_n629), .A3(new_n530), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n529), .B2(new_n530), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n630), .A2(new_n631), .B1(new_n536), .B2(new_n259), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G200), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n301), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n550), .A2(new_n633), .B1(new_n558), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n627), .A2(new_n628), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n550), .A2(new_n556), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n558), .A2(new_n559), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT26), .B1(new_n639), .B2(new_n526), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n558), .A2(new_n634), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n636), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT84), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n609), .A2(new_n473), .A3(new_n481), .A4(new_n488), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n526), .A2(new_n635), .A3(new_n570), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n616), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n636), .A2(new_n640), .A3(new_n647), .A4(new_n641), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n643), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n626), .B1(new_n438), .B2(new_n650), .ZN(G369));
  NOR2_X1   g0451(.A1(new_n359), .A2(G20), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n262), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n608), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n616), .A2(new_n609), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n585), .A2(new_n608), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT85), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n481), .A2(new_n473), .A3(new_n488), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n658), .A2(new_n472), .ZN(new_n668));
  MUX2_X1   g0468(.A(new_n667), .B(new_n489), .S(new_n668), .Z(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n658), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n663), .B2(new_n665), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n585), .A2(new_n608), .A3(new_n673), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(G399));
  NOR2_X1   g0479(.A1(new_n229), .A2(new_n263), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G1), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n540), .A2(G116), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n223), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n645), .A2(new_n616), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n667), .B1(new_n585), .B2(new_n608), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT89), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n627), .A2(KEYINPUT26), .A3(new_n635), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT88), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n628), .B1(new_n639), .B2(new_n526), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n627), .A2(KEYINPUT88), .A3(KEYINPUT26), .A4(new_n635), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n644), .A2(new_n695), .A3(new_n616), .A4(new_n645), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n688), .A2(new_n641), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n697), .A2(KEYINPUT90), .A3(new_n673), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT90), .B1(new_n697), .B2(new_n673), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT29), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n649), .A2(new_n673), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT87), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT87), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(new_n705), .A3(new_n702), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n700), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n579), .A2(new_n581), .A3(new_n524), .A4(new_n521), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n474), .A2(G179), .A3(new_n475), .A4(new_n554), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n579), .A2(new_n449), .A3(new_n581), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n521), .A2(new_n524), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n632), .A2(new_n329), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n712), .A2(new_n482), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT86), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n711), .A2(KEYINPUT86), .A3(new_n715), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n709), .A2(new_n710), .A3(new_n708), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT31), .B(new_n658), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n616), .A2(new_n609), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n489), .A3(new_n571), .A4(new_n673), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n658), .B1(new_n716), .B2(new_n721), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n707), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n685), .B1(new_n730), .B2(G1), .ZN(G364));
  INV_X1    g0531(.A(new_n670), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n652), .A2(G45), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n681), .A2(G1), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n669), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n226), .A2(new_n270), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n329), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n252), .B1(new_n741), .B2(G322), .ZN(new_n742));
  INV_X1    g0542(.A(G329), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n226), .A2(G190), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n742), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n226), .B1(new_n745), .B2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(G294), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n329), .A2(new_n367), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n738), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G326), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n367), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n744), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n738), .A2(new_n755), .ZN(new_n759));
  INV_X1    g0559(.A(G303), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n744), .A2(new_n739), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n759), .A2(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n751), .A2(new_n744), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT33), .B(G317), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n758), .B(new_n763), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n750), .A2(new_n754), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n746), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G159), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G97), .B2(new_n749), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n314), .B1(new_n741), .B2(G58), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n761), .A2(KEYINPUT91), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n761), .A2(KEYINPUT91), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G77), .ZN(new_n778));
  INV_X1    g0578(.A(new_n759), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G87), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n351), .B2(new_n752), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G68), .B2(new_n765), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n772), .A2(new_n773), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n756), .A2(new_n315), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n768), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n225), .B1(G20), .B2(new_n301), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n786), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n224), .A2(new_n445), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n229), .A2(new_n252), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(new_n445), .C2(new_n247), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n229), .A2(new_n314), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G355), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G116), .C2(new_n228), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n785), .A2(new_n786), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n789), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n669), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n737), .B1(new_n734), .B2(new_n799), .ZN(G396));
  AOI21_X1  g0600(.A(new_n314), .B1(new_n769), .B2(G132), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n801), .B1(new_n351), .B2(new_n759), .C1(new_n201), .C2(new_n748), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G137), .A2(new_n753), .B1(new_n741), .B2(G143), .ZN(new_n803));
  INV_X1    g0603(.A(G159), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n273), .B2(new_n764), .C1(new_n776), .C2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT34), .Z(new_n806));
  INV_X1    g0606(.A(new_n756), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n802), .B(new_n806), .C1(G68), .C2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G303), .A2(new_n753), .B1(new_n807), .B2(G87), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n776), .B2(new_n463), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n314), .B1(new_n746), .B2(new_n762), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G107), .B2(new_n779), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(new_n467), .B2(new_n748), .C1(new_n757), .C2(new_n764), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n810), .B(new_n813), .C1(G294), .C2(new_n741), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n786), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n786), .A2(new_n787), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n734), .B1(new_n216), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT92), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n328), .A2(new_n658), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT93), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n331), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n320), .A2(new_n328), .A3(KEYINPUT93), .A4(new_n330), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n435), .B(new_n819), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n331), .A2(new_n673), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n815), .B(new_n818), .C1(new_n788), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n434), .B1(new_n821), .B2(new_n823), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n701), .A2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(KEYINPUT94), .B(new_n826), .C1(new_n830), .C2(new_n819), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT94), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n825), .B2(new_n827), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n832), .B1(new_n701), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(new_n729), .Z(new_n839));
  OAI21_X1  g0639(.A(new_n829), .B1(new_n839), .B2(new_n735), .ZN(G384));
  OAI21_X1  g0640(.A(new_n621), .B1(new_n624), .B2(new_n623), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n415), .A2(new_n416), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n656), .B(KEYINPUT96), .Z(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n408), .A3(new_n426), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n844), .A2(new_n408), .A3(new_n849), .A4(new_n426), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n656), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n404), .B2(new_n407), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n408), .A2(new_n426), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(new_n850), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT95), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n431), .B2(new_n854), .ZN(new_n859));
  INV_X1    g0659(.A(new_n854), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n841), .A2(KEYINPUT95), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n857), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n852), .B1(new_n862), .B2(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n726), .A2(KEYINPUT98), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n658), .B(new_n864), .C1(new_n716), .C2(new_n721), .ZN(new_n865));
  INV_X1    g0665(.A(new_n864), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n725), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n724), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n364), .B(new_n658), .C1(new_n350), .C2(new_n369), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n364), .A2(new_n658), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n370), .B(new_n870), .C1(new_n871), .C2(new_n363), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n868), .A2(new_n873), .A3(new_n828), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT40), .B1(new_n863), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT40), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n868), .A2(new_n873), .A3(new_n876), .A4(new_n828), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n879), .B(new_n857), .C1(new_n859), .C2(new_n861), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n859), .A2(new_n861), .ZN(new_n881));
  INV_X1    g0681(.A(new_n857), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n878), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n437), .A2(new_n868), .ZN(new_n886));
  XOR2_X1   g0686(.A(new_n885), .B(new_n886), .Z(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(G330), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n700), .A2(new_n437), .A3(new_n704), .A4(new_n706), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n626), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT97), .Z(new_n891));
  XNOR2_X1  g0691(.A(new_n888), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n881), .A2(new_n882), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n879), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n880), .B2(new_n852), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n365), .A2(new_n658), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n624), .A2(new_n623), .A3(new_n843), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n822), .A2(new_n824), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n673), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n701), .B2(new_n831), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(new_n873), .C1(new_n880), .C2(new_n883), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n892), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n262), .B2(new_n652), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n463), .B1(new_n564), .B2(KEYINPUT35), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n909), .B(new_n227), .C1(KEYINPUT35), .C2(new_n564), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT36), .ZN(new_n911));
  OAI21_X1  g0711(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n223), .A2(new_n912), .B1(G50), .B2(new_n202), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(G1), .A3(new_n359), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n908), .A2(new_n911), .A3(new_n914), .ZN(G367));
  OAI211_X1 g0715(.A(new_n526), .B(new_n570), .C1(new_n568), .C2(new_n673), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(new_n609), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n658), .B1(new_n917), .B2(new_n526), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT42), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n627), .A2(new_n658), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n919), .B1(new_n676), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n662), .B(KEYINPUT85), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n924), .A2(KEYINPUT42), .A3(new_n675), .A4(new_n921), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n918), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n548), .A2(new_n549), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n635), .B1(new_n928), .B2(new_n673), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT99), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n641), .A2(new_n928), .A3(new_n673), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(KEYINPUT99), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT100), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT43), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n926), .A2(new_n935), .A3(KEYINPUT43), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n927), .B(new_n934), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n671), .A2(new_n921), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n938), .ZN(new_n942));
  INV_X1    g0742(.A(new_n934), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n936), .A3(new_n943), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n939), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n941), .B1(new_n939), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n680), .B(KEYINPUT41), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT103), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n676), .A2(new_n677), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n922), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT44), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n951), .A2(new_n950), .A3(new_n922), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI211_X1 g0756(.A(KEYINPUT103), .B(new_n921), .C1(new_n676), .C2(new_n677), .ZN(new_n957));
  OAI21_X1  g0757(.A(KEYINPUT44), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n676), .A2(new_n677), .A3(new_n921), .ZN(new_n960));
  XNOR2_X1  g0760(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n960), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT45), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n965), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(new_n968), .A3(new_n963), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n671), .B1(new_n959), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n956), .A2(new_n958), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n972), .A2(new_n672), .A3(new_n969), .A4(new_n966), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n676), .A2(KEYINPUT104), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n732), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n670), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n924), .A2(new_n675), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n977), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n730), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n971), .A2(new_n973), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n949), .B1(new_n983), .B2(new_n730), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n733), .A2(G1), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n947), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n314), .B1(new_n748), .B2(new_n315), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n759), .A2(new_n463), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT46), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(G311), .C2(new_n753), .ZN(new_n990));
  INV_X1    g0790(.A(G294), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n991), .A2(new_n764), .B1(new_n740), .B2(new_n760), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n756), .A2(new_n467), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n777), .C2(G283), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n990), .B(new_n994), .C1(new_n995), .C2(new_n746), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n756), .A2(new_n216), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n748), .A2(new_n202), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n252), .B1(new_n764), .B2(new_n804), .C1(new_n273), .C2(new_n740), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G143), .C2(new_n753), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G58), .A2(new_n779), .B1(new_n769), .B2(G137), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n351), .C2(new_n776), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n996), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n786), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n792), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n790), .B1(new_n228), .B2(new_n321), .C1(new_n243), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n735), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT105), .Z(new_n1009));
  OAI211_X1 g0809(.A(new_n1005), .B(new_n1009), .C1(new_n798), .C2(new_n934), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n986), .A2(KEYINPUT106), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT106), .B1(new_n986), .B2(new_n1010), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(KEYINPUT107), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n982), .B2(new_n681), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n981), .A2(KEYINPUT107), .A3(new_n680), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n730), .C2(new_n980), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n980), .A2(new_n985), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G322), .A2(new_n753), .B1(new_n765), .B2(G311), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n995), .B2(new_n740), .C1(new_n776), .C2(new_n760), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n757), .B2(new_n748), .C1(new_n991), .C2(new_n759), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT49), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n769), .A2(G326), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n252), .B1(new_n807), .B2(G116), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n764), .A2(new_n278), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n779), .A2(G77), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n761), .B2(new_n202), .C1(new_n273), .C2(new_n746), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G159), .B2(new_n753), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n314), .B(new_n993), .C1(G50), .C2(new_n741), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n321), .C2(new_n748), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1030), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1006), .B1(new_n240), .B2(G45), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n683), .B2(new_n794), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n278), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n351), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n683), .B1(new_n1041), .B2(KEYINPUT50), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1042), .B(new_n445), .C1(KEYINPUT50), .C2(new_n1041), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G68), .B2(G77), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1039), .A2(new_n1044), .B1(G107), .B2(new_n228), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1037), .A2(new_n786), .B1(new_n790), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n735), .C1(new_n924), .C2(new_n798), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1019), .A2(new_n1020), .A3(new_n1047), .ZN(G393));
  NAND2_X1  g0848(.A1(new_n971), .A2(new_n973), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n981), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(new_n680), .A3(new_n983), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n971), .A2(new_n985), .A3(new_n973), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G50), .A2(new_n765), .B1(new_n769), .B2(G143), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n202), .B2(new_n759), .C1(new_n209), .C2(new_n756), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n748), .A2(new_n216), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(new_n314), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n752), .A2(new_n273), .B1(new_n740), .B2(new_n804), .ZN(new_n1057));
  XOR2_X1   g0857(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n1058));
  XNOR2_X1  g0858(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1056), .B(new_n1059), .C1(new_n278), .C2(new_n776), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT109), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G303), .A2(new_n765), .B1(new_n769), .B2(G322), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n757), .B2(new_n759), .C1(new_n991), .C2(new_n761), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G116), .B2(new_n749), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n752), .A2(new_n995), .B1(new_n740), .B2(new_n762), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n314), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1061), .B1(new_n784), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n734), .B1(new_n1068), .B2(new_n786), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n790), .B1(new_n467), .B2(new_n228), .C1(new_n250), .C2(new_n1006), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n798), .C2(new_n921), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1051), .A2(new_n1052), .A3(new_n1071), .ZN(G390));
  AND4_X1   g0872(.A1(G330), .A2(new_n728), .A3(new_n828), .A4(new_n873), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT111), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n865), .B1(new_n617), .B2(new_n658), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n867), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n836), .B(G330), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n873), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n828), .B1(new_n698), .B2(new_n699), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1077), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1080), .A2(new_n903), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n874), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n728), .A2(G330), .A3(new_n828), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1084), .A2(G330), .B1(new_n1085), .B2(new_n1078), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n904), .ZN(new_n1087));
  OAI21_X1  g0887(.A(KEYINPUT110), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT110), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1085), .A2(new_n1078), .ZN(new_n1090));
  INV_X1    g0890(.A(G330), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n874), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1089), .B(new_n904), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1083), .A2(new_n1088), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n886), .A2(G330), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n889), .A2(new_n1095), .A3(new_n626), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n880), .A2(new_n852), .B1(new_n365), .B2(new_n658), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1081), .A2(new_n903), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n873), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n899), .B1(new_n904), .B2(new_n873), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n896), .B2(new_n898), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1100), .A2(new_n1102), .A3(new_n1073), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1092), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n863), .A2(new_n899), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n903), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n697), .A2(new_n673), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT90), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n697), .A2(KEYINPUT90), .A3(new_n673), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1106), .B1(new_n1111), .B2(new_n828), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1105), .B1(new_n1112), .B2(new_n1078), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1101), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n880), .A2(new_n883), .A3(new_n897), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1104), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1097), .B1(new_n1103), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1092), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1073), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1113), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1120), .A2(new_n1122), .A3(new_n1096), .A4(new_n1094), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1119), .A2(new_n680), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(KEYINPUT112), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT112), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1119), .A2(new_n1126), .A3(new_n1123), .A4(new_n680), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1120), .A2(new_n1122), .A3(new_n985), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n787), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n816), .A2(new_n278), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n777), .A2(G97), .B1(G283), .B2(new_n753), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n315), .B2(new_n764), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT113), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n740), .A2(new_n463), .B1(new_n756), .B2(new_n202), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1055), .B(new_n1135), .C1(G294), .C2(new_n769), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1134), .A2(new_n314), .A3(new_n780), .A4(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G128), .A2(new_n753), .B1(new_n807), .B2(G50), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n769), .A2(G125), .ZN(new_n1139));
  INV_X1    g0939(.A(G132), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1138), .B(new_n1139), .C1(new_n1140), .C2(new_n740), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n314), .B(new_n1141), .C1(G159), .C2(new_n749), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT54), .B(G143), .Z(new_n1143));
  NAND2_X1  g0943(.A1(new_n777), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n765), .A2(G137), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n779), .A2(G150), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1137), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT114), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n734), .B1(new_n1150), .B2(new_n786), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1130), .A2(new_n1131), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1129), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1128), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT115), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT115), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1128), .A2(new_n1157), .A3(new_n1154), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(G378));
  NAND2_X1  g0959(.A1(new_n1123), .A2(new_n1096), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n289), .A2(new_n853), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT55), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n300), .B2(new_n306), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n300), .A2(new_n1164), .A3(new_n306), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1163), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1163), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1169), .A2(new_n1165), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1162), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1169), .B2(new_n1165), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1166), .A2(new_n1167), .A3(new_n1163), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(new_n1161), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n885), .B2(G330), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1091), .B(new_n1176), .C1(new_n875), .C2(new_n884), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n906), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n852), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n895), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n876), .B1(new_n1182), .B2(new_n1084), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n877), .B1(new_n894), .B2(new_n895), .ZN(new_n1184));
  OAI21_X1  g0984(.A(G330), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1176), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n885), .A2(G330), .A3(new_n1177), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT119), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1180), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n906), .B(KEYINPUT119), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1160), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1123), .A2(new_n1096), .B1(new_n1180), .B2(new_n1189), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n681), .B1(new_n1196), .B2(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1191), .A2(new_n985), .A3(new_n1192), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1177), .A2(new_n787), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n816), .A2(new_n351), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n753), .A2(G116), .B1(new_n769), .B2(G283), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n467), .B2(new_n764), .C1(new_n315), .C2(new_n740), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n756), .A2(new_n201), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n252), .A2(new_n263), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1032), .B(new_n1205), .C1(new_n321), .C2(new_n761), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1203), .A2(new_n998), .A3(new_n1204), .A4(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT58), .Z(new_n1208));
  INV_X1    g1008(.A(new_n761), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n779), .A2(new_n1143), .B1(new_n1209), .B2(G137), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n741), .A2(G128), .B1(new_n749), .B2(G150), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n753), .A2(G125), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n765), .A2(G132), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n807), .A2(G159), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT117), .B(G124), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G33), .B(G41), .C1(new_n769), .C2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n351), .B1(G33), .B2(G41), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1208), .B(new_n1221), .C1(new_n1205), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n734), .B1(new_n1223), .B2(new_n786), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1200), .A2(new_n1201), .A3(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1199), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1198), .A2(new_n1226), .ZN(G375));
  NOR2_X1   g1027(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT120), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n948), .A3(new_n1097), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT121), .Z(new_n1231));
  NAND2_X1  g1031(.A1(new_n1094), .A2(new_n985), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n873), .A2(new_n788), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT122), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n816), .A2(new_n202), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(KEYINPUT122), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n748), .A2(new_n321), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n314), .B1(new_n746), .B2(new_n760), .C1(new_n216), .C2(new_n756), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(G97), .C2(new_n779), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n463), .A2(new_n764), .B1(new_n740), .B2(new_n757), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n777), .B2(G107), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(new_n991), .C2(new_n752), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n752), .A2(new_n1140), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT123), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G50), .B2(new_n749), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n741), .A2(G137), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n765), .A2(new_n1143), .B1(new_n769), .B2(G128), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n314), .B(new_n1204), .C1(G150), .C2(new_n1209), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n759), .A2(new_n804), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1243), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT124), .Z(new_n1253));
  AOI21_X1  g1053(.A(new_n734), .B1(new_n1253), .B2(new_n786), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1232), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1231), .A2(new_n1257), .ZN(G381));
  INV_X1    g1058(.A(G390), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1012), .A2(new_n1014), .A3(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1260), .A2(G381), .A3(G384), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1262), .B(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1124), .A2(new_n1154), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(G375), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1264), .A2(new_n1267), .ZN(G407));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n657), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G213), .B(new_n1269), .C1(new_n1264), .C2(new_n1267), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n657), .A2(G213), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1097), .A2(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1229), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n680), .A3(new_n1275), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1276), .A2(G384), .A3(new_n1257), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1276), .B2(new_n1257), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G375), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1193), .A2(new_n949), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1225), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1180), .A2(new_n1189), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n985), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1265), .B1(new_n1281), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1272), .B(new_n1279), .C1(new_n1280), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G393), .B(G396), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1011), .A2(new_n1013), .A3(G390), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n986), .A2(new_n1010), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(G390), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1289), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1291), .A2(G390), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1289), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1292), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1157), .B1(new_n1128), .B2(new_n1154), .ZN(new_n1299));
  AOI211_X1 g1099(.A(KEYINPUT115), .B(new_n1153), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1198), .B(new_n1226), .C1(new_n1299), .C2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1285), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1272), .A4(new_n1279), .ZN(new_n1304));
  AND4_X1   g1104(.A1(new_n1271), .A2(new_n1288), .A3(new_n1298), .A4(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1272), .B1(new_n1280), .B2(new_n1285), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1303), .A2(KEYINPUT126), .A3(new_n1272), .ZN(new_n1309));
  INV_X1    g1109(.A(G2897), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1272), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1279), .A2(new_n1311), .ZN(new_n1312));
  OAI22_X1  g1112(.A1(new_n1277), .A2(new_n1278), .B1(new_n1310), .B2(new_n1272), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1308), .A2(new_n1309), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT127), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1308), .A2(new_n1309), .A3(KEYINPUT127), .A4(new_n1314), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1305), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT61), .B1(new_n1286), .B2(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1314), .A2(new_n1306), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1320), .B(new_n1321), .C1(KEYINPUT62), .C2(new_n1286), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1298), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1319), .A2(new_n1324), .ZN(G405));
  AOI21_X1  g1125(.A(new_n1265), .B1(new_n1198), .B2(new_n1226), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1301), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1279), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(new_n1323), .ZN(G402));
endmodule


