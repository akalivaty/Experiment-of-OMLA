//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G141gat), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT80), .B(G141gat), .Z(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(new_n203), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n211), .A2(KEYINPUT81), .B1(KEYINPUT2), .B2(new_n210), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n206), .B(new_n212), .C1(KEYINPUT81), .C2(new_n211), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n210), .B1(KEYINPUT79), .B2(KEYINPUT2), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n217));
  OAI22_X1  g016(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n214), .A2(new_n215), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n210), .B(new_n209), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G211gat), .B(G218gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224));
  INV_X1    g023(.A(G211gat), .ZN(new_n225));
  INV_X1    g024(.A(G218gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n222), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT75), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n222), .A2(KEYINPUT74), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n223), .A2(new_n227), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(KEYINPUT74), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT29), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n221), .B1(new_n234), .B2(KEYINPUT3), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT85), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g036(.A(KEYINPUT85), .B(new_n221), .C1(new_n234), .C2(KEYINPUT3), .ZN(new_n238));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n229), .A2(new_n233), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n213), .A2(new_n220), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n239), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n237), .A2(new_n238), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n221), .ZN(new_n248));
  INV_X1    g047(.A(new_n231), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n249), .A2(new_n222), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n229), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n244), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n248), .B1(new_n252), .B2(new_n242), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n240), .B1(new_n244), .B2(new_n243), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n239), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n202), .B1(new_n256), .B2(G22gat), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G50gat), .ZN(new_n259));
  XOR2_X1   g058(.A(G78gat), .B(G106gat), .Z(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G22gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n263), .B1(new_n247), .B2(new_n255), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n247), .A2(new_n255), .A3(new_n263), .ZN(new_n265));
  OAI22_X1  g064(.A1(new_n257), .A2(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n264), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n255), .A3(new_n263), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(new_n202), .A3(new_n268), .A4(new_n261), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G113gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(G120gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(new_n271), .B2(G120gat), .ZN(new_n275));
  INV_X1    g074(.A(G120gat), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n273), .B(new_n275), .C1(G113gat), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n276), .A2(G113gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n272), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n279), .A2(new_n283), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G183gat), .B2(G190gat), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT64), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n291), .ZN(new_n293));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .A4(new_n289), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(KEYINPUT23), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n302), .A2(new_n303), .B1(new_n298), .B2(KEYINPUT23), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n292), .A2(new_n297), .A3(new_n299), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT25), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n299), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n294), .B1(new_n311), .B2(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n313), .A2(KEYINPUT68), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT68), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n312), .B(KEYINPUT69), .C1(new_n315), .C2(new_n316), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n310), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n308), .A2(new_n309), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT27), .B(G183gat), .ZN(new_n323));
  INV_X1    g122(.A(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n325), .B(KEYINPUT28), .Z(new_n326));
  NAND2_X1  g125(.A1(new_n302), .A2(new_n303), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  OR3_X1    g127(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n313), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n288), .B1(new_n322), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G227gat), .ZN(new_n334));
  INV_X1    g133(.A(G233gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n305), .A2(new_n307), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT67), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n304), .A2(new_n299), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n291), .B(KEYINPUT68), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT69), .B1(new_n340), .B2(new_n312), .ZN(new_n341));
  INV_X1    g140(.A(new_n320), .ZN(new_n342));
  OAI211_X1 g141(.A(KEYINPUT25), .B(new_n339), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(new_n287), .A3(new_n331), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n333), .A2(new_n336), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT72), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT72), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n333), .A2(new_n349), .A3(new_n336), .A4(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G15gat), .B(G43gat), .Z(new_n355));
  XNOR2_X1  g154(.A(G71gat), .B(G99gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n333), .A2(new_n346), .ZN(new_n359));
  INV_X1    g158(.A(new_n336), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n361), .A2(KEYINPUT34), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(KEYINPUT34), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT32), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n348), .B2(new_n350), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT33), .B1(new_n348), .B2(new_n350), .ZN(new_n367));
  INV_X1    g166(.A(new_n357), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n358), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n270), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n345), .B2(new_n331), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(KEYINPUT76), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n345), .A2(new_n331), .ZN(new_n379));
  INV_X1    g178(.A(new_n376), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n345), .B2(new_n331), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n383), .B2(KEYINPUT76), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(new_n240), .ZN(new_n385));
  INV_X1    g184(.A(new_n382), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(KEYINPUT77), .A3(new_n376), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n382), .B2(new_n380), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n387), .A2(new_n389), .A3(new_n240), .A4(new_n381), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n375), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n390), .B(new_n374), .C1(new_n384), .C2(new_n240), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(KEYINPUT30), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n383), .A2(KEYINPUT76), .ZN(new_n395));
  INV_X1    g194(.A(new_n378), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n241), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n390), .A4(new_n374), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n213), .A2(new_n220), .A3(new_n286), .A4(new_n280), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(new_n243), .A3(new_n287), .ZN(new_n405));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n403), .A2(new_n405), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n409), .A2(KEYINPUT5), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n221), .A2(new_n287), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n401), .ZN(new_n412));
  INV_X1    g211(.A(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT5), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n406), .B1(new_n411), .B2(new_n401), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT83), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n416), .B(new_n419), .C1(new_n409), .C2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n409), .A2(new_n420), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n410), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n428), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n410), .B(new_n427), .C1(new_n421), .C2(new_n422), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n394), .A2(new_n400), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n364), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n436));
  AOI221_X4 g235(.A(new_n365), .B1(KEYINPUT33), .B2(new_n357), .C1(new_n348), .C2(new_n350), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n364), .B1(new_n358), .B2(new_n369), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT73), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n371), .A2(new_n434), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT35), .ZN(new_n444));
  INV_X1    g243(.A(new_n270), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(KEYINPUT35), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT91), .ZN(new_n447));
  INV_X1    g246(.A(new_n370), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(new_n441), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n438), .A2(KEYINPUT91), .A3(new_n370), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n446), .A2(new_n449), .A3(new_n434), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT39), .B1(new_n412), .B2(new_n413), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n453), .A2(KEYINPUT88), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(KEYINPUT88), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n403), .A2(new_n405), .A3(new_n408), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n413), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n457), .A2(KEYINPUT39), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT40), .A4(new_n427), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n460), .B(KEYINPUT89), .Z(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n459), .A3(new_n427), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n462), .A2(new_n463), .B1(new_n423), .B2(new_n428), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n461), .A2(new_n394), .A3(new_n400), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n398), .A2(new_n466), .A3(new_n467), .A4(new_n390), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n390), .B(new_n467), .C1(new_n384), .C2(new_n240), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT90), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n467), .B1(new_n397), .B2(new_n240), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n387), .A2(new_n389), .A3(new_n241), .A4(new_n381), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT38), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n375), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n433), .A2(new_n429), .A3(new_n393), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n374), .B1(new_n468), .B2(new_n470), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT37), .B1(new_n385), .B2(new_n391), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n465), .B(new_n270), .C1(new_n477), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n394), .A2(new_n400), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n433), .A2(new_n429), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n270), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n370), .A2(KEYINPUT36), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n440), .A3(new_n442), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT36), .B1(new_n438), .B2(new_n370), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n485), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT87), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n482), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g291(.A(KEYINPUT87), .B(new_n485), .C1(new_n487), .C2(new_n489), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n452), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n495));
  INV_X1    g294(.A(G36gat), .ZN(new_n496));
  AND2_X1   g295(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G29gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n504));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n504), .A2(new_n505), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT17), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G1gat), .B2(new_n510), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n513), .A2(G8gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(G8gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT93), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n516), .A2(KEYINPUT93), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n509), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n508), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT18), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n508), .B(new_n516), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n520), .B(KEYINPUT13), .Z(new_n525));
  AOI22_X1  g324(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n519), .A2(KEYINPUT18), .A3(new_n520), .A4(new_n521), .ZN(new_n527));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G169gat), .B(G197gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT12), .Z(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n526), .A2(new_n527), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n526), .B2(new_n527), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n495), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n526), .A2(new_n527), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n533), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n526), .A2(new_n527), .A3(new_n534), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(KEYINPUT94), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n494), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G71gat), .B(G78gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT21), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G127gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n515), .B(new_n514), .C1(new_n550), .C2(new_n551), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT95), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(new_n207), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n560), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n558), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT41), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT96), .ZN(new_n568));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT97), .B(G85gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT98), .B(G92gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT7), .ZN(new_n575));
  INV_X1    g374(.A(G99gat), .ZN(new_n576));
  INV_X1    g375(.A(G106gat), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT8), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n508), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n566), .B2(new_n565), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n579), .B(new_n580), .Z(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n509), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n570), .B1(new_n588), .B2(KEYINPUT99), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n585), .B(new_n587), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n564), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n584), .A2(new_n550), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n549), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n549), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n602), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n596), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(KEYINPUT100), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n596), .B1(new_n598), .B2(new_n600), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  OR4_X1    g412(.A1(new_n605), .A2(new_n608), .A3(new_n609), .A4(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n613), .B1(new_n603), .B2(new_n609), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT101), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n595), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n544), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n484), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G1gat), .ZN(G1324gat));
  INV_X1    g422(.A(new_n483), .ZN(new_n624));
  INV_X1    g423(.A(new_n619), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n494), .A2(new_n624), .A3(new_n543), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT102), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n358), .A2(new_n369), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT73), .B1(new_n628), .B2(new_n435), .ZN(new_n629));
  AOI211_X1 g428(.A(new_n439), .B(new_n364), .C1(new_n358), .C2(new_n369), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n488), .B1(new_n631), .B2(new_n486), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT87), .B1(new_n632), .B2(new_n485), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n487), .A2(new_n489), .ZN(new_n634));
  INV_X1    g433(.A(new_n485), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n491), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n636), .A3(new_n482), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n542), .B1(new_n637), .B2(new_n452), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n624), .A4(new_n625), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n627), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT103), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n627), .A2(new_n640), .A3(G8gat), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n620), .A2(KEYINPUT42), .A3(new_n624), .A4(new_n643), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n649), .A3(KEYINPUT104), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT42), .B1(new_n641), .B2(new_n643), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n648), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(G1325gat));
  INV_X1    g454(.A(new_n620), .ZN(new_n656));
  OAI21_X1  g455(.A(G15gat), .B1(new_n656), .B2(new_n634), .ZN(new_n657));
  INV_X1    g456(.A(G15gat), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n449), .A2(new_n450), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n620), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(G1326gat));
  OAI21_X1  g460(.A(KEYINPUT105), .B1(new_n656), .B2(new_n270), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n620), .A2(new_n663), .A3(new_n445), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n662), .B2(new_n664), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(G1327gat));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n485), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT106), .B1(new_n434), .B2(new_n270), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n482), .A2(new_n634), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n452), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n594), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n494), .A2(KEYINPUT44), .A3(new_n594), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n564), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n539), .A2(new_n540), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n679), .A2(new_n681), .A3(new_n617), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT107), .B1(new_n683), .B2(new_n484), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n678), .A2(new_n685), .A3(new_n621), .A4(new_n682), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(G29gat), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n679), .A2(new_n617), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n594), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n544), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n500), .A3(new_n621), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT45), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(new_n692), .ZN(G1328gat));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n496), .A3(new_n624), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT46), .Z(new_n695));
  OAI21_X1  g494(.A(G36gat), .B1(new_n683), .B2(new_n483), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(G1329gat));
  NAND4_X1  g496(.A1(new_n678), .A2(G43gat), .A3(new_n632), .A4(new_n682), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT47), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(KEYINPUT108), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n638), .A2(new_n659), .A3(new_n594), .A4(new_n688), .ZN(new_n701));
  INV_X1    g500(.A(G43gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(KEYINPUT108), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT109), .Z(new_n705));
  AND3_X1   g504(.A1(new_n698), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n698), .B2(new_n703), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(G1330gat));
  NAND4_X1  g507(.A1(new_n676), .A2(new_n677), .A3(new_n445), .A4(new_n682), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G50gat), .ZN(new_n710));
  INV_X1    g509(.A(G50gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n690), .A2(new_n711), .A3(new_n445), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT48), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716));
  AOI211_X1 g515(.A(KEYINPUT110), .B(new_n716), .C1(new_n710), .C2(new_n712), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n715), .A2(new_n717), .ZN(G1331gat));
  NOR4_X1   g517(.A1(new_n564), .A2(new_n618), .A3(new_n594), .A4(new_n680), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n673), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n621), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g522(.A1(new_n720), .A2(new_n483), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n720), .B2(new_n634), .ZN(new_n729));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n659), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n720), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g532(.A1(new_n720), .A2(new_n270), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT111), .B(G78gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1335gat));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n679), .A2(new_n680), .A3(new_n618), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n676), .A2(new_n677), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(new_n484), .ZN(new_n741));
  INV_X1    g540(.A(new_n571), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n739), .A2(KEYINPUT112), .A3(new_n621), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n679), .A2(new_n680), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n674), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n673), .A2(KEYINPUT51), .A3(new_n594), .A4(new_n746), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n750), .A2(new_n621), .A3(new_n571), .A4(new_n617), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n744), .A2(new_n751), .ZN(G1336gat));
  NOR3_X1   g551(.A1(new_n483), .A2(new_n618), .A3(G92gat), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT113), .Z(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n739), .A2(new_n624), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n572), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n572), .B1(new_n739), .B2(new_n624), .ZN(new_n759));
  INV_X1    g558(.A(new_n755), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(G1337gat));
  OAI21_X1  g561(.A(G99gat), .B1(new_n740), .B2(new_n634), .ZN(new_n763));
  INV_X1    g562(.A(new_n750), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n659), .A2(new_n576), .A3(new_n617), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(G1338gat));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n445), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT114), .B(G106gat), .Z(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n618), .A2(new_n270), .A3(G106gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n750), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n770), .ZN(new_n775));
  INV_X1    g574(.A(new_n768), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n739), .B2(new_n445), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT53), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(G1339gat));
  OAI21_X1  g578(.A(KEYINPUT54), .B1(new_n606), .B2(new_n596), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n608), .A2(new_n605), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n613), .B1(new_n607), .B2(KEYINPUT54), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n680), .A2(new_n784), .A3(new_n614), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n524), .A2(new_n525), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n532), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n540), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n617), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n594), .B1(new_n786), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n594), .A2(new_n790), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n784), .A2(new_n614), .A3(new_n785), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n564), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n595), .A2(new_n681), .A3(new_n618), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n445), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n624), .A2(new_n484), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n798), .A2(new_n659), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(new_n543), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n484), .B1(new_n796), .B2(new_n797), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n631), .A2(new_n371), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n483), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n680), .A2(new_n271), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT116), .Z(new_n806));
  OAI22_X1  g605(.A1(new_n801), .A2(new_n271), .B1(new_n804), .B2(new_n806), .ZN(G1340gat));
  INV_X1    g606(.A(new_n804), .ZN(new_n808));
  AOI21_X1  g607(.A(G120gat), .B1(new_n808), .B2(new_n617), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n618), .A2(new_n276), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n800), .B2(new_n810), .ZN(G1341gat));
  NAND3_X1  g610(.A1(new_n800), .A2(G127gat), .A3(new_n679), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(KEYINPUT117), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(KEYINPUT117), .ZN(new_n814));
  AOI21_X1  g613(.A(G127gat), .B1(new_n808), .B2(new_n679), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(G1342gat));
  INV_X1    g615(.A(new_n594), .ZN(new_n817));
  OR3_X1    g616(.A1(new_n804), .A2(G134gat), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT118), .Z(new_n820));
  NAND2_X1  g619(.A1(new_n800), .A2(new_n594), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n818), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(G1343gat));
  OAI21_X1  g622(.A(new_n791), .B1(new_n542), .B2(new_n794), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n817), .ZN(new_n825));
  INV_X1    g624(.A(new_n795), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n827), .A2(new_n564), .B1(new_n681), .B2(new_n625), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n445), .A2(KEYINPUT57), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n270), .B1(new_n796), .B2(new_n797), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n828), .A2(new_n829), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n634), .A2(new_n799), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT119), .Z(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n205), .B1(new_n836), .B2(new_n542), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n542), .A2(G141gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n802), .A2(new_n445), .A3(new_n634), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT122), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(KEYINPUT122), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n483), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n833), .A2(new_n680), .A3(new_n835), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(new_n205), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n845), .B2(new_n205), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n840), .A2(new_n624), .A3(new_n839), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n844), .B1(new_n850), .B2(new_n838), .ZN(G1344gat));
  INV_X1    g650(.A(new_n843), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n203), .A3(new_n617), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n618), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(KEYINPUT59), .A3(new_n203), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n827), .A2(new_n564), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n625), .A2(new_n542), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n270), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n830), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n859), .A2(KEYINPUT57), .B1(new_n860), .B2(new_n831), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n617), .A3(new_n835), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n856), .B1(new_n862), .B2(G148gat), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n853), .B1(new_n855), .B2(new_n863), .ZN(G1345gat));
  OAI21_X1  g663(.A(G155gat), .B1(new_n836), .B2(new_n564), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n679), .A2(new_n207), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n843), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n867), .B(new_n868), .ZN(G1346gat));
  NOR3_X1   g668(.A1(new_n836), .A2(new_n208), .A3(new_n817), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n594), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n208), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n621), .A2(new_n483), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n803), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n796), .B2(new_n797), .ZN(new_n875));
  AOI21_X1  g674(.A(G169gat), .B1(new_n875), .B2(new_n680), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n659), .A2(new_n873), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT124), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(new_n798), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n878), .A2(KEYINPUT124), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n543), .A2(G169gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(G1348gat));
  INV_X1    g683(.A(G176gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n875), .A2(new_n885), .A3(new_n617), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n882), .A2(new_n617), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n885), .ZN(G1349gat));
  NAND3_X1  g687(.A1(new_n880), .A2(new_n679), .A3(new_n881), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G183gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n323), .A3(new_n679), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n324), .A3(new_n594), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n881), .A2(new_n594), .A3(new_n798), .A4(new_n879), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n895), .A2(new_n896), .A3(G190gat), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n895), .B2(G190gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n899), .B(new_n900), .ZN(G1351gat));
  NAND2_X1  g700(.A1(new_n634), .A2(new_n873), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n861), .B2(KEYINPUT126), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904));
  OAI221_X1 g703(.A(new_n904), .B1(new_n860), .B2(new_n831), .C1(new_n859), .C2(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G197gat), .B1(new_n906), .B2(new_n542), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n860), .A2(new_n902), .ZN(new_n908));
  INV_X1    g707(.A(G197gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n680), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(G1352gat));
  NAND3_X1  g710(.A1(new_n903), .A2(new_n617), .A3(new_n905), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n903), .A2(KEYINPUT127), .A3(new_n617), .A4(new_n905), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(G204gat), .A3(new_n915), .ZN(new_n916));
  NOR4_X1   g715(.A1(new_n860), .A2(G204gat), .A3(new_n618), .A4(new_n902), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT62), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1353gat));
  NOR2_X1   g718(.A1(new_n902), .A2(new_n564), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n225), .B1(new_n861), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT63), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n830), .A2(new_n920), .A3(new_n225), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1354gat));
  NOR3_X1   g723(.A1(new_n906), .A2(new_n226), .A3(new_n817), .ZN(new_n925));
  AOI21_X1  g724(.A(G218gat), .B1(new_n908), .B2(new_n594), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(G1355gat));
endmodule


