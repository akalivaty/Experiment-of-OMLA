//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n216), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n214), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XOR2_X1   g0035(.A(G107), .B(G116), .Z(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND3_X1  g0042(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G1), .A2(G13), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(new_n208), .B2(G20), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n248), .A2(new_n250), .B1(new_n249), .B2(new_n244), .ZN(new_n251));
  OAI21_X1  g0051(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n209), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n209), .A2(KEYINPUT68), .A3(G33), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n256), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n247), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n251), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G1), .A3(G13), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G77), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G222), .A2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G223), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n246), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n276), .A2(new_n281), .B1(new_n286), .B2(G226), .ZN(new_n287));
  OAI21_X1  g0087(.A(G274), .B1(new_n282), .B2(new_n246), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT67), .B1(new_n288), .B2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n285), .A2(new_n269), .A3(new_n290), .A4(G274), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n266), .A2(new_n267), .B1(G200), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n294), .B1(new_n267), .B2(new_n266), .C1(new_n295), .C2(new_n293), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n266), .C1(G179), .C2(new_n293), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT74), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G97), .ZN(new_n303));
  INV_X1    g0103(.A(G232), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G1698), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G226), .B2(G1698), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n306), .B2(new_n274), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(new_n283), .B1(new_n286), .B2(G238), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n292), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n292), .A3(new_n310), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n298), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n302), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n308), .A2(new_n292), .A3(new_n310), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n310), .B1(new_n308), .B2(new_n292), .ZN(new_n318));
  OAI21_X1  g0118(.A(G169), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n309), .A2(KEYINPUT72), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT13), .B1(new_n309), .B2(KEYINPUT72), .ZN(new_n322));
  OAI211_X1 g0122(.A(G179), .B(new_n313), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n314), .A2(new_n315), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n316), .A2(new_n320), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n259), .A2(G77), .A3(new_n260), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n247), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(KEYINPUT11), .A3(new_n247), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT73), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n243), .A2(G68), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT12), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n248), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(new_n336), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n325), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n341), .ZN(new_n343));
  OAI211_X1 g0143(.A(G190), .B(new_n313), .C1(new_n321), .C2(new_n322), .ZN(new_n344));
  OAI21_X1  g0144(.A(G200), .B1(new_n317), .B2(new_n318), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT70), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n277), .A2(G238), .A3(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G107), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n277), .A2(new_n279), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n350), .B1(new_n351), .B2(new_n277), .C1(new_n352), .C2(new_n304), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n283), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n289), .A2(new_n291), .B1(new_n286), .B2(G244), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n275), .B1(new_n208), .B2(G20), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n248), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT69), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n244), .A2(new_n275), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n262), .A2(new_n255), .B1(new_n209), .B2(new_n275), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n257), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n247), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n349), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n367), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(KEYINPUT70), .C1(new_n357), .C2(new_n356), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n354), .A2(new_n355), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n368), .B(new_n370), .C1(new_n295), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n298), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n367), .C1(G179), .C2(new_n371), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n301), .A2(new_n348), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT81), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n262), .B1(new_n208), .B2(G20), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(new_n248), .B1(new_n244), .B2(new_n262), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT77), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n270), .B2(KEYINPUT3), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT76), .B1(new_n272), .B2(G33), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(new_n270), .A3(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n272), .A2(KEYINPUT77), .A3(G33), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n381), .A2(new_n382), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(G20), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n387), .B1(new_n277), .B2(G20), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G68), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n203), .A3(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(G20), .B1(G159), .B2(new_n254), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT16), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n274), .B2(new_n209), .ZN(new_n400));
  INV_X1    g0200(.A(new_n388), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n277), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT16), .A3(new_n398), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n247), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n379), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n269), .A2(G232), .A3(new_n284), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT78), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT78), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n269), .A2(new_n284), .A3(new_n409), .A4(G232), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n292), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT79), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT79), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n292), .A3(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G226), .B2(new_n279), .ZN(new_n417));
  INV_X1    g0217(.A(G87), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n417), .A2(new_n274), .B1(new_n270), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(G179), .B1(new_n419), .B2(new_n283), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n408), .A2(new_n410), .B1(new_n289), .B2(new_n291), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n283), .ZN(new_n423));
  AOI21_X1  g0223(.A(G169), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n406), .A2(KEYINPUT18), .A3(new_n421), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT80), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n411), .A2(new_n292), .A3(new_n414), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n414), .B1(new_n411), .B2(new_n292), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n424), .B1(new_n431), .B2(new_n420), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n432), .A2(KEYINPUT80), .A3(KEYINPUT18), .A4(new_n406), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n421), .A2(new_n425), .ZN(new_n435));
  INV_X1    g0235(.A(new_n379), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n274), .A2(new_n388), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n202), .B1(new_n390), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n397), .A2(G20), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n254), .A2(G159), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n265), .B1(new_n442), .B2(KEYINPUT16), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT16), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n202), .B1(new_n389), .B2(new_n390), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n441), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n436), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n434), .B1(new_n435), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n433), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n377), .B1(new_n428), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n426), .A2(new_n427), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT81), .A3(new_n448), .A4(new_n433), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT83), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT82), .A2(G190), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT82), .A2(G190), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n419), .B2(new_n283), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n453), .B1(new_n431), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n413), .A2(new_n453), .A3(new_n415), .A4(new_n457), .ZN(new_n459));
  INV_X1    g0259(.A(new_n423), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n357), .B1(new_n460), .B2(new_n412), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n447), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT84), .A2(KEYINPUT17), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT84), .A2(KEYINPUT17), .ZN(new_n467));
  OAI221_X1 g0267(.A(new_n447), .B1(new_n467), .B2(new_n464), .C1(new_n458), .C2(new_n462), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(new_n452), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n376), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n208), .A2(G33), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n243), .A2(new_n473), .A3(new_n246), .A4(new_n245), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G116), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n244), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n245), .A2(new_n246), .B1(G20), .B2(new_n477), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n209), .C1(G33), .C2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT20), .B1(new_n479), .B2(new_n482), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n476), .B(new_n478), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT21), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n277), .A2(G264), .A3(G1698), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n277), .A2(G257), .A3(new_n279), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n274), .A2(G303), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n283), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n208), .A2(G45), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n283), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n494), .A2(new_n493), .ZN(new_n496));
  INV_X1    g0296(.A(new_n288), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n495), .A2(G270), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n486), .B(new_n298), .C1(new_n491), .C2(new_n498), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n491), .A2(new_n498), .A3(G179), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n485), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G200), .ZN(new_n503));
  INV_X1    g0303(.A(new_n485), .ZN(new_n504));
  INV_X1    g0304(.A(new_n456), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n503), .B(new_n504), .C1(new_n505), .C2(new_n502), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n485), .A3(G169), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT87), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n507), .A2(new_n508), .A3(new_n486), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n507), .B2(new_n486), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n501), .B(new_n506), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  INV_X1    g0312(.A(G244), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n352), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n277), .A2(G250), .A3(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n514), .A2(new_n480), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n283), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n495), .A2(G257), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n496), .A2(new_n497), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT85), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(G200), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n521), .B1(new_n517), .B2(new_n283), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT85), .B1(new_n526), .B2(new_n357), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n243), .A2(G97), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n474), .B2(new_n481), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n254), .A2(G77), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n351), .A2(KEYINPUT6), .A3(G97), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n481), .A2(new_n351), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n205), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n534), .B2(KEYINPUT6), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G20), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n400), .B1(new_n388), .B2(new_n386), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n531), .B(new_n536), .C1(new_n537), .C2(new_n351), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n530), .B1(new_n538), .B2(new_n247), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n526), .A2(G190), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n525), .A2(new_n527), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n247), .ZN(new_n542));
  INV_X1    g0342(.A(new_n530), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n523), .A2(new_n298), .ZN(new_n545));
  INV_X1    g0345(.A(G179), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n526), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g0349(.A(KEYINPUT90), .B(G294), .Z(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G33), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n277), .A2(G257), .A3(G1698), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n277), .A2(G250), .A3(new_n279), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n283), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n495), .A2(G264), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n546), .A3(new_n520), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n520), .A3(new_n556), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n298), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n277), .A2(new_n209), .A3(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n277), .A2(new_n564), .A3(new_n209), .A4(G87), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT89), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(KEYINPUT89), .A2(KEYINPUT23), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(G20), .A3(new_n351), .A4(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n567), .B(new_n568), .C1(new_n209), .C2(G107), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  OR3_X1    g0373(.A1(new_n573), .A2(KEYINPUT88), .A3(G20), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT88), .B1(new_n573), .B2(G20), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n571), .A2(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n561), .B1(new_n566), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n566), .A2(new_n561), .A3(new_n576), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n265), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n244), .A2(KEYINPUT25), .A3(new_n351), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT25), .B1(new_n244), .B2(new_n351), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n582), .A2(new_n583), .B1(new_n351), .B2(new_n474), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n558), .B(new_n560), .C1(new_n580), .C2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n492), .A2(G250), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n269), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n288), .B2(new_n492), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n277), .A2(G244), .A3(G1698), .ZN(new_n589));
  INV_X1    g0389(.A(G238), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n573), .C1(new_n352), .C2(new_n590), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n295), .B(new_n588), .C1(new_n283), .C2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n277), .A2(new_n209), .A3(G68), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n209), .B1(new_n303), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G87), .B2(new_n206), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n594), .B1(new_n257), .B2(new_n481), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(new_n247), .B1(new_n244), .B2(new_n364), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT86), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n475), .B2(G87), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n474), .A2(KEYINPUT86), .A3(new_n418), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n592), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n588), .B1(new_n283), .B2(new_n591), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n474), .A2(new_n364), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n605), .A2(new_n546), .B1(new_n599), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n298), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n604), .A2(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n579), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n247), .B1(new_n612), .B2(new_n577), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n557), .A2(G190), .A3(new_n520), .ZN(new_n614));
  INV_X1    g0414(.A(new_n584), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n559), .A2(G200), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n585), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  NOR4_X1   g0418(.A1(new_n472), .A2(new_n511), .A3(new_n549), .A4(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n374), .A2(KEYINPUT93), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n374), .A2(KEYINPUT93), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n347), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(new_n342), .B1(new_n468), .B2(new_n466), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n448), .A2(new_n426), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n297), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n300), .ZN(new_n627));
  INV_X1    g0427(.A(new_n588), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n591), .A2(KEYINPUT91), .A3(new_n283), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT91), .B1(new_n591), .B2(new_n283), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n298), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(G200), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n609), .A2(new_n632), .B1(new_n633), .B2(new_n604), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n541), .A3(new_n548), .A4(new_n617), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT92), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n560), .B1(G179), .B2(new_n559), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n613), .B2(new_n615), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n636), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n507), .A2(new_n486), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT87), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n507), .A2(new_n508), .A3(new_n486), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(new_n585), .A3(KEYINPUT92), .A4(new_n501), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n635), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n632), .A2(new_n609), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n634), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n648), .A2(new_n611), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n647), .B(new_n650), .C1(new_n651), .C2(new_n649), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n627), .B1(new_n472), .B2(new_n653), .ZN(G369));
  INV_X1    g0454(.A(new_n511), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT94), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n660));
  INV_X1    g0460(.A(G213), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT95), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT95), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n659), .A2(new_n665), .A3(new_n662), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n664), .A2(G343), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n485), .ZN(new_n668));
  MUX2_X1   g0468(.A(new_n637), .B(new_n655), .S(new_n668), .Z(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n667), .B1(new_n580), .B2(new_n584), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n639), .B1(new_n617), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n585), .A2(new_n667), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n617), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n585), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n667), .B1(new_n644), .B2(new_n501), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n212), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n215), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n526), .A2(new_n500), .A3(new_n557), .A4(new_n605), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n605), .A2(new_n555), .A3(new_n556), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n526), .A3(new_n500), .A4(KEYINPUT30), .ZN(new_n693));
  AOI21_X1  g0493(.A(G179), .B1(new_n491), .B2(new_n498), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n631), .A2(new_n523), .A3(new_n559), .A4(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n696), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT31), .B1(new_n696), .B2(new_n667), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n585), .A2(new_n611), .A3(new_n617), .ZN(new_n700));
  INV_X1    g0500(.A(new_n549), .ZN(new_n701));
  INV_X1    g0501(.A(new_n667), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n655), .A4(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n688), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n635), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n637), .A2(new_n639), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT96), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT96), .B1(new_n635), .B2(new_n706), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n634), .A2(new_n648), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT26), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n651), .A2(new_n649), .B1(new_n609), .B2(new_n632), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n709), .A2(new_n710), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .A3(new_n702), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n653), .B2(new_n667), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n704), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n687), .B1(new_n718), .B2(G1), .ZN(G364));
  AND2_X1   g0519(.A1(new_n209), .A2(G13), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n208), .B1(new_n720), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n682), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n670), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(G330), .B2(new_n669), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n723), .B(KEYINPUT97), .Z(new_n726));
  NOR2_X1   g0526(.A1(new_n681), .A2(new_n274), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G355), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G116), .B2(new_n212), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n681), .A2(new_n277), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G45), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n216), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n241), .A2(new_n732), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n729), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n246), .B1(G20), .B2(new_n298), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n726), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n209), .A2(G179), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n418), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n209), .A2(new_n546), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(G68), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n209), .A2(new_n546), .A3(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n295), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n743), .A2(new_n295), .A3(G200), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n749), .B1(new_n275), .B2(new_n751), .C1(new_n351), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n456), .A2(new_n750), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n274), .B(new_n753), .C1(G58), .C2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n747), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(KEYINPUT98), .A3(new_n456), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT98), .B1(new_n757), .B2(new_n456), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G50), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT99), .B1(G179), .B2(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(KEYINPUT99), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n209), .B1(new_n768), .B2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n767), .A2(new_n209), .A3(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G159), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT32), .Z(new_n774));
  NAND4_X1  g0574(.A1(new_n756), .A2(new_n763), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n550), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n769), .A2(new_n776), .B1(new_n777), .B2(new_n751), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n762), .B2(G326), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT100), .Z(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n274), .B1(new_n752), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n772), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(new_n744), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n755), .A2(G322), .B1(G303), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(KEYINPUT33), .A2(G317), .ZN(new_n786));
  AND2_X1   g0586(.A1(KEYINPUT33), .A2(G317), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n748), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n783), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n775), .B1(new_n780), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n742), .B1(new_n790), .B2(new_n739), .ZN(new_n791));
  INV_X1    g0591(.A(new_n738), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n669), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n725), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  NAND2_X1  g0595(.A1(new_n667), .A2(new_n367), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n372), .A2(new_n374), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n621), .A2(new_n367), .A3(new_n620), .A4(new_n667), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n653), .B2(new_n667), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n799), .B(new_n702), .C1(new_n646), .C2(new_n652), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n704), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n723), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  INV_X1    g0606(.A(new_n726), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n739), .A2(new_n736), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n275), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n739), .ZN(new_n810));
  INV_X1    g0610(.A(new_n751), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G159), .A2(new_n811), .B1(new_n748), .B2(G150), .ZN(new_n812));
  INV_X1    g0612(.A(G143), .ZN(new_n813));
  INV_X1    g0613(.A(G137), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n812), .B1(new_n813), .B2(new_n754), .C1(new_n761), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT34), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n752), .A2(new_n202), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n274), .B(new_n819), .C1(G50), .C2(new_n784), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  INV_X1    g0621(.A(new_n772), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n201), .B2(new_n769), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n817), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G303), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n771), .B1(new_n825), .B2(new_n761), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n274), .B1(new_n351), .B2(new_n744), .C1(new_n822), .C2(new_n777), .ZN(new_n827));
  INV_X1    g0627(.A(G294), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n754), .A2(new_n828), .B1(new_n477), .B2(new_n751), .ZN(new_n829));
  INV_X1    g0629(.A(new_n748), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n830), .A2(new_n781), .B1(new_n418), .B2(new_n752), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n826), .A2(new_n827), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n809), .B1(new_n810), .B2(new_n833), .C1(new_n799), .C2(new_n737), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n806), .A2(new_n834), .ZN(G384));
  NOR3_X1   g0635(.A1(new_n246), .A2(new_n209), .A3(new_n477), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n535), .B(KEYINPUT101), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT35), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT36), .ZN(new_n842));
  INV_X1    g0642(.A(new_n215), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n843), .A2(G77), .A3(new_n395), .A4(new_n396), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n249), .A2(G68), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n208), .B(G13), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n379), .B1(new_n849), .B2(new_n405), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n664), .A2(new_n666), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n451), .A2(new_n448), .A3(new_n433), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n854), .A2(new_n377), .B1(new_n468), .B2(new_n466), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(new_n855), .B2(new_n452), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n406), .B1(new_n432), .B2(new_n852), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n463), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n850), .B1(new_n432), .B2(new_n852), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n857), .B1(new_n463), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n848), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n853), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n470), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT38), .B1(new_n859), .B2(new_n861), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT104), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT104), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n869), .B(new_n866), .C1(new_n470), .C2(new_n864), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n863), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  NOR4_X1   g0672(.A1(new_n618), .A2(new_n549), .A3(new_n511), .A4(new_n667), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n696), .A2(new_n667), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT31), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n696), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n872), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n343), .A2(new_n702), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n346), .B2(new_n325), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n882));
  INV_X1    g0682(.A(new_n880), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n342), .A2(new_n347), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT102), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(new_n880), .C1(new_n346), .C2(new_n325), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n699), .A2(KEYINPUT105), .A3(new_n703), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n879), .A2(new_n887), .A3(new_n799), .A4(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT40), .B1(new_n871), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n865), .A2(new_n867), .ZN(new_n892));
  INV_X1    g0692(.A(new_n859), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n463), .A2(new_n858), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n406), .A2(new_n852), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n469), .B2(new_n624), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n848), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n889), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n891), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT105), .B1(new_n699), .B2(new_n703), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n699), .A2(KEYINPUT105), .A3(new_n703), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n472), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n688), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n904), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n625), .A2(new_n851), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n374), .A2(new_n667), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n802), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n887), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT103), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n912), .A2(KEYINPUT103), .A3(new_n887), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n871), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n856), .A2(new_n866), .ZN(new_n918));
  INV_X1    g0718(.A(new_n899), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n919), .B2(new_n896), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n918), .A2(new_n920), .A3(KEYINPUT39), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n871), .B2(KEYINPUT39), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n342), .A2(new_n667), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n910), .B(new_n917), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n472), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n715), .A3(new_n717), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n627), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n925), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n909), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n208), .B2(new_n720), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n909), .A2(new_n929), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n847), .B1(new_n931), .B2(new_n932), .ZN(G367));
  INV_X1    g0733(.A(KEYINPUT108), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n682), .B(KEYINPUT41), .Z(new_n935));
  INV_X1    g0735(.A(KEYINPUT45), .ZN(new_n936));
  INV_X1    g0736(.A(new_n673), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n637), .A2(new_n702), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n672), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n544), .A2(new_n667), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n541), .A2(new_n548), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n648), .A2(new_n667), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n936), .B1(new_n939), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n939), .A2(KEYINPUT44), .A3(new_n944), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT44), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n679), .B2(new_n943), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n670), .A2(new_n674), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n938), .B1(new_n672), .B2(new_n673), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n937), .A2(new_n677), .A3(new_n678), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n670), .B(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n675), .A2(new_n947), .A3(new_n951), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n718), .A2(new_n954), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n935), .B1(new_n960), .B2(new_n718), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(new_n722), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n941), .A2(new_n585), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n667), .B1(new_n963), .B2(new_n548), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n672), .A2(new_n673), .A3(new_n938), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n943), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n966), .B2(KEYINPUT42), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT42), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n674), .A2(new_n968), .A3(new_n678), .A4(new_n943), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT106), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n667), .A2(new_n603), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n634), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n647), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n965), .A2(KEYINPUT106), .A3(new_n968), .A4(new_n943), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n967), .A2(new_n971), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT42), .B1(new_n956), .B2(new_n944), .ZN(new_n978));
  INV_X1    g0778(.A(new_n964), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n971), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n974), .B(KEYINPUT43), .Z(new_n981));
  AOI22_X1  g0781(.A1(new_n977), .A2(KEYINPUT107), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n976), .A2(new_n979), .A3(new_n978), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT107), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n983), .A2(new_n984), .A3(new_n975), .A4(new_n971), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n675), .A2(new_n944), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n982), .A2(new_n987), .A3(new_n985), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n934), .B1(new_n962), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n977), .A2(KEYINPUT107), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n980), .A2(new_n981), .ZN(new_n994));
  AND4_X1   g0794(.A1(new_n987), .A2(new_n993), .A3(new_n985), .A4(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n987), .B1(new_n982), .B2(new_n985), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(KEYINPUT108), .C1(new_n722), .C2(new_n961), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n740), .B1(new_n212), .B2(new_n364), .C1(new_n731), .C2(new_n233), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n726), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n274), .B1(new_n830), .B2(new_n776), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n772), .A2(G317), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n744), .A2(new_n477), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(KEYINPUT46), .B2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1002), .B(new_n1005), .C1(KEYINPUT46), .C2(new_n1004), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n752), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n811), .A2(G283), .B1(new_n1007), .B2(G97), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n825), .B2(new_n754), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G107), .B2(new_n770), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1006), .B(new_n1010), .C1(new_n777), .C2(new_n761), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n277), .B1(new_n275), .B2(new_n752), .C1(new_n822), .C2(new_n814), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n751), .A2(new_n249), .B1(new_n744), .B2(new_n201), .ZN(new_n1013));
  INV_X1    g0813(.A(G159), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n830), .A2(new_n1014), .B1(new_n253), .B2(new_n754), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n770), .A2(G68), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n813), .C2(new_n761), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT47), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1001), .B1(new_n1020), .B2(new_n739), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n974), .A2(new_n792), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n999), .A2(new_n1023), .ZN(G387));
  XOR2_X1   g0824(.A(new_n682), .B(KEYINPUT110), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n718), .B2(new_n958), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n718), .B2(new_n958), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n958), .A2(new_n722), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n684), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n727), .A2(new_n1030), .B1(new_n351), .B2(new_n681), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n230), .A2(new_n732), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n263), .A2(new_n249), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n684), .B(new_n732), .C1(new_n202), .C2(new_n275), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n730), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1031), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n807), .B1(new_n1037), .B2(new_n740), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n274), .B1(new_n752), .B2(new_n477), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n755), .A2(G317), .B1(G303), .B2(new_n811), .ZN(new_n1040));
  INV_X1    g0840(.A(G322), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1040), .B1(new_n777), .B2(new_n830), .C1(new_n761), .C2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n770), .A2(G283), .B1(new_n550), .B2(new_n784), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1039), .B(new_n1049), .C1(G326), .C2(new_n772), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n274), .B1(new_n1007), .B2(G97), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n275), .B2(new_n744), .C1(new_n822), .C2(new_n253), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT109), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n769), .A2(new_n364), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n755), .A2(G50), .B1(G68), .B2(new_n811), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n262), .B2(new_n830), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(G159), .C2(new_n762), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1050), .A2(new_n1051), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1038), .B1(new_n674), .B2(new_n792), .C1(new_n1059), .C2(new_n810), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1029), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1028), .A2(new_n1061), .ZN(G393));
  NAND2_X1  g0862(.A1(new_n954), .A2(new_n959), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n721), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n761), .A2(new_n253), .B1(new_n1014), .B2(new_n754), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT51), .Z(new_n1066));
  NOR2_X1   g0866(.A1(new_n769), .A2(new_n275), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n263), .A2(new_n811), .B1(new_n748), .B2(G50), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n202), .B2(new_n744), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n277), .B1(new_n418), .B2(new_n752), .C1(new_n822), .C2(new_n813), .ZN(new_n1070));
  OR4_X1    g0870(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n811), .A2(G294), .B1(new_n784), .B2(G283), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n825), .B2(new_n830), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n274), .B1(new_n351), .B2(new_n752), .C1(new_n822), .C2(new_n1041), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(G116), .C2(new_n770), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n762), .A2(G317), .B1(G311), .B2(new_n755), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT52), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1080), .A2(KEYINPUT111), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(KEYINPUT111), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1071), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n739), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n740), .B1(new_n481), .B2(new_n212), .C1(new_n731), .C2(new_n237), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n726), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n738), .B2(new_n944), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1064), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n718), .A2(new_n958), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1063), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n960), .A3(new_n1025), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1088), .A2(new_n1091), .A3(KEYINPUT112), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT112), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(G390));
  NAND2_X1  g0895(.A1(new_n913), .A2(new_n924), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT39), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n892), .A2(new_n900), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n869), .B1(new_n856), .B2(new_n866), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n865), .A2(KEYINPUT104), .A3(new_n867), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n862), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n865), .A2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1099), .A2(new_n1100), .B1(new_n1102), .B2(new_n848), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1096), .B(new_n1098), .C1(new_n1103), .C2(new_n1097), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n901), .A2(new_n924), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n887), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n714), .A2(new_n702), .A3(new_n799), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n911), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n884), .A2(new_n886), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n800), .B1(new_n1110), .B2(new_n882), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(KEYINPUT113), .A3(new_n704), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT113), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n887), .A2(new_n799), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n804), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1104), .A2(new_n1109), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n906), .A2(new_n905), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(G330), .A3(new_n1111), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT114), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1107), .A2(new_n911), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1115), .B2(new_n1112), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n879), .A2(G330), .A3(new_n888), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1106), .B1(new_n1125), .B2(new_n800), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1106), .B1(new_n804), .B2(new_n800), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1125), .B2(new_n1114), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1124), .A2(new_n1126), .B1(new_n912), .B2(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1125), .A2(new_n472), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n927), .A2(new_n1130), .A3(new_n627), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1122), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1128), .A2(new_n912), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1131), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n1122), .C1(new_n1117), .C2(new_n1120), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1133), .A2(new_n1139), .A3(new_n1025), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1104), .A2(new_n1109), .A3(new_n1116), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n922), .B2(new_n1096), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1141), .B1(new_n1143), .B2(new_n1119), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1098), .B1(new_n1103), .B2(new_n1097), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n737), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n808), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n744), .A2(new_n253), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT53), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1149), .B1(new_n1014), .B2(new_n769), .C1(new_n761), .C2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n748), .A2(G137), .B1(new_n1007), .B2(G50), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n821), .B2(new_n754), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  INV_X1    g0954(.A(G125), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n277), .B1(new_n751), .B2(new_n1154), .C1(new_n822), .C2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1151), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT115), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(KEYINPUT115), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1067), .B1(new_n762), .B2(G283), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n819), .B1(G97), .B2(new_n811), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n755), .A2(G116), .B1(G107), .B2(new_n748), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n277), .B(new_n745), .C1(new_n772), .C2(G294), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1158), .A2(new_n1159), .A3(new_n1164), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n726), .B1(new_n263), .B2(new_n1147), .C1(new_n1165), .C2(new_n810), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n1144), .A2(new_n721), .B1(new_n1146), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1140), .A2(new_n1168), .ZN(G378));
  OAI21_X1  g0969(.A(new_n1017), .B1(new_n761), .B2(new_n477), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT116), .Z(new_n1171));
  AOI22_X1  g0971(.A1(new_n748), .A2(G97), .B1(new_n1007), .B2(G58), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n351), .B2(new_n754), .C1(new_n364), .C2(new_n751), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n277), .A2(G41), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n275), .B2(new_n744), .C1(new_n822), .C2(new_n781), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1171), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1174), .ZN(new_n1177));
  INV_X1    g0977(.A(G41), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G50), .B1(new_n270), .B2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1176), .A2(KEYINPUT58), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n755), .A2(G128), .B1(G137), .B2(new_n811), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1154), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n748), .A2(G132), .B1(new_n784), .B2(new_n1182), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n253), .B2(new_n769), .C1(new_n1155), .C2(new_n761), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n270), .B(new_n1178), .C1(new_n752), .C2(new_n1014), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n772), .B2(G124), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1180), .B1(KEYINPUT58), .B2(new_n1176), .C1(new_n1186), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n739), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n722), .B(new_n682), .C1(new_n249), .C2(new_n808), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n852), .A2(new_n266), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT55), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n301), .B(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1197));
  XOR2_X1   g0997(.A(new_n1196), .B(new_n1197), .Z(new_n1198));
  OAI211_X1 g0998(.A(new_n1192), .B(new_n1193), .C1(new_n1198), .C2(new_n737), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT118), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1118), .A2(new_n1111), .A3(KEYINPUT40), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n918), .A2(new_n920), .ZN(new_n1203));
  OAI21_X1  g1003(.A(G330), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1196), .B(new_n1197), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n891), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n902), .B1(new_n1103), .B2(new_n889), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n688), .B1(new_n903), .B2(new_n901), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1198), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1201), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n925), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n925), .B(new_n1201), .C1(new_n1206), .C2(new_n1209), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1200), .B1(new_n1214), .B2(new_n722), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1141), .B(new_n1136), .C1(new_n1143), .C2(new_n1119), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1137), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT57), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1216), .A2(new_n1137), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1145), .A2(new_n923), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n917), .A2(new_n910), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n1206), .C2(new_n1209), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1207), .A2(new_n1208), .A3(new_n1198), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1205), .B1(new_n891), .B2(new_n1204), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n925), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(KEYINPUT57), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1025), .B1(new_n1219), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1215), .B1(new_n1218), .B2(new_n1227), .ZN(G375));
  INV_X1    g1028(.A(new_n935), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1134), .A2(new_n1135), .A3(new_n1131), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1138), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1106), .A2(new_n736), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1055), .B1(G283), .B2(new_n755), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT119), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n811), .A2(G107), .B1(new_n784), .B2(G97), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n477), .B2(new_n830), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n274), .B1(new_n275), .B2(new_n752), .C1(new_n822), .C2(new_n825), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(G294), .C2(new_n762), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n748), .A2(new_n1182), .B1(new_n784), .B2(G159), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n814), .B2(new_n754), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n277), .B1(new_n201), .B2(new_n752), .C1(new_n822), .C2(new_n1150), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(G132), .C2(new_n762), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n769), .A2(new_n249), .B1(new_n253), .B2(new_n751), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT120), .Z(new_n1244));
  AOI22_X1  g1044(.A1(new_n1234), .A2(new_n1238), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n726), .B1(G68), .B2(new_n1147), .C1(new_n1245), .C2(new_n810), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT121), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1136), .A2(new_n722), .B1(new_n1232), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1231), .A2(new_n1248), .ZN(G381));
  NAND3_X1  g1049(.A1(new_n1028), .A2(new_n794), .A3(new_n1061), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(G384), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1251), .ZN(new_n1252));
  OR3_X1    g1052(.A1(new_n1252), .A2(G378), .A3(G375), .ZN(G407));
  AOI21_X1  g1053(.A(new_n1026), .B1(new_n1121), .B2(new_n1132), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1167), .B1(new_n1254), .B2(new_n1139), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n661), .A2(G343), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G375), .C2(new_n1257), .ZN(G409));
  NAND2_X1  g1058(.A1(G393), .A2(G396), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1250), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1260), .A2(KEYINPUT123), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(KEYINPUT123), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n999), .A2(new_n1023), .A3(new_n1094), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n992), .A2(new_n998), .B1(new_n1022), .B2(new_n1021), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(new_n1094), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1263), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G387), .A2(G390), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n1265), .A3(new_n1271), .A4(new_n1264), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT126), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1215), .C1(new_n1218), .C2(new_n1227), .ZN(new_n1275));
  AOI221_X4 g1075(.A(new_n935), .B1(new_n1216), .B2(new_n1137), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1222), .A2(new_n722), .A3(new_n1225), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1199), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1255), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1256), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1230), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1284), .A2(new_n1138), .A3(new_n1025), .A4(new_n1285), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1286), .A2(G384), .A3(new_n1248), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G384), .B1(new_n1286), .B2(new_n1248), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT122), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G2897), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1281), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  OAI221_X1 g1092(.A(KEYINPUT122), .B1(new_n1290), .B2(new_n1281), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT122), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1292), .A2(new_n1293), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1280), .A2(new_n1281), .A3(new_n1295), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1274), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1287), .A2(new_n1288), .A3(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1280), .A2(new_n1281), .A3(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1256), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1309), .B2(new_n1295), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1303), .B1(new_n1311), .B2(new_n1297), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1298), .A2(new_n1304), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1273), .B1(new_n1309), .B2(new_n1305), .ZN(new_n1314));
  AND4_X1   g1114(.A1(new_n1303), .A2(new_n1297), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1302), .B1(new_n1312), .B2(new_n1315), .ZN(G405));
  XNOR2_X1  g1116(.A(G375), .B(G378), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1295), .A2(KEYINPUT127), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1317), .B(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(new_n1274), .ZN(G402));
endmodule


