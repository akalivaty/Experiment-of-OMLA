//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OR3_X1    g0007(.A1(new_n207), .A2(KEYINPUT65), .A3(G13), .ZN(new_n208));
  OAI21_X1  g0008(.A(KEYINPUT65), .B1(new_n207), .B2(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n206), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n214), .A2(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT66), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(new_n202), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(new_n216), .B2(new_n202), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT67), .Z(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n214), .A2(KEYINPUT0), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n215), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT68), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  INV_X1    g0029(.A(G87), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n206), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n232));
  INV_X1    g0032(.A(G77), .ZN(new_n233));
  INV_X1    g0033(.A(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G107), .ZN(new_n235));
  OAI221_X1 g0035(.A(new_n232), .B1(new_n233), .B2(new_n234), .C1(new_n235), .C2(new_n213), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n207), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n226), .A2(new_n238), .ZN(G361));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  INV_X1    g0045(.A(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT2), .B(G226), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n244), .B(new_n249), .Z(G358));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT71), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(G68), .B(G77), .Z(new_n255));
  XOR2_X1   g0055(.A(G50), .B(G58), .Z(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT73), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT73), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n261), .A2(new_n267), .A3(G226), .A4(new_n268), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n261), .A2(new_n267), .A3(G232), .A4(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G97), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n272), .A2(KEYINPUT79), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  OAI211_X1 g0074(.A(G1), .B(G13), .C1(new_n263), .C2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n272), .B2(KEYINPUT79), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n275), .A2(new_n279), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(new_n229), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT13), .B1(new_n277), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n273), .B2(new_n276), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G200), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT80), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n286), .A2(KEYINPUT80), .A3(new_n287), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n292), .A2(new_n285), .A3(G190), .A4(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n295), .A2(G50), .B1(G20), .B2(new_n228), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT74), .B1(new_n263), .B2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT74), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(new_n221), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n296), .B1(new_n300), .B2(new_n233), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n220), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n309), .A2(new_n221), .A3(G1), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n311), .A2(KEYINPUT12), .A3(G68), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT12), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n310), .B2(new_n228), .ZN(new_n314));
  INV_X1    g0114(.A(new_n303), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n278), .A2(G20), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n312), .A2(new_n314), .B1(new_n228), .B2(new_n317), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n307), .A2(new_n308), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n290), .A2(new_n294), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n288), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n286), .A2(new_n287), .ZN(new_n323));
  OAI211_X1 g0123(.A(KEYINPUT14), .B(G169), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT14), .B1(new_n289), .B2(G169), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n292), .A2(new_n285), .A3(new_n293), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n319), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n321), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT84), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT72), .B(G226), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n282), .B1(new_n283), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n261), .A2(new_n267), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(G222), .A3(new_n268), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n261), .A2(new_n267), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G77), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(G1698), .ZN(new_n339));
  INV_X1    g0139(.A(G223), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n336), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n334), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G190), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n295), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT8), .B(G58), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n300), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n303), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n310), .A2(new_n303), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n316), .A2(G50), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G50), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n349), .A2(new_n351), .B1(new_n352), .B2(new_n310), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT9), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n348), .A2(KEYINPUT9), .A3(new_n353), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n344), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G200), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n343), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT10), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n356), .A2(new_n357), .ZN(new_n362));
  INV_X1    g0162(.A(new_n360), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT10), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n344), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n343), .A2(new_n327), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n354), .B1(new_n343), .B2(G169), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n343), .A2(G169), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n372), .A2(KEYINPUT75), .A3(new_n354), .A4(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n335), .A2(G232), .A3(new_n268), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n337), .A2(G107), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n375), .B(new_n376), .C1(new_n339), .C2(new_n229), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n342), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n282), .B1(new_n283), .B2(new_n234), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(new_n383), .A3(new_n380), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(G200), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n383), .B1(new_n378), .B2(new_n380), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT76), .B(new_n379), .C1(new_n377), .C2(new_n342), .ZN(new_n387));
  OAI21_X1  g0187(.A(G190), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n295), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n346), .A2(new_n389), .B1(new_n221), .B2(new_n233), .ZN(new_n390));
  XOR2_X1   g0190(.A(KEYINPUT15), .B(G87), .Z(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(new_n299), .A3(new_n297), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n392), .B2(KEYINPUT77), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(KEYINPUT77), .B2(new_n392), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n303), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n310), .A2(new_n233), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n317), .B2(new_n233), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT78), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(new_n401), .A3(new_n398), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n385), .A2(new_n388), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n382), .A2(new_n404), .A3(new_n384), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n327), .B1(new_n386), .B2(new_n387), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n399), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n366), .A2(new_n374), .A3(new_n403), .A4(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT83), .ZN(new_n409));
  INV_X1    g0209(.A(new_n349), .ZN(new_n410));
  INV_X1    g0210(.A(new_n346), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n316), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n410), .A2(new_n412), .B1(new_n311), .B2(new_n411), .ZN(new_n413));
  INV_X1    g0213(.A(G58), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n228), .ZN(new_n415));
  OAI21_X1  g0215(.A(G20), .B1(new_n415), .B2(new_n202), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n295), .A2(G159), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n259), .A2(new_n260), .A3(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT7), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n264), .A2(new_n221), .A3(new_n266), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT81), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n422), .B1(new_n421), .B2(new_n423), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n420), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n418), .B1(new_n426), .B2(G68), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n315), .B1(new_n427), .B2(KEYINPUT16), .ZN(new_n428));
  INV_X1    g0228(.A(new_n418), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n421), .A2(new_n423), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n337), .A2(new_n221), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(new_n423), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n429), .B1(new_n432), .B2(new_n228), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT16), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n413), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n340), .A2(new_n268), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n437), .B1(G226), .B2(new_n268), .C1(new_n259), .C2(new_n260), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G87), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n275), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n283), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n281), .B1(new_n442), .B2(G232), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(G179), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n282), .B1(new_n283), .B2(new_n246), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT82), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(KEYINPUT82), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n409), .B(KEYINPUT18), .C1(new_n436), .C2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT81), .B1(new_n419), .B2(KEYINPUT7), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n430), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(KEYINPUT16), .B(new_n429), .C1(new_n455), .C2(new_n228), .ZN(new_n456));
  AOI21_X1  g0256(.A(G20), .B1(new_n261), .B2(new_n267), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n420), .B1(new_n457), .B2(KEYINPUT7), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n418), .B1(new_n458), .B2(G68), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n456), .B(new_n303), .C1(KEYINPUT16), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n413), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n440), .A2(new_n445), .ZN(new_n462));
  INV_X1    g0262(.A(G190), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(G200), .B2(new_n462), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT17), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n456), .A2(new_n303), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n459), .A2(KEYINPUT16), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n461), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n444), .A2(KEYINPUT82), .A3(new_n446), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT82), .B1(new_n444), .B2(new_n446), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT18), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n409), .A2(KEYINPUT18), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n472), .A2(new_n475), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n452), .A2(new_n468), .A3(new_n469), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n408), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n331), .A2(new_n332), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n332), .B1(new_n331), .B2(new_n481), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT85), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT4), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n234), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n335), .A2(new_n486), .A3(new_n268), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n335), .A2(G250), .A3(G1698), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n261), .A2(new_n267), .A3(new_n268), .A4(new_n488), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT85), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n264), .A2(new_n266), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G244), .A3(new_n268), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(new_n487), .B1(G33), .B2(G283), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n489), .A2(new_n490), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n342), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT5), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT86), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(G41), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n274), .A2(KEYINPUT86), .A3(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G45), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G1), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G274), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n502), .A2(new_n505), .A3(new_n342), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n504), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n275), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n212), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n497), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n404), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n496), .B2(new_n342), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n327), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n310), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n278), .A2(G33), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n349), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G97), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n521), .A2(new_n516), .A3(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n524), .A2(new_n221), .B1(new_n233), .B2(new_n389), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n458), .B2(G107), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n517), .B(new_n520), .C1(new_n526), .C2(new_n315), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n513), .A2(new_n515), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n514), .A2(G190), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n520), .A2(new_n517), .ZN(new_n530));
  INV_X1    g0330(.A(new_n526), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n303), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n529), .B(new_n532), .C1(new_n359), .C2(new_n514), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n300), .B2(new_n516), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n493), .A2(new_n221), .A3(G68), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n221), .B1(new_n271), .B2(new_n534), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n230), .A2(new_n516), .A3(new_n235), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n391), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n540), .A2(new_n303), .B1(new_n310), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n519), .A2(G87), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n229), .A2(G1698), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n493), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G116), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n342), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n275), .A2(new_n508), .A3(G250), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n505), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(G190), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n548), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n493), .B2(new_n545), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n275), .B1(new_n556), .B2(new_n547), .ZN(new_n557));
  OAI21_X1  g0357(.A(G200), .B1(new_n557), .B2(new_n552), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n519), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n542), .B1(new_n541), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n550), .A2(G179), .A3(new_n553), .ZN(new_n562));
  OAI21_X1  g0362(.A(G169), .B1(new_n557), .B2(new_n552), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n544), .A2(new_n559), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n528), .A2(new_n533), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n528), .A2(new_n533), .A3(KEYINPUT87), .A4(new_n565), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT88), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n213), .A2(G1698), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n493), .B(new_n571), .C1(G257), .C2(G1698), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G303), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n261), .B2(new_n267), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n570), .B(new_n342), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n509), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n506), .B1(new_n577), .B2(G270), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n337), .A2(G303), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n275), .B1(new_n580), .B2(new_n572), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n581), .A2(new_n570), .ZN(new_n582));
  OAI21_X1  g0382(.A(G200), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n311), .A2(G116), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n519), .B2(G116), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G283), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n586), .B(new_n221), .C1(G33), .C2(new_n516), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n587), .B(new_n303), .C1(new_n221), .C2(G116), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n579), .ZN(new_n593));
  INV_X1    g0393(.A(new_n582), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n583), .B(new_n592), .C1(new_n595), .C2(new_n463), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n579), .A2(new_n582), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n591), .A2(G169), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n404), .B1(new_n585), .B2(new_n590), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(KEYINPUT21), .C1(new_n582), .C2(new_n579), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(G179), .A3(new_n591), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n596), .A2(new_n600), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n493), .A2(new_n221), .A3(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT22), .ZN(new_n606));
  OR3_X1    g0406(.A1(new_n230), .A2(KEYINPUT22), .A3(G20), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n337), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT24), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT89), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n221), .B2(G107), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n611), .A2(KEYINPUT23), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(KEYINPUT23), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(new_n221), .B2(new_n555), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n608), .B2(new_n614), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n303), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n310), .A2(KEYINPUT25), .A3(new_n235), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT25), .B1(new_n310), .B2(new_n235), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n560), .A2(new_n235), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n212), .A2(G1698), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G250), .B2(G1698), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n259), .A2(new_n260), .ZN(new_n626));
  INV_X1    g0426(.A(G294), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n625), .A2(new_n626), .B1(new_n263), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n342), .ZN(new_n629));
  OAI211_X1 g0429(.A(G264), .B(new_n275), .C1(new_n502), .C2(new_n508), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n507), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n404), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n507), .A2(new_n629), .A3(new_n327), .A4(new_n630), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n623), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n631), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G190), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n631), .A2(G200), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n617), .A2(new_n638), .A3(new_n622), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n604), .A2(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n485), .A2(new_n568), .A3(new_n569), .A4(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n447), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n436), .A2(KEYINPUT18), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n476), .B1(new_n472), .B2(new_n447), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n407), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n329), .A2(new_n330), .B1(new_n320), .B2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n469), .A2(new_n468), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n652), .A2(new_n366), .B1(new_n371), .B2(new_n373), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n513), .A2(new_n515), .A3(new_n527), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT92), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT26), .A4(new_n565), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n565), .A2(new_n513), .A3(new_n515), .A4(new_n527), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT92), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n404), .B1(new_n550), .B2(new_n553), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n557), .A2(new_n327), .A3(new_n552), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT90), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n562), .A2(new_n563), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n561), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n544), .A2(new_n559), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n658), .B1(new_n668), .B2(new_n528), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n656), .A2(new_n659), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n636), .A2(KEYINPUT91), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n623), .A2(new_n673), .A3(new_n635), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n665), .A2(new_n561), .B1(new_n544), .B2(new_n559), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n528), .A2(new_n533), .A3(new_n676), .A4(new_n640), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n666), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n653), .B1(new_n484), .B2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n278), .A2(new_n221), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n592), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n671), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n604), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n687), .B1(new_n617), .B2(new_n622), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n641), .A2(new_n692), .B1(new_n636), .B2(new_n687), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n686), .ZN(new_n696));
  INV_X1    g0496(.A(new_n641), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n673), .B1(new_n623), .B2(new_n635), .ZN(new_n698));
  AOI211_X1 g0498(.A(KEYINPUT91), .B(new_n634), .C1(new_n617), .C2(new_n622), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n686), .B(KEYINPUT93), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n696), .A2(new_n697), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n694), .A2(new_n703), .ZN(G399));
  NOR2_X1   g0504(.A1(new_n211), .A2(G41), .ZN(new_n705));
  NOR4_X1   g0505(.A1(new_n705), .A2(new_n278), .A3(G116), .A4(new_n538), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n218), .B2(new_n705), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n550), .A2(new_n553), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n595), .A2(new_n327), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n512), .A2(new_n712), .A3(new_n631), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT94), .B1(new_n514), .B2(new_n637), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n595), .A2(new_n327), .ZN(new_n716));
  AND4_X1   g0516(.A1(new_n550), .A2(new_n553), .A3(new_n629), .A4(new_n630), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n514), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT30), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NOR4_X1   g0521(.A1(new_n718), .A2(new_n595), .A3(new_n721), .A4(new_n327), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n715), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n709), .B1(new_n723), .B2(new_n687), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n642), .A2(new_n568), .A3(new_n569), .A4(new_n702), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n701), .A2(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n716), .A2(new_n719), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n713), .A2(new_n714), .ZN(new_n730));
  INV_X1    g0530(.A(new_n711), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n722), .B1(new_n733), .B2(KEYINPUT95), .ZN(new_n734));
  OR3_X1    g0534(.A1(new_n715), .A2(new_n720), .A3(KEYINPUT95), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n726), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  INV_X1    g0538(.A(new_n666), .ZN(new_n739));
  AND4_X1   g0539(.A1(new_n528), .A2(new_n533), .A3(new_n676), .A4(new_n640), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n695), .B1(new_n699), .B2(new_n698), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n656), .A2(new_n659), .A3(new_n669), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n701), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n677), .B1(new_n636), .B2(new_n695), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT26), .B1(new_n668), .B2(new_n528), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n747), .B(new_n666), .C1(KEYINPUT26), .C2(new_n657), .ZN(new_n748));
  OAI211_X1 g0548(.A(KEYINPUT29), .B(new_n687), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n738), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n708), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n309), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n278), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n705), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n691), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G330), .B2(new_n690), .ZN(new_n758));
  OAI21_X1  g0558(.A(G20), .B1(KEYINPUT97), .B2(G169), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(KEYINPUT97), .A2(G169), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n220), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n221), .A2(new_n463), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n327), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n221), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G322), .A2(new_n767), .B1(new_n771), .B2(G329), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n359), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n764), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G326), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n327), .A2(new_n359), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n764), .A2(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n772), .B1(new_n574), .B2(new_n774), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n768), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(KEYINPUT33), .A2(G317), .ZN(new_n781));
  AND2_X1   g0581(.A1(KEYINPUT33), .A2(G317), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(new_n768), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n768), .A2(new_n765), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n783), .B1(new_n784), .B2(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n221), .B1(new_n769), .B2(G190), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n337), .B1(new_n627), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n778), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT98), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n785), .A2(new_n235), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n777), .A2(new_n352), .B1(new_n766), .B2(new_n414), .ZN(new_n794));
  INV_X1    g0594(.A(new_n787), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n793), .B(new_n794), .C1(G77), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n789), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G97), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n228), .A2(new_n779), .B1(new_n774), .B2(new_n230), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n337), .ZN(new_n800));
  INV_X1    g0600(.A(G159), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n770), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT32), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n796), .A2(new_n798), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n791), .B1(new_n792), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n804), .A2(new_n792), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n763), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n762), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n257), .A2(G45), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT96), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n219), .A2(new_n503), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n211), .A2(new_n493), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n211), .A2(new_n337), .ZN(new_n818));
  INV_X1    g0618(.A(G116), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(G355), .B1(new_n819), .B2(new_n211), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n812), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n756), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n807), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n810), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n690), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n758), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  AND4_X1   g0627(.A1(new_n399), .A2(new_n405), .A3(new_n406), .A4(new_n687), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n399), .A2(new_n686), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n403), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n407), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n744), .B(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n756), .B1(new_n738), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n738), .B2(new_n832), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G143), .A2(new_n767), .B1(new_n795), .B2(G159), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n777), .C1(new_n837), .C2(new_n779), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT100), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n797), .A2(G58), .ZN(new_n841));
  INV_X1    g0641(.A(new_n774), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n626), .B1(new_n842), .B2(G50), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n785), .A2(new_n228), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G132), .B2(new_n771), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n840), .A2(new_n841), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n839), .A2(KEYINPUT34), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n785), .A2(new_n230), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G116), .B2(new_n795), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n627), .B2(new_n766), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n235), .A2(new_n774), .B1(new_n779), .B2(new_n784), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n777), .A2(new_n574), .B1(new_n770), .B2(new_n786), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n337), .A3(new_n798), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n846), .A2(new_n847), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n762), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n763), .A2(new_n809), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT99), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n822), .B1(new_n859), .B2(new_n233), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n856), .B(new_n860), .C1(new_n831), .C2(new_n809), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n834), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  INV_X1    g0663(.A(new_n524), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT35), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(KEYINPUT35), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(G116), .A3(new_n222), .A4(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n218), .B(G77), .C1(new_n414), .C2(new_n228), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n201), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n278), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n684), .B1(new_n460), .B2(new_n461), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n647), .B2(new_n650), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n436), .A2(KEYINPUT102), .A3(new_n465), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n466), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n684), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n472), .B1(new_n447), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n875), .B1(new_n436), .B2(new_n465), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT37), .B1(new_n472), .B2(new_n475), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n883), .A2(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n874), .B1(new_n877), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n429), .B1(new_n455), .B2(new_n228), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n434), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n413), .B1(new_n428), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n684), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n480), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n466), .B1(new_n891), .B2(new_n684), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n891), .A2(new_n644), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT37), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n885), .A2(new_n876), .A3(new_n466), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n893), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n887), .A2(new_n888), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n893), .A2(new_n898), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n874), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n888), .B1(new_n902), .B2(new_n899), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT103), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(G169), .B1(new_n322), .B2(new_n323), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT14), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n292), .A2(new_n285), .A3(new_n293), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n907), .A2(new_n324), .B1(new_n908), .B2(G179), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n909), .A2(new_n319), .A3(new_n686), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n898), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n893), .B2(new_n898), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT39), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT103), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n887), .A2(new_n888), .A3(new_n899), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n904), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n647), .A2(new_n881), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n831), .B(new_n702), .C1(new_n670), .C2(new_n678), .ZN(new_n919));
  INV_X1    g0719(.A(new_n828), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n319), .A2(new_n687), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n320), .B(new_n922), .C1(new_n909), .C2(new_n319), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n329), .A2(new_n921), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n919), .A2(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n902), .A2(new_n899), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n918), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n917), .A2(KEYINPUT104), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT104), .B1(new_n917), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n745), .B(new_n749), .C1(new_n482), .C2(new_n483), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n653), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n831), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n923), .B2(new_n924), .ZN(new_n935));
  OAI211_X1 g0735(.A(KEYINPUT31), .B(new_n686), .C1(new_n733), .C2(new_n722), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n724), .A2(new_n725), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n887), .A2(new_n899), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n935), .A2(KEYINPUT106), .A3(new_n937), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n940), .A2(KEYINPUT40), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n935), .A2(new_n926), .A3(new_n937), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT105), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n485), .A2(new_n937), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(G330), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n933), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n278), .B2(new_n753), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n933), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n873), .B1(new_n956), .B2(new_n957), .ZN(G367));
  OAI211_X1 g0758(.A(new_n528), .B(new_n533), .C1(new_n532), .C2(new_n702), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n654), .A2(new_n701), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n696), .A2(new_n697), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n528), .B1(new_n959), .B2(new_n636), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n702), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n666), .A2(new_n544), .A3(new_n687), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n676), .B1(new_n544), .B2(new_n687), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT43), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n967), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n964), .A2(new_n972), .A3(new_n971), .A4(new_n966), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n694), .A2(new_n961), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n705), .B(KEYINPUT41), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n962), .B1(new_n693), .B2(new_n696), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(new_n691), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n738), .A2(new_n750), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n700), .A2(new_n702), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n962), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n986), .B2(new_n961), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n959), .A2(new_n960), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(KEYINPUT44), .A3(new_n961), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT44), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n703), .B2(new_n988), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n990), .A2(new_n994), .A3(new_n694), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n694), .B1(new_n990), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g0796(.A(KEYINPUT107), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(KEYINPUT107), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n983), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n980), .B1(new_n999), .B2(new_n751), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n979), .B1(new_n1000), .B2(new_n755), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n244), .A2(new_n816), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n811), .B1(new_n210), .B2(new_n541), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n756), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G58), .A2(new_n842), .B1(new_n771), .B2(G137), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT108), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT108), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n837), .A2(new_n766), .B1(new_n779), .B2(new_n801), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n777), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1008), .B1(G143), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n785), .A2(new_n233), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n201), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n795), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n335), .C1(new_n228), .C2(new_n789), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n842), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT46), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n774), .B2(new_n819), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1016), .B(new_n1018), .C1(new_n235), .C2(new_n789), .ZN(new_n1019));
  INV_X1    g0819(.A(G317), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n785), .A2(new_n516), .B1(new_n770), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n626), .B1(new_n777), .B2(new_n786), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G294), .A2(new_n780), .B1(new_n767), .B2(G303), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n784), .C2(new_n787), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1011), .A2(new_n1015), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1004), .B1(new_n1027), .B2(new_n762), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n970), .B2(new_n824), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT109), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1001), .A2(new_n1030), .ZN(G387));
  OR2_X1    g0831(.A1(new_n693), .A2(new_n824), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n816), .B1(new_n249), .B2(new_n503), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n538), .A2(G116), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n818), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n346), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT50), .B1(new_n346), .B2(G50), .ZN(new_n1038));
  AOI21_X1  g0838(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1037), .A2(new_n1034), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1036), .A2(new_n1040), .B1(new_n235), .B2(new_n211), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n756), .B1(new_n1041), .B2(new_n812), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n777), .A2(new_n801), .B1(new_n774), .B2(new_n233), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n785), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n626), .B(new_n1043), .C1(G97), .C2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G68), .A2(new_n795), .B1(new_n771), .B2(G150), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G50), .A2(new_n767), .B1(new_n780), .B2(new_n411), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n797), .A2(new_n391), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n842), .A2(G294), .B1(new_n797), .B2(G283), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G317), .A2(new_n767), .B1(new_n795), .B2(G303), .ZN(new_n1051));
  INV_X1    g0851(.A(G322), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1051), .B1(new_n786), .B2(new_n779), .C1(new_n1052), .C2(new_n777), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT49), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n626), .B1(new_n770), .B2(new_n775), .C1(new_n819), .C2(new_n785), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT110), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1056), .A2(KEYINPUT49), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1049), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1042), .B1(new_n1062), .B2(new_n762), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n982), .A2(new_n755), .B1(new_n1032), .B2(new_n1063), .ZN(new_n1064));
  OR3_X1    g0864(.A1(new_n983), .A2(G41), .A3(new_n211), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n751), .A2(new_n982), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  NOR2_X1   g0867(.A1(new_n995), .A2(new_n996), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n999), .B(new_n705), .C1(new_n983), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n961), .A2(new_n810), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n254), .A2(new_n211), .A3(new_n493), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n811), .B1(new_n516), .B2(new_n210), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n756), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n777), .A2(new_n837), .B1(new_n766), .B2(new_n801), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT112), .Z(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n780), .A2(new_n1013), .B1(new_n795), .B2(new_n411), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G68), .A2(new_n842), .B1(new_n771), .B2(G143), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n789), .A2(new_n233), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n848), .A2(new_n1080), .A3(new_n626), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n777), .A2(new_n1020), .B1(new_n766), .B2(new_n786), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT52), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n793), .B1(G283), .B2(new_n842), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1052), .B2(new_n770), .ZN(new_n1087));
  OR3_X1    g0887(.A1(new_n1085), .A2(new_n335), .A3(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n779), .A2(new_n574), .B1(new_n787), .B2(new_n627), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G116), .B2(new_n797), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT113), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n1082), .A2(new_n1083), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1073), .B1(new_n1092), .B2(new_n762), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1068), .A2(new_n755), .B1(new_n1070), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1069), .A2(new_n1094), .ZN(G390));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n925), .B2(new_n910), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n910), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n828), .B1(new_n744), .B2(new_n831), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n909), .A2(new_n922), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n331), .B2(new_n922), .ZN(new_n1101));
  OAI211_X1 g0901(.A(KEYINPUT114), .B(new_n1098), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1097), .B(new_n1102), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n830), .A2(new_n407), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n687), .B(new_n1106), .C1(new_n746), .C2(new_n748), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1107), .A2(new_n920), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(new_n1101), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n941), .A2(new_n1098), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n737), .A2(G330), .A3(new_n935), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1105), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n904), .A2(new_n916), .B1(new_n1115), .B2(new_n1096), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1111), .B1(new_n1116), .B2(new_n1102), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n935), .A2(G330), .A3(new_n937), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1114), .B(new_n755), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n808), .B1(new_n1104), .B2(new_n1103), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n756), .B1(new_n858), .B2(new_n411), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n779), .A2(new_n235), .B1(new_n787), .B2(new_n516), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G283), .B2(new_n1009), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n844), .B1(G87), .B2(new_n842), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G116), .A2(new_n767), .B1(new_n771), .B2(G294), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n335), .A2(new_n1080), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n774), .A2(new_n837), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT54), .B(G143), .Z(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT115), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n795), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1044), .A2(new_n1013), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G132), .A2(new_n767), .B1(new_n780), .B2(G137), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1009), .A2(G128), .B1(new_n771), .B2(G125), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(new_n335), .C1(new_n801), .C2(new_n789), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1127), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1121), .B1(new_n1139), .B2(new_n762), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1120), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT117), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1119), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT118), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1114), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1145));
  OAI211_X1 g0945(.A(G330), .B(new_n937), .C1(new_n482), .C2(new_n483), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n931), .A2(new_n1146), .A3(new_n653), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n831), .C1(new_n726), .C2(new_n736), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1101), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1118), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1099), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n937), .A2(G330), .A3(new_n831), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1101), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1113), .A2(new_n1108), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1147), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1145), .A2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1114), .B(new_n1156), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n705), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT118), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1119), .A2(new_n1142), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1144), .A2(new_n1160), .A3(new_n1162), .ZN(G378));
  OAI211_X1 g0963(.A(new_n943), .B(G330), .C1(new_n948), .C2(new_n949), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n366), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n369), .A2(new_n370), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n354), .A2(new_n881), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  OR3_X1    g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n928), .A2(new_n929), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT104), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1104), .A2(new_n1103), .A3(new_n1098), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n927), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n917), .A2(KEYINPUT104), .A3(new_n927), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1175), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1164), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1176), .B1(new_n928), .B2(new_n929), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1181), .A2(new_n1182), .A3(new_n1175), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1164), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1184), .A2(new_n755), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n756), .B1(new_n858), .B2(new_n1013), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G50), .B1(new_n266), .B2(new_n274), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n785), .A2(new_n414), .B1(new_n770), .B2(new_n784), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n274), .B(new_n626), .C1(new_n774), .C2(new_n233), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G68), .C2(new_n797), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1009), .A2(G116), .B1(new_n795), .B2(new_n391), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G97), .A2(new_n780), .B1(new_n767), .B2(G107), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1191), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1132), .A2(new_n842), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n797), .A2(G150), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G125), .A2(new_n1009), .B1(new_n767), .B2(G128), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G132), .A2(new_n780), .B1(new_n795), .B2(G137), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT59), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(KEYINPUT119), .A2(G124), .ZN(new_n1206));
  AND2_X1   g1006(.A1(KEYINPUT119), .A2(G124), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n771), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1044), .A2(G159), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1208), .A2(new_n1209), .A3(new_n263), .A4(new_n274), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1199), .B1(new_n1198), .B2(new_n1197), .C1(new_n1205), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1190), .B1(new_n1211), .B2(new_n762), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1175), .B2(new_n809), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1189), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1147), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1159), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1184), .A2(new_n1188), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT57), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1184), .A2(new_n1217), .A3(KEYINPUT57), .A4(new_n1188), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n705), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1215), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT120), .Z(G375));
  NAND2_X1  g1024(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1101), .A2(new_n808), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n756), .B1(new_n858), .B2(G68), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1009), .A2(G132), .B1(new_n771), .B2(G128), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n836), .B2(new_n766), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n780), .B2(new_n1132), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n774), .A2(new_n801), .B1(new_n787), .B2(new_n837), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n626), .B(new_n1231), .C1(G58), .C2(new_n1044), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(new_n352), .C2(new_n789), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n774), .A2(new_n516), .B1(new_n770), .B2(new_n574), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT121), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n766), .A2(new_n784), .B1(new_n787), .B2(new_n235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G294), .B2(new_n1009), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1012), .B1(G116), .B2(new_n780), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1237), .A2(new_n337), .A3(new_n1048), .A4(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1233), .B1(new_n1235), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1227), .B1(new_n1240), .B2(new_n762), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT122), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1225), .A2(new_n755), .B1(new_n1226), .B2(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1156), .A2(new_n980), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1225), .A2(new_n1216), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT123), .Z(G381));
  XNOR2_X1  g1047(.A(new_n1223), .B(KEYINPUT120), .ZN(new_n1248));
  INV_X1    g1048(.A(G378), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  INV_X1    g1052(.A(G390), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n862), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(G381), .A2(G387), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(G407));
  NAND2_X1  g1056(.A1(new_n685), .A2(G213), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT124), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1251), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(G407), .A2(new_n1259), .A3(G213), .ZN(G409));
  XNOR2_X1  g1060(.A(G393), .B(G396), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1001), .A2(G390), .A3(new_n1030), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G390), .B1(new_n1001), .B2(new_n1030), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1264), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(G393), .B(new_n826), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1262), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1223), .A2(G378), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1218), .A2(new_n980), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1272), .A2(new_n1214), .A3(G378), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1152), .A2(new_n1147), .A3(KEYINPUT60), .A4(new_n1155), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1275), .A2(new_n705), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1156), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1278), .B2(new_n1245), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(G384), .A3(new_n1243), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1279), .B2(new_n1243), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1271), .A2(new_n1274), .A3(new_n1257), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n705), .A3(new_n1221), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1249), .B1(new_n1286), .B2(new_n1215), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1287), .A2(new_n1258), .A3(new_n1273), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1282), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1280), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(new_n1270), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1270), .A2(new_n1284), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1257), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(G2897), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1283), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT126), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1258), .A2(G2897), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1296), .B(new_n1297), .C1(new_n1283), .C2(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1289), .A2(new_n1280), .A3(new_n1295), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1298), .B1(new_n1289), .B2(new_n1280), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT126), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1293), .B1(new_n1303), .B2(new_n1288), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1269), .B1(new_n1292), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT125), .ZN(new_n1306));
  NOR4_X1   g1106(.A1(new_n1287), .A2(new_n1273), .A3(new_n1294), .A4(new_n1290), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(KEYINPUT63), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1284), .A2(KEYINPUT125), .A3(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1271), .A2(new_n1257), .A3(new_n1274), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(new_n1302), .A3(new_n1299), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1265), .A2(new_n1268), .A3(new_n1293), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1290), .A2(new_n1309), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1288), .B2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1308), .A2(new_n1310), .A3(new_n1312), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1305), .A2(new_n1316), .ZN(G405));
  NOR3_X1   g1117(.A1(new_n1263), .A2(new_n1261), .A3(new_n1264), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1267), .B1(new_n1266), .B2(new_n1262), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1290), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1265), .A2(new_n1283), .A3(new_n1268), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1321), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1325), .A2(new_n1250), .A3(new_n1271), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1250), .B2(new_n1271), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


