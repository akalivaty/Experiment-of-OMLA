//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  INV_X1    g008(.A(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(new_n210), .A3(new_n211), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n206), .B1(new_n208), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT67), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(KEYINPUT23), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n205), .B1(new_n217), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n211), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n212), .A2(KEYINPUT69), .A3(new_n230), .A4(new_n207), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n231), .A2(new_n206), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n230), .A3(new_n207), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n233), .A2(new_n234), .B1(new_n225), .B2(new_n222), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(KEYINPUT68), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT23), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n232), .A2(new_n235), .A3(KEYINPUT25), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n229), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT26), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n239), .A2(new_n243), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n220), .A2(KEYINPUT26), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n244), .A2(new_n245), .B1(G183gat), .B2(G190gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT27), .B(G183gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n211), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT28), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n248), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n242), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT73), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n257));
  XNOR2_X1  g056(.A(G127gat), .B(G134gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n259), .A2(KEYINPUT1), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n258), .B(new_n260), .C1(new_n256), .C2(KEYINPUT1), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n262), .A2(KEYINPUT72), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT72), .B1(new_n262), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n229), .A2(new_n241), .B1(new_n246), .B2(new_n251), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n255), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(KEYINPUT73), .A3(new_n266), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n270), .A2(G227gat), .A3(G233gat), .A4(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT33), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n204), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(KEYINPUT32), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n272), .B(KEYINPUT32), .C1(new_n273), .C2(new_n204), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n271), .ZN(new_n279));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT34), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n278), .A2(KEYINPUT74), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n283), .B1(new_n278), .B2(KEYINPUT74), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT36), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n278), .A2(new_n283), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n281), .B(KEYINPUT34), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n277), .A3(new_n276), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT76), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n287), .A2(new_n289), .A3(new_n293), .A4(new_n290), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n286), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G197gat), .B(G204gat), .Z(new_n299));
  AOI21_X1  g098(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G211gat), .B(G218gat), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n299), .B2(new_n300), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT77), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n307), .B(new_n302), .C1(new_n299), .C2(new_n300), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n268), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n242), .A2(new_n313), .A3(new_n252), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n310), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n268), .A2(new_n313), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n317), .B(new_n309), .C1(new_n268), .C2(new_n311), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(KEYINPUT78), .B(new_n310), .C1(new_n312), .C2(new_n314), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n298), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n321), .A2(KEYINPUT30), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n298), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n321), .A2(KEYINPUT79), .A3(KEYINPUT30), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT79), .B1(new_n321), .B2(KEYINPUT30), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327));
  INV_X1    g126(.A(G85gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT0), .B(G57gat), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n329), .B(new_n330), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT82), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT80), .B(G141gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G141gat), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT81), .B1(new_n337), .B2(G148gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT81), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(new_n335), .A3(G141gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n333), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n338), .A2(new_n340), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n343), .B(KEYINPUT82), .C1(new_n335), .C2(new_n334), .ZN(new_n344));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  INV_X1    g144(.A(G155gat), .ZN(new_n346));
  INV_X1    g145(.A(G162gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n345), .B1(new_n348), .B2(KEYINPUT2), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n342), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n262), .A2(new_n263), .ZN(new_n351));
  XNOR2_X1  g150(.A(G141gat), .B(G148gat), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n348), .B(new_n345), .C1(new_n352), .C2(KEYINPUT2), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n350), .B(new_n353), .C1(new_n264), .C2(new_n265), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT5), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n350), .A2(new_n353), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g163(.A(new_n351), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT83), .B(KEYINPUT3), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n353), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n357), .A2(new_n362), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n369), .B(new_n371), .C1(new_n372), .C2(new_n355), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n363), .A2(new_n365), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n354), .ZN(new_n375));
  INV_X1    g174(.A(new_n362), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n361), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n332), .B1(new_n370), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n369), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n376), .B1(new_n380), .B2(new_n359), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n332), .B1(new_n381), .B2(KEYINPUT39), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT87), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n384), .B(new_n332), .C1(new_n381), .C2(KEYINPUT39), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT39), .B1(new_n375), .B2(new_n376), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n383), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT40), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n379), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n383), .A2(KEYINPUT40), .A3(new_n385), .A4(new_n390), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n326), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G228gat), .ZN(new_n396));
  INV_X1    g195(.A(G233gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n309), .B1(new_n368), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n304), .B1(KEYINPUT84), .B2(new_n305), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n305), .A2(KEYINPUT84), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n404), .A2(new_n367), .B1(new_n353), .B2(new_n350), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n401), .A2(new_n399), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n306), .A2(new_n400), .A3(new_n308), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n363), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT85), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n368), .A2(new_n400), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n310), .ZN(new_n414));
  AND4_X1   g213(.A1(KEYINPUT85), .A2(new_n414), .A3(new_n411), .A4(new_n398), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n406), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT31), .B(G50gat), .Z(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(G22gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT86), .ZN(new_n421));
  INV_X1    g220(.A(new_n417), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n422), .B(new_n406), .C1(new_n412), .C2(new_n415), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n418), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n418), .B2(new_n423), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n379), .A2(KEYINPUT6), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT90), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n379), .A2(new_n429), .A3(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n319), .A2(new_n320), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT37), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n298), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT38), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n379), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n370), .A2(new_n378), .A3(new_n332), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n321), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n431), .A2(new_n437), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n315), .A2(new_n318), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT38), .B1(new_n444), .B2(KEYINPUT37), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n434), .A2(new_n298), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT89), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n395), .B(new_n426), .C1(new_n443), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n427), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n321), .A2(KEYINPUT30), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n321), .A2(KEYINPUT79), .A3(KEYINPUT30), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n449), .A2(new_n454), .A3(new_n322), .A4(new_n323), .ZN(new_n455));
  INV_X1    g254(.A(new_n421), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n414), .A2(new_n411), .A3(new_n398), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT85), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n422), .B1(new_n459), .B2(new_n406), .ZN(new_n460));
  INV_X1    g259(.A(new_n423), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n418), .A2(new_n421), .A3(new_n423), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n295), .A2(new_n448), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n426), .B1(new_n284), .B2(new_n285), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT35), .B1(new_n467), .B2(new_n455), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n370), .A2(new_n378), .A3(new_n332), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(new_n379), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n428), .A2(new_n430), .B1(new_n470), .B2(new_n439), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n464), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT35), .ZN(new_n473));
  INV_X1    g272(.A(new_n326), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n287), .A2(new_n289), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n466), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(G15gat), .A2(G22gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(G15gat), .A2(G22gat), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT93), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G15gat), .ZN(new_n482));
  INV_X1    g281(.A(G22gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n485));
  NAND2_X1  g284(.A1(G15gat), .A2(G22gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G1gat), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n481), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n481), .A2(new_n487), .B1(KEYINPUT16), .B2(new_n488), .ZN(new_n490));
  OAI21_X1  g289(.A(G8gat), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n481), .A2(new_n487), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(KEYINPUT16), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n481), .A2(new_n487), .A3(new_n488), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G57gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G64gat), .ZN(new_n500));
  INV_X1    g299(.A(G64gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G57gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G71gat), .ZN(new_n504));
  INV_X1    g303(.A(G78gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G71gat), .A2(G78gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT9), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n503), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(new_n510), .B2(new_n503), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n498), .B1(KEYINPUT21), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G211gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G127gat), .B(G155gat), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n513), .A2(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(new_n520), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n518), .B(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT96), .B(G183gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n522), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527));
  INV_X1    g326(.A(G29gat), .ZN(new_n528));
  INV_X1    g327(.A(G36gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G29gat), .A2(G36gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G50gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G43gat), .ZN(new_n536));
  INV_X1    g335(.A(G43gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(G50gat), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n536), .A2(new_n538), .A3(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n530), .A2(KEYINPUT92), .A3(new_n531), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT92), .B1(new_n530), .B2(new_n531), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n533), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT15), .B1(new_n536), .B2(new_n538), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n538), .A3(KEYINPUT15), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n540), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G92gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n328), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n550), .A2(new_n553), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G99gat), .B(G106gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n328), .B2(new_n554), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n548), .A2(new_n566), .B1(KEYINPUT41), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n532), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n530), .A2(KEYINPUT92), .A3(new_n531), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n539), .A2(new_n544), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n533), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(KEYINPUT17), .A3(new_n540), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n559), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n563), .A2(new_n558), .A3(new_n564), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT17), .B1(new_n574), .B2(new_n540), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n568), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n567), .A2(KEYINPUT41), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n581), .B(new_n582), .Z(new_n583));
  XOR2_X1   g382(.A(G190gat), .B(G218gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT97), .ZN(new_n585));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n583), .B(new_n587), .Z(new_n588));
  NOR2_X1   g387(.A1(new_n526), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n507), .B(new_n506), .C1(new_n590), .C2(new_n509), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n503), .A2(new_n508), .A3(new_n510), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n591), .B(new_n592), .C1(new_n560), .C2(new_n565), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n577), .B(new_n576), .C1(new_n511), .C2(new_n512), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT100), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n596), .B(KEYINPUT101), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT10), .B1(new_n593), .B2(new_n594), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n604), .B2(new_n566), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n603), .A2(new_n578), .A3(KEYINPUT98), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n598), .B1(new_n600), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n606), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT98), .B1(new_n603), .B2(new_n578), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT99), .B1(new_n618), .B2(new_n596), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620));
  INV_X1    g419(.A(new_n596), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n607), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n598), .B(new_n613), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n612), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n498), .B(new_n548), .ZN(new_n626));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n489), .A2(new_n490), .A3(G8gat), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT17), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n548), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n634), .A3(new_n575), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT94), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n498), .A2(new_n548), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .A4(new_n627), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT95), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT18), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT94), .B1(new_n639), .B2(KEYINPUT18), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n491), .A2(new_n497), .B1(new_n574), .B2(new_n540), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n580), .A2(new_n498), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n575), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n644), .B2(new_n627), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n629), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT91), .ZN(new_n647));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648));
  INV_X1    g447(.A(G197gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT11), .B(G169gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n646), .B2(new_n647), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n478), .A2(new_n589), .A3(new_n625), .A4(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n449), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(new_n488), .ZN(G1324gat));
  NOR2_X1   g462(.A1(new_n661), .A2(new_n474), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(G8gat), .B1(new_n661), .B2(new_n474), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(KEYINPUT42), .A3(new_n665), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(G1325gat));
  INV_X1    g470(.A(new_n661), .ZN(new_n672));
  AOI21_X1  g471(.A(G15gat), .B1(new_n672), .B2(new_n475), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n661), .A2(new_n295), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(G15gat), .B2(new_n674), .ZN(G1326gat));
  NOR2_X1   g474(.A1(new_n661), .A2(new_n426), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT43), .B(G22gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  INV_X1    g477(.A(new_n588), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n466), .B2(new_n477), .ZN(new_n680));
  INV_X1    g479(.A(new_n526), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n654), .A2(new_n655), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n681), .A2(new_n624), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n449), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n528), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n680), .A2(new_n689), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT44), .B(new_n679), .C1(new_n466), .C2(new_n477), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n683), .B(KEYINPUT103), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n449), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n688), .A2(new_n695), .ZN(G1328gat));
  OAI21_X1  g495(.A(G36gat), .B1(new_n694), .B2(new_n474), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n684), .A2(G36gat), .A3(new_n474), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(G1329gat));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n537), .A3(new_n475), .ZN(new_n701));
  INV_X1    g500(.A(new_n295), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n693), .B(new_n702), .C1(new_n690), .C2(new_n691), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n701), .B1(new_n704), .B2(new_n537), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT47), .B1(new_n701), .B2(KEYINPUT104), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1330gat));
  INV_X1    g506(.A(KEYINPUT48), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n693), .B(new_n464), .C1(new_n690), .C2(new_n691), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G50gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n685), .A2(new_n535), .A3(new_n464), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT105), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(KEYINPUT105), .B2(new_n710), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(new_n708), .ZN(G1331gat));
  AOI211_X1 g514(.A(new_n625), .B(new_n656), .C1(new_n466), .C2(new_n477), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n716), .A2(new_n589), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n449), .B(KEYINPUT106), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n717), .A2(new_n326), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n717), .A2(new_n724), .A3(new_n326), .A4(new_n721), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1333gat));
  NAND4_X1  g527(.A1(new_n716), .A2(new_n702), .A3(G71gat), .A4(new_n589), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n717), .ZN(new_n732));
  INV_X1    g531(.A(new_n475), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n504), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n731), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n731), .B2(new_n734), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n464), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(G78gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  NAND2_X1  g540(.A1(new_n526), .A2(new_n682), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT111), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n624), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n692), .A2(new_n686), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n692), .A2(KEYINPUT112), .A3(new_n686), .A4(new_n744), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(G85gat), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n478), .B2(new_n588), .ZN(new_n751));
  AOI211_X1 g550(.A(KEYINPUT113), .B(new_n679), .C1(new_n466), .C2(new_n477), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n743), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT51), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n755), .B(new_n743), .C1(new_n751), .C2(new_n752), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n624), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n686), .A2(new_n328), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n749), .B1(new_n757), .B2(new_n758), .ZN(G1336gat));
  NAND3_X1  g558(.A1(new_n692), .A2(new_n326), .A3(new_n744), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n474), .A2(G92gat), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n754), .A2(new_n624), .A3(new_n756), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n692), .A2(new_n702), .A3(new_n744), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G99gat), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n757), .A2(G99gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n733), .ZN(G1338gat));
  NOR2_X1   g571(.A1(new_n426), .A2(G106gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n754), .A2(new_n624), .A3(new_n756), .A4(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n464), .B(new_n744), .C1(new_n690), .C2(new_n691), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT114), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n778), .A3(G106gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT53), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n774), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n607), .B2(new_n600), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n622), .B2(new_n619), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n607), .A2(new_n600), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n613), .B1(new_n790), .B2(new_n785), .ZN(new_n791));
  OAI211_X1 g590(.A(KEYINPUT116), .B(new_n786), .C1(new_n622), .C2(new_n619), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n789), .A2(KEYINPUT55), .A3(new_n791), .A4(new_n792), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n656), .A2(new_n623), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n629), .B(new_n653), .C1(new_n640), .C2(new_n645), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n644), .A2(new_n627), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n626), .A2(new_n628), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n652), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n624), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n797), .A2(new_n798), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n798), .B1(new_n797), .B2(new_n804), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n588), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n795), .A2(new_n623), .A3(new_n796), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n588), .A3(new_n803), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n526), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  NOR4_X1   g612(.A1(new_n526), .A2(new_n588), .A3(new_n624), .A4(new_n656), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n804), .B1(new_n808), .B2(new_n682), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n798), .A3(new_n804), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n679), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n681), .B1(new_n820), .B2(new_n810), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT118), .B1(new_n821), .B2(new_n814), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n326), .A2(new_n449), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n816), .A2(new_n822), .A3(new_n426), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n733), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n682), .ZN(new_n827));
  INV_X1    g626(.A(new_n467), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n816), .A2(new_n822), .A3(new_n828), .A4(new_n718), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n829), .A2(G113gat), .A3(new_n326), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n682), .B2(new_n830), .ZN(G1340gat));
  INV_X1    g630(.A(new_n829), .ZN(new_n832));
  INV_X1    g631(.A(G120gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n624), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT119), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n474), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n824), .A2(new_n733), .A3(new_n625), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n833), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT120), .ZN(G1341gat));
  INV_X1    g638(.A(G127gat), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n826), .A2(new_n840), .A3(new_n526), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n832), .A2(new_n474), .A3(new_n681), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n840), .B2(new_n842), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n825), .B2(new_n588), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n326), .A2(new_n679), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n844), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n847), .B1(new_n829), .B2(new_n849), .ZN(new_n850));
  OR3_X1    g649(.A1(new_n829), .A2(new_n847), .A3(new_n849), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n846), .A2(KEYINPUT122), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n850), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n845), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(G1343gat));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n816), .A2(new_n822), .A3(new_n857), .A4(new_n464), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n295), .A2(new_n823), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n793), .A2(KEYINPUT123), .A3(KEYINPUT55), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n656), .A2(new_n860), .A3(new_n623), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n795), .A2(new_n796), .B1(KEYINPUT123), .B2(new_n793), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n804), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n679), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n681), .B1(new_n864), .B2(new_n810), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n464), .B1(new_n865), .B2(new_n814), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n859), .B1(new_n866), .B2(KEYINPUT57), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n334), .B1(new_n868), .B2(new_n682), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n702), .A2(new_n426), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n816), .A2(new_n822), .A3(new_n718), .A4(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n326), .A2(new_n682), .A3(G141gat), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT58), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n813), .B1(new_n812), .B2(new_n815), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n821), .A2(KEYINPUT118), .A3(new_n814), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n879), .A2(KEYINPUT124), .A3(new_n718), .A4(new_n870), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n871), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n873), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n869), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n871), .A2(new_n881), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n881), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n884), .B(new_n872), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n876), .B1(new_n885), .B2(new_n890), .ZN(G1344gat));
  AOI21_X1  g690(.A(new_n326), .B1(new_n880), .B2(new_n882), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n335), .A3(new_n624), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n816), .A2(new_n822), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT57), .B1(new_n895), .B2(new_n426), .ZN(new_n896));
  INV_X1    g695(.A(new_n859), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n866), .A2(KEYINPUT57), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n896), .A2(new_n624), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n894), .B1(new_n868), .B2(new_n625), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n335), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n893), .B1(new_n900), .B2(new_n902), .ZN(G1345gat));
  NAND3_X1  g702(.A1(new_n892), .A2(new_n346), .A3(new_n681), .ZN(new_n904));
  OAI21_X1  g703(.A(G155gat), .B1(new_n868), .B2(new_n526), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  OAI211_X1 g705(.A(new_n347), .B(new_n848), .C1(new_n886), .C2(new_n887), .ZN(new_n907));
  OAI21_X1  g706(.A(G162gat), .B1(new_n868), .B2(new_n679), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n718), .A2(new_n474), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n475), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n879), .A2(new_n426), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n682), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n816), .A2(new_n822), .A3(new_n449), .A4(new_n828), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n474), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n218), .A3(new_n656), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(G1348gat));
  NOR3_X1   g720(.A1(new_n916), .A2(new_n219), .A3(new_n625), .ZN(new_n922));
  AOI21_X1  g721(.A(G176gat), .B1(new_n919), .B2(new_n624), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1349gat));
  OAI21_X1  g723(.A(G183gat), .B1(new_n916), .B2(new_n526), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n247), .A3(new_n681), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT60), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n919), .A2(new_n211), .A3(new_n588), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n933));
  INV_X1    g732(.A(new_n913), .ZN(new_n934));
  NOR4_X1   g733(.A1(new_n895), .A2(new_n464), .A3(new_n934), .A4(new_n914), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n588), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n936), .B2(G190gat), .ZN(new_n937));
  AOI211_X1 g736(.A(KEYINPUT61), .B(new_n211), .C1(new_n935), .C2(new_n588), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(G1351gat));
  NOR2_X1   g738(.A1(new_n895), .A2(new_n686), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(new_n326), .A3(new_n870), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n649), .A3(new_n656), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n896), .A2(new_n898), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n910), .A2(new_n295), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n943), .A2(new_n656), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n945), .B2(new_n649), .ZN(G1352gat));
  AND2_X1   g745(.A1(new_n940), .A2(new_n870), .ZN(new_n947));
  XNOR2_X1  g746(.A(KEYINPUT127), .B(G204gat), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n947), .A2(new_n326), .A3(new_n624), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n896), .A2(new_n624), .A3(new_n898), .A4(new_n944), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n948), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n941), .A2(new_n954), .A3(new_n624), .A4(new_n949), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n515), .A3(new_n681), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n896), .A2(new_n681), .A3(new_n898), .A4(new_n944), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  INV_X1    g760(.A(G218gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n941), .A2(new_n962), .A3(new_n588), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n943), .A2(new_n588), .A3(new_n944), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(new_n962), .ZN(G1355gat));
endmodule


