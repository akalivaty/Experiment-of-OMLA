//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT27), .B(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT28), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n208), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n213), .B1(new_n211), .B2(new_n212), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n209), .A2(new_n210), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n224));
  OR2_X1    g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT23), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT25), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(new_n226), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(new_n220), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n236), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n219), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT1), .B1(new_n240), .B2(KEYINPUT67), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(KEYINPUT67), .B2(new_n240), .ZN(new_n242));
  NOR2_X1   g041(.A1(G127gat), .A2(G134gat), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT66), .B(G127gat), .Z(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(G134gat), .ZN(new_n245));
  INV_X1    g044(.A(G113gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G120gat), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT68), .B(G120gat), .Z(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n246), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n250), .A2(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(KEYINPUT69), .ZN(new_n252));
  AND2_X1   g051(.A1(G127gat), .A2(G134gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n252), .C1(new_n243), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n242), .A2(new_n245), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n235), .B1(new_n222), .B2(new_n221), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n232), .B1(new_n258), .B2(new_n224), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n233), .A2(KEYINPUT25), .ZN(new_n260));
  OAI22_X1  g059(.A1(new_n259), .A2(KEYINPUT25), .B1(new_n236), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n250), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n245), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n255), .A2(new_n249), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(new_n267), .A3(new_n219), .ZN(new_n268));
  INV_X1    g067(.A(G227gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n257), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT33), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n205), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT34), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n268), .ZN(new_n276));
  INV_X1    g075(.A(new_n271), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI211_X1 g077(.A(KEYINPUT34), .B(new_n271), .C1(new_n257), .C2(new_n268), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n274), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n272), .A2(KEYINPUT32), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n284), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n286), .B2(new_n280), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G78gat), .B(G106gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT31), .B(G50gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G22gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT79), .ZN(new_n295));
  XOR2_X1   g094(.A(G141gat), .B(G148gat), .Z(new_n296));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT2), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n297), .A2(new_n301), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n297), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(new_n300), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n296), .B(new_n298), .C1(new_n306), .C2(new_n302), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n295), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI211_X1 g109(.A(KEYINPUT79), .B(KEYINPUT3), .C1(new_n304), .C2(new_n307), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n294), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT70), .B(G197gat), .ZN(new_n315));
  INV_X1    g114(.A(G204gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n323), .B1(new_n317), .B2(new_n321), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT84), .B(new_n294), .C1(new_n310), .C2(new_n311), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n314), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(G228gat), .A2(G233gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n294), .B1(new_n325), .B2(new_n326), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n309), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n304), .A2(new_n307), .A3(KEYINPUT78), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT78), .B1(new_n304), .B2(new_n307), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n331), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT85), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n329), .A2(new_n338), .A3(KEYINPUT85), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n312), .A2(new_n327), .ZN(new_n344));
  INV_X1    g143(.A(new_n333), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n345), .B2(new_n308), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n331), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n293), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n329), .A2(new_n338), .A3(KEYINPUT85), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT85), .B1(new_n329), .B2(new_n338), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n347), .B(new_n293), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n292), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G22gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(new_n351), .A3(new_n291), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n288), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n308), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(KEYINPUT3), .A3(new_n334), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n267), .C1(new_n310), .C2(new_n311), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n308), .A2(new_n265), .A3(new_n266), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT4), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n256), .A2(new_n365), .A3(new_n308), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT80), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n363), .B2(KEYINPUT4), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n361), .B(new_n362), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT5), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n359), .A2(new_n334), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n363), .B1(new_n372), .B2(new_n256), .ZN(new_n373));
  INV_X1    g172(.A(new_n362), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n371), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n256), .B1(new_n337), .B2(KEYINPUT3), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n310), .A2(new_n311), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT5), .B1(new_n364), .B2(new_n366), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  XOR2_X1   g181(.A(G1gat), .B(G29gat), .Z(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G57gat), .B(G85gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT6), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n376), .A2(new_n389), .A3(new_n381), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(KEYINPUT82), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT82), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n370), .A2(new_n375), .B1(new_n379), .B2(new_n380), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n388), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n393), .A2(new_n396), .A3(new_n389), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n239), .A2(new_n294), .ZN(new_n400));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT73), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT71), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n239), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n261), .A2(KEYINPUT71), .A3(new_n219), .ZN(new_n405));
  INV_X1    g204(.A(new_n401), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT73), .A4(new_n406), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n327), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n405), .A3(new_n294), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n401), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n239), .A2(KEYINPUT72), .A3(new_n406), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT72), .B1(new_n239), .B2(new_n406), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n327), .ZN(new_n419));
  XOR2_X1   g218(.A(G64gat), .B(G92gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT76), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n412), .A2(new_n419), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n327), .B1(new_n408), .B2(new_n409), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n411), .B1(new_n414), .B2(new_n417), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n425), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n419), .ZN(new_n433));
  INV_X1    g232(.A(new_n425), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n428), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n399), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n390), .A2(KEYINPUT82), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n393), .A2(new_n392), .A3(new_n389), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n397), .B1(new_n441), .B2(new_n388), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n428), .A2(new_n432), .A3(new_n435), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT83), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n357), .A2(new_n438), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT35), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT87), .B1(new_n393), .B2(new_n389), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n382), .A2(new_n448), .A3(new_n387), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n441), .A2(new_n396), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT35), .B(new_n443), .C1(new_n450), .C2(new_n398), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n357), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n285), .A2(KEYINPUT36), .A3(new_n287), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT36), .B1(new_n285), .B2(new_n287), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n364), .A2(new_n366), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n362), .B1(new_n361), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n387), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT39), .B1(new_n373), .B2(new_n374), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n462), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n459), .B(new_n464), .C1(new_n457), .C2(new_n460), .ZN(new_n465));
  AND4_X1   g264(.A1(new_n447), .A2(new_n463), .A3(new_n449), .A4(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n353), .A2(new_n356), .B1(new_n466), .B2(new_n443), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n434), .B1(new_n433), .B2(KEYINPUT37), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT37), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n431), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT38), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n425), .B1(new_n431), .B2(new_n469), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n410), .B2(new_n327), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n418), .A2(new_n411), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT38), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n472), .A2(new_n475), .B1(new_n431), .B2(new_n425), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n450), .A2(new_n471), .A3(new_n476), .A4(new_n398), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n455), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n353), .A2(new_n356), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n437), .B1(new_n399), .B2(new_n436), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT83), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n446), .A2(new_n452), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(G1gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT16), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n485), .A2(G1gat), .ZN(new_n489));
  OAI21_X1  g288(.A(G8gat), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n487), .ZN(new_n491));
  INV_X1    g290(.A(G8gat), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n491), .B(new_n492), .C1(G1gat), .C2(new_n485), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT88), .ZN(new_n497));
  INV_X1    g296(.A(G29gat), .ZN(new_n498));
  INV_X1    g297(.A(G36gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT14), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT14), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT15), .A4(new_n503), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n496), .B(new_n497), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT89), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(new_n511), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n494), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n521), .A2(KEYINPUT90), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT90), .B1(new_n521), .B2(new_n522), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n515), .A2(KEYINPUT18), .A3(new_n518), .A4(new_n520), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n494), .B(new_n519), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n517), .B(KEYINPUT13), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G197gat), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT11), .B(G169gat), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT12), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n526), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n522), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n529), .A3(new_n526), .ZN(new_n538));
  INV_X1    g337(.A(new_n534), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n525), .A2(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n484), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  INV_X1    g342(.A(G85gat), .ZN(new_n544));
  INV_X1    g343(.A(G92gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G99gat), .B(G106gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(G85gat), .A2(G92gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n546), .A2(new_n547), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT95), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n543), .A2(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n544), .A2(new_n545), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(new_n550), .A3(new_n556), .A4(new_n551), .ZN(new_n557));
  INV_X1    g356(.A(new_n547), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(new_n553), .A3(new_n552), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n542), .B1(new_n561), .B2(new_n519), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n562), .B(KEYINPUT96), .Z(new_n563));
  INV_X1    g362(.A(new_n561), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n513), .B2(new_n514), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n567), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G190gat), .B(G218gat), .Z(new_n571));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n568), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n568), .B2(new_n570), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G64gat), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n577), .A2(G57gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(G57gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G78gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT92), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(G71gat), .B2(G78gat), .ZN(new_n587));
  AND3_X1   g386(.A1(KEYINPUT91), .A2(G71gat), .A3(G78gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT91), .B1(G71gat), .B2(G78gat), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n585), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n581), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(KEYINPUT91), .A2(G71gat), .A3(G78gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(KEYINPUT93), .A3(new_n587), .A4(new_n585), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n582), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n581), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n490), .B(new_n493), .C1(new_n603), .C2(new_n604), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT94), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n609), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n576), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n582), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n585), .A2(new_n587), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT93), .B1(new_n621), .B2(new_n596), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n590), .A2(new_n591), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n624), .A2(new_n601), .A3(new_n554), .A4(new_n560), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n559), .A2(new_n552), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n598), .B2(new_n602), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n624), .B2(new_n601), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n561), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n619), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n618), .B1(new_n625), .B2(new_n628), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT97), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n636), .B1(new_n635), .B2(new_n640), .ZN(new_n643));
  INV_X1    g442(.A(new_n640), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT98), .B1(new_n634), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n634), .A2(KEYINPUT98), .A3(new_n644), .ZN(new_n646));
  OAI22_X1  g445(.A1(new_n642), .A2(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n617), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n541), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n442), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n443), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n649), .ZN(new_n654));
  OAI21_X1  g453(.A(G8gat), .B1(new_n654), .B2(new_n436), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n653), .ZN(new_n656));
  MUX2_X1   g455(.A(new_n653), .B(new_n656), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g456(.A(new_n455), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n288), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n654), .B2(new_n660), .ZN(G1326gat));
  NAND2_X1  g460(.A1(new_n649), .A2(new_n480), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n616), .A2(new_n647), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n525), .A2(new_n536), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n538), .A2(new_n539), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n484), .A2(new_n576), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n498), .A3(new_n442), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT45), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n484), .B2(new_n576), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n574), .A2(new_n575), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n478), .A2(new_n483), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n445), .A2(KEYINPUT35), .B1(new_n451), .B2(new_n357), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT44), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n669), .B(KEYINPUT100), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n674), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n674), .A2(new_n678), .A3(KEYINPUT101), .A4(new_n679), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n682), .A2(new_n442), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n672), .B1(new_n684), .B2(new_n498), .ZN(G1328gat));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n499), .A3(new_n443), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT46), .Z(new_n687));
  AND3_X1   g486(.A1(new_n682), .A2(new_n443), .A3(new_n683), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n499), .B2(new_n688), .ZN(G1329gat));
  INV_X1    g488(.A(new_n670), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(G43gat), .A3(new_n288), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G43gat), .B1(new_n680), .B2(new_n658), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n682), .A2(new_n455), .A3(new_n683), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n691), .B1(new_n696), .B2(G43gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n697), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g497(.A1(new_n576), .A2(G50gat), .ZN(new_n699));
  AND4_X1   g498(.A1(new_n480), .A2(new_n541), .A3(new_n665), .A4(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT48), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G50gat), .B1(new_n680), .B2(new_n479), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n682), .A2(new_n480), .A3(new_n683), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n705), .A2(new_n706), .A3(G50gat), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n705), .B2(G50gat), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n707), .A2(new_n708), .A3(new_n700), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n704), .B1(new_n709), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g509(.A(new_n647), .ZN(new_n711));
  NOR4_X1   g510(.A1(new_n484), .A2(new_n668), .A3(new_n617), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n442), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n443), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT49), .B(G64gat), .Z(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT103), .ZN(G1333gat));
  NAND3_X1  g518(.A1(new_n712), .A2(G71gat), .A3(new_n455), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT104), .ZN(new_n721));
  INV_X1    g520(.A(new_n288), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n712), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(G71gat), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g524(.A1(new_n712), .A2(new_n480), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n668), .A3(new_n616), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n674), .A2(new_n678), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n674), .A2(new_n678), .A3(KEYINPUT105), .A4(new_n728), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n731), .A2(new_n442), .A3(new_n732), .ZN(new_n733));
  OR4_X1    g532(.A1(new_n484), .A2(new_n668), .A3(new_n616), .A4(new_n576), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT51), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n442), .A2(new_n544), .A3(new_n647), .ZN(new_n736));
  OAI22_X1  g535(.A1(new_n733), .A2(new_n544), .B1(new_n735), .B2(new_n736), .ZN(G1336gat));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738));
  OAI21_X1  g537(.A(G92gat), .B1(new_n729), .B2(new_n436), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n443), .A2(new_n545), .A3(new_n647), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n738), .B(new_n739), .C1(new_n735), .C2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n731), .A2(new_n443), .A3(new_n732), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(new_n743), .A3(G92gat), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(G92gat), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n734), .A2(KEYINPUT107), .A3(KEYINPUT51), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n734), .B2(KEYINPUT107), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n746), .A2(new_n747), .A3(new_n740), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n741), .B1(new_n749), .B2(new_n738), .ZN(G1337gat));
  NAND3_X1  g549(.A1(new_n731), .A2(new_n455), .A3(new_n732), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G99gat), .ZN(new_n752));
  OR3_X1    g551(.A1(new_n288), .A2(new_n711), .A3(G99gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n735), .B2(new_n753), .ZN(G1338gat));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  OAI21_X1  g554(.A(G106gat), .B1(new_n729), .B2(new_n479), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n479), .A2(G106gat), .A3(new_n711), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n755), .B(new_n756), .C1(new_n735), .C2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n746), .A2(new_n747), .A3(new_n757), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n731), .A2(new_n480), .A3(new_n732), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(G106gat), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n761), .B2(new_n755), .ZN(G1339gat));
  NOR3_X1   g561(.A1(new_n617), .A2(new_n668), .A3(new_n647), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n646), .A2(new_n645), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n644), .B1(new_n632), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n629), .A2(new_n631), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n765), .B1(new_n768), .B2(new_n618), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n618), .B1(new_n630), .B2(new_n561), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n629), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n629), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT108), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n769), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT109), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n770), .A2(new_n771), .A3(new_n629), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n771), .B1(new_n770), .B2(new_n629), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n769), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n767), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n764), .B1(new_n782), .B2(KEYINPUT55), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n779), .B2(new_n769), .ZN(new_n784));
  AND4_X1   g583(.A1(new_n780), .A2(new_n769), .A3(new_n772), .A4(new_n774), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n766), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n523), .A2(new_n524), .A3(new_n535), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n518), .B1(new_n515), .B2(new_n520), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n790), .A2(new_n791), .B1(new_n527), .B2(new_n528), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n533), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(KEYINPUT111), .B(new_n533), .C1(new_n792), .C2(new_n793), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n789), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n788), .A3(new_n675), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n540), .B1(new_n786), .B2(new_n787), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n800), .A2(new_n783), .B1(new_n647), .B2(new_n798), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n801), .B2(new_n675), .ZN(new_n802));
  INV_X1    g601(.A(new_n616), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT112), .B(new_n763), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n783), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n798), .A2(new_n647), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n675), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n799), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n763), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n804), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n480), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n399), .A2(new_n443), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n722), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n246), .A3(new_n540), .ZN(new_n817));
  INV_X1    g616(.A(new_n357), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n813), .A2(new_n399), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n819), .A2(KEYINPUT113), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(KEYINPUT113), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n436), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(new_n540), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n817), .B1(new_n823), .B2(new_n246), .ZN(G1340gat));
  OAI21_X1  g623(.A(G120gat), .B1(new_n816), .B2(new_n711), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n711), .A2(new_n248), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT114), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n822), .B2(new_n827), .ZN(G1341gat));
  OAI21_X1  g627(.A(new_n244), .B1(new_n816), .B2(new_n803), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n803), .A2(new_n244), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n822), .B2(new_n830), .ZN(G1342gat));
  NOR2_X1   g630(.A1(new_n576), .A2(G134gat), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OR3_X1    g632(.A1(new_n822), .A2(KEYINPUT56), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n816), .B2(new_n576), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT56), .B1(new_n822), .B2(new_n833), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n658), .A2(new_n815), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n786), .A2(new_n787), .B1(new_n645), .B2(new_n646), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n668), .B1(new_n782), .B2(KEYINPUT55), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n807), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n576), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n616), .B1(new_n843), .B2(new_n799), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT112), .B1(new_n844), .B2(new_n763), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n763), .B1(new_n802), .B2(new_n803), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n805), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n848), .B2(new_n480), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n479), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT115), .B(new_n852), .C1(new_n844), .C2(new_n763), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n839), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G141gat), .B1(new_n857), .B2(new_n540), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n455), .A2(new_n479), .A3(new_n443), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n848), .A2(new_n442), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(G141gat), .A3(new_n540), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(KEYINPUT58), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n480), .B1(new_n804), .B2(new_n812), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n856), .B1(new_n851), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT116), .B1(new_n865), .B2(new_n838), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n867), .B(new_n839), .C1(new_n849), .C2(new_n856), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n668), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n861), .B1(new_n869), .B2(G141gat), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(G1344gat));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n647), .A3(new_n868), .ZN(new_n873));
  INV_X1    g672(.A(G148gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(KEYINPUT59), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(KEYINPUT117), .A3(new_n875), .ZN(new_n879));
  XOR2_X1   g678(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n880));
  XNOR2_X1  g679(.A(new_n763), .B(KEYINPUT119), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n851), .B(new_n480), .C1(new_n881), .C2(new_n844), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n838), .A2(new_n711), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n479), .B1(new_n845), .B2(new_n847), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n851), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n880), .B1(new_n885), .B2(G148gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n878), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n860), .A2(G148gat), .A3(new_n711), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1345gat));
  NAND4_X1  g690(.A1(new_n866), .A2(G155gat), .A3(new_n616), .A4(new_n868), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n860), .A2(new_n803), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(G155gat), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT121), .ZN(G1346gat));
  NOR3_X1   g694(.A1(new_n860), .A2(G162gat), .A3(new_n576), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT122), .Z(new_n897));
  INV_X1    g696(.A(G162gat), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n866), .A2(new_n675), .A3(new_n868), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n436), .A2(new_n442), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n479), .A2(new_n848), .A3(new_n722), .A4(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(G169gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(new_n540), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n813), .A2(new_n442), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT123), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n818), .A2(new_n436), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(new_n668), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n909), .B2(new_n904), .ZN(G1348gat));
  NAND3_X1  g709(.A1(new_n902), .A2(G176gat), .A3(new_n647), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT124), .ZN(new_n912));
  INV_X1    g711(.A(G176gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n907), .A2(new_n647), .A3(new_n908), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(G1349gat));
  NAND2_X1  g714(.A1(new_n902), .A2(new_n616), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT125), .B1(new_n916), .B2(G183gat), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n907), .A2(new_n908), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n616), .A2(new_n206), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n920), .B(new_n922), .ZN(G1350gat));
  AOI21_X1  g722(.A(new_n207), .B1(new_n902), .B2(new_n675), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT61), .Z(new_n925));
  NAND2_X1  g724(.A1(new_n675), .A2(new_n207), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n918), .B2(new_n926), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n864), .A2(KEYINPUT57), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n928), .A2(new_n658), .A3(new_n882), .A4(new_n901), .ZN(new_n929));
  INV_X1    g728(.A(G197gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(new_n540), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n455), .A2(new_n479), .A3(new_n436), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n907), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n668), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n930), .ZN(G1352gat));
  NOR2_X1   g735(.A1(new_n711), .A2(G204gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n929), .B2(new_n711), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(G1353gat));
  NAND3_X1  g742(.A1(new_n934), .A2(new_n319), .A3(new_n616), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n929), .A2(new_n803), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1354gat));
  OAI21_X1  g748(.A(G218gat), .B1(new_n929), .B2(new_n576), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n576), .A2(G218gat), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n933), .B2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(G1355gat));
endmodule


