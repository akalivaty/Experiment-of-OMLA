

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n733), .A2(n732), .ZN(n721) );
  NOR2_X1 U554 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U555 ( .A1(G8), .A2(n726), .ZN(n761) );
  INV_X1 U556 ( .A(G651), .ZN(n527) );
  INV_X2 U557 ( .A(n670), .ZN(n774) );
  NOR2_X2 U558 ( .A1(n679), .A2(n678), .ZN(n684) );
  NOR2_X4 U559 ( .A1(G2105), .A2(n543), .ZN(n907) );
  NAND2_X1 U560 ( .A1(n642), .A2(n641), .ZN(n726) );
  BUF_X1 U561 ( .A(n647), .Z(n520) );
  NOR2_X1 U562 ( .A1(G543), .A2(n527), .ZN(n529) );
  XOR2_X2 U563 ( .A(n656), .B(n655), .Z(n670) );
  NOR2_X4 U564 ( .A1(n586), .A2(n527), .ZN(n645) );
  XOR2_X2 U565 ( .A(KEYINPUT0), .B(G543), .Z(n586) );
  XNOR2_X1 U566 ( .A(n529), .B(n528), .ZN(n647) );
  NAND2_X1 U567 ( .A1(n522), .A2(n993), .ZN(n750) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  NOR2_X2 U569 ( .A1(n557), .A2(n556), .ZN(G160) );
  XOR2_X1 U570 ( .A(n649), .B(n648), .Z(n521) );
  OR2_X1 U571 ( .A1(n749), .A2(n761), .ZN(n522) );
  INV_X1 U572 ( .A(KEYINPUT103), .ZN(n685) );
  XNOR2_X1 U573 ( .A(n714), .B(KEYINPUT30), .ZN(n715) );
  INV_X1 U574 ( .A(KEYINPUT29), .ZN(n706) );
  INV_X1 U575 ( .A(KEYINPUT66), .ZN(n540) );
  OR2_X1 U576 ( .A1(n751), .A2(n750), .ZN(n758) );
  AND2_X1 U577 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U578 ( .A(n540), .B(KEYINPUT17), .ZN(n541) );
  XNOR2_X1 U579 ( .A(n542), .B(n541), .ZN(n551) );
  BUF_X1 U580 ( .A(n551), .Z(n908) );
  XNOR2_X1 U581 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n769) );
  NOR2_X1 U582 ( .A1(n548), .A2(n547), .ZN(G164) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n796) );
  NAND2_X1 U584 ( .A1(n796), .A2(G89), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(KEYINPUT4), .ZN(n525) );
  NAND2_X1 U586 ( .A1(G76), .A2(n645), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U588 ( .A(KEYINPUT5), .B(n526), .ZN(n535) );
  XNOR2_X1 U589 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n528) );
  NAND2_X1 U590 ( .A1(G63), .A2(n520), .ZN(n531) );
  NOR2_X4 U591 ( .A1(G651), .A2(n586), .ZN(n799) );
  NAND2_X1 U592 ( .A1(G51), .A2(n799), .ZN(n530) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n533) );
  XOR2_X1 U594 ( .A(KEYINPUT82), .B(KEYINPUT6), .Z(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U597 ( .A(KEYINPUT7), .B(n536), .ZN(G168) );
  INV_X1 U598 ( .A(G2104), .ZN(n543) );
  AND2_X1 U599 ( .A1(n543), .A2(G2105), .ZN(n902) );
  NAND2_X1 U600 ( .A1(G126), .A2(n902), .ZN(n538) );
  AND2_X1 U601 ( .A1(G2104), .A2(G2105), .ZN(n903) );
  NAND2_X1 U602 ( .A1(G114), .A2(n903), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(KEYINPUT96), .B(n539), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n551), .A2(G138), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G102), .A2(n907), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT97), .B(n546), .Z(n547) );
  NAND2_X1 U609 ( .A1(G101), .A2(n907), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n549), .B(KEYINPUT65), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT23), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G137), .A2(n908), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G125), .A2(n902), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G113), .A2(n903), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G72), .A2(n645), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G85), .A2(n796), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G60), .A2(n520), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G47), .A2(n799), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U623 ( .A1(n563), .A2(n562), .ZN(G290) );
  XNOR2_X1 U624 ( .A(KEYINPUT9), .B(KEYINPUT71), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G77), .A2(n645), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G90), .A2(n796), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U628 ( .A(n567), .B(n566), .ZN(n574) );
  NAND2_X1 U629 ( .A1(n799), .A2(G52), .ZN(n568) );
  XNOR2_X1 U630 ( .A(KEYINPUT69), .B(n568), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n520), .A2(G64), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT68), .B(n569), .Z(n570) );
  NOR2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT70), .B(n572), .Z(n573) );
  NOR2_X1 U635 ( .A1(n574), .A2(n573), .ZN(G171) );
  NAND2_X1 U636 ( .A1(n799), .A2(G50), .ZN(n581) );
  NAND2_X1 U637 ( .A1(G75), .A2(n645), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G62), .A2(n520), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G88), .A2(n796), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT87), .B(n577), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U644 ( .A(KEYINPUT88), .B(n582), .ZN(G303) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(G49), .A2(n799), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G74), .A2(G651), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U649 ( .A1(n520), .A2(n585), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n586), .A2(G87), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(G288) );
  NAND2_X1 U652 ( .A1(G86), .A2(n796), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G61), .A2(n520), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G73), .A2(n645), .ZN(n591) );
  XOR2_X1 U656 ( .A(KEYINPUT2), .B(n591), .Z(n592) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U658 ( .A1(n799), .A2(G48), .ZN(n594) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(G305) );
  INV_X1 U660 ( .A(G303), .ZN(G166) );
  NOR2_X1 U661 ( .A1(G164), .A2(G1384), .ZN(n596) );
  XNOR2_X1 U662 ( .A(KEYINPUT64), .B(n596), .ZN(n641) );
  NAND2_X1 U663 ( .A1(G40), .A2(G160), .ZN(n597) );
  XOR2_X1 U664 ( .A(KEYINPUT98), .B(n597), .Z(n642) );
  INV_X1 U665 ( .A(n642), .ZN(n598) );
  NOR2_X1 U666 ( .A1(n641), .A2(n598), .ZN(n636) );
  INV_X1 U667 ( .A(n636), .ZN(n633) );
  XNOR2_X1 U668 ( .A(G2067), .B(KEYINPUT37), .ZN(n608) );
  NAND2_X1 U669 ( .A1(G128), .A2(n902), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G116), .A2(n903), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n601), .B(KEYINPUT35), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G104), .A2(n907), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G140), .A2(n908), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT34), .B(n604), .Z(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U678 ( .A(n607), .B(KEYINPUT36), .Z(n884) );
  AND2_X1 U679 ( .A1(n608), .A2(n884), .ZN(n952) );
  NOR2_X1 U680 ( .A1(n608), .A2(n884), .ZN(n946) );
  XOR2_X1 U681 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n629) );
  NAND2_X1 U682 ( .A1(G129), .A2(n902), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G141), .A2(n908), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n907), .A2(G105), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT38), .B(n611), .Z(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n903), .A2(G117), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n881) );
  NOR2_X1 U690 ( .A1(G1996), .A2(n881), .ZN(n930) );
  NAND2_X1 U691 ( .A1(G95), .A2(n907), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G131), .A2(n908), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G119), .A2(n902), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G107), .A2(n903), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n886) );
  AND2_X1 U698 ( .A1(n886), .A2(G1991), .ZN(n623) );
  AND2_X1 U699 ( .A1(n881), .A2(G1996), .ZN(n622) );
  NOR2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n933) );
  NOR2_X1 U701 ( .A1(n933), .A2(n633), .ZN(n638) );
  NOR2_X1 U702 ( .A1(G1986), .A2(G290), .ZN(n625) );
  NOR2_X1 U703 ( .A1(G1991), .A2(n886), .ZN(n624) );
  XNOR2_X1 U704 ( .A(KEYINPUT106), .B(n624), .ZN(n941) );
  NOR2_X1 U705 ( .A1(n625), .A2(n941), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n638), .A2(n626), .ZN(n627) );
  NOR2_X1 U707 ( .A1(n930), .A2(n627), .ZN(n628) );
  XOR2_X1 U708 ( .A(n629), .B(n628), .Z(n630) );
  NOR2_X1 U709 ( .A1(n946), .A2(n630), .ZN(n631) );
  NOR2_X1 U710 ( .A1(n952), .A2(n631), .ZN(n632) );
  NOR2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n634), .B(KEYINPUT108), .ZN(n768) );
  INV_X1 U713 ( .A(n946), .ZN(n635) );
  XOR2_X1 U714 ( .A(G1986), .B(G290), .Z(n980) );
  NAND2_X1 U715 ( .A1(n635), .A2(n980), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n640) );
  INV_X1 U717 ( .A(n638), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n766) );
  NOR2_X1 U719 ( .A1(G1966), .A2(n761), .ZN(n722) );
  XNOR2_X1 U720 ( .A(KEYINPUT15), .B(KEYINPUT81), .ZN(n656) );
  NAND2_X1 U721 ( .A1(G92), .A2(n796), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n643), .B(KEYINPUT78), .ZN(n654) );
  NAND2_X1 U723 ( .A1(G54), .A2(n799), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(KEYINPUT80), .ZN(n652) );
  NAND2_X1 U725 ( .A1(G79), .A2(n645), .ZN(n646) );
  XNOR2_X1 U726 ( .A(KEYINPUT79), .B(n646), .ZN(n650) );
  INV_X1 U727 ( .A(KEYINPUT77), .ZN(n649) );
  NAND2_X1 U728 ( .A1(G66), .A2(n647), .ZN(n648) );
  NOR2_X1 U729 ( .A1(n650), .A2(n521), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U731 ( .A1(G2067), .A2(n774), .ZN(n658) );
  XNOR2_X1 U732 ( .A(KEYINPUT26), .B(KEYINPUT102), .ZN(n677) );
  NAND2_X1 U733 ( .A1(G1996), .A2(n677), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n659), .A2(n688), .ZN(n676) );
  NAND2_X1 U736 ( .A1(n520), .A2(G56), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT14), .B(n660), .Z(n666) );
  NAND2_X1 U738 ( .A1(n796), .A2(G81), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(KEYINPUT12), .ZN(n663) );
  NAND2_X1 U740 ( .A1(G68), .A2(n645), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U742 ( .A(KEYINPUT13), .B(n664), .Z(n665) );
  NOR2_X1 U743 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n667), .B(KEYINPUT76), .ZN(n669) );
  NAND2_X1 U745 ( .A1(G43), .A2(n799), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n669), .A2(n668), .ZN(n1000) );
  NAND2_X1 U747 ( .A1(G1348), .A2(n774), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n671), .A2(n677), .ZN(n672) );
  NOR2_X1 U749 ( .A1(G1341), .A2(n672), .ZN(n673) );
  NOR2_X1 U750 ( .A1(n688), .A2(n673), .ZN(n674) );
  NOR2_X1 U751 ( .A1(n1000), .A2(n674), .ZN(n675) );
  NAND2_X1 U752 ( .A1(n676), .A2(n675), .ZN(n679) );
  NOR2_X1 U753 ( .A1(G1996), .A2(n677), .ZN(n678) );
  NAND2_X1 U754 ( .A1(G1348), .A2(n726), .ZN(n681) );
  INV_X1 U755 ( .A(n726), .ZN(n688) );
  NAND2_X1 U756 ( .A1(n688), .A2(G2067), .ZN(n680) );
  NAND2_X1 U757 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U758 ( .A1(n682), .A2(n774), .ZN(n683) );
  NOR2_X1 U759 ( .A1(n684), .A2(n683), .ZN(n686) );
  XNOR2_X1 U760 ( .A(n686), .B(n685), .ZN(n701) );
  NAND2_X1 U761 ( .A1(G1956), .A2(n726), .ZN(n687) );
  XNOR2_X1 U762 ( .A(KEYINPUT101), .B(n687), .ZN(n691) );
  NAND2_X1 U763 ( .A1(n688), .A2(G2072), .ZN(n689) );
  XNOR2_X1 U764 ( .A(KEYINPUT27), .B(n689), .ZN(n690) );
  NOR2_X1 U765 ( .A1(n691), .A2(n690), .ZN(n702) );
  NAND2_X1 U766 ( .A1(G65), .A2(n520), .ZN(n693) );
  NAND2_X1 U767 ( .A1(G53), .A2(n799), .ZN(n692) );
  NAND2_X1 U768 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U769 ( .A(n694), .B(KEYINPUT73), .ZN(n696) );
  NAND2_X1 U770 ( .A1(G78), .A2(n645), .ZN(n695) );
  NAND2_X1 U771 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U772 ( .A1(n796), .A2(G91), .ZN(n697) );
  XOR2_X1 U773 ( .A(KEYINPUT72), .B(n697), .Z(n698) );
  NOR2_X1 U774 ( .A1(n699), .A2(n698), .ZN(n979) );
  NAND2_X1 U775 ( .A1(n702), .A2(n979), .ZN(n700) );
  NAND2_X1 U776 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U777 ( .A1(n702), .A2(n979), .ZN(n703) );
  XOR2_X1 U778 ( .A(n703), .B(KEYINPUT28), .Z(n704) );
  NAND2_X1 U779 ( .A1(n705), .A2(n704), .ZN(n707) );
  XNOR2_X1 U780 ( .A(n707), .B(n706), .ZN(n712) );
  INV_X1 U781 ( .A(G1961), .ZN(n863) );
  NAND2_X1 U782 ( .A1(n726), .A2(n863), .ZN(n709) );
  XNOR2_X1 U783 ( .A(G2078), .B(KEYINPUT25), .ZN(n958) );
  NAND2_X1 U784 ( .A1(n688), .A2(n958), .ZN(n708) );
  NAND2_X1 U785 ( .A1(n709), .A2(n708), .ZN(n716) );
  AND2_X1 U786 ( .A1(n716), .A2(G171), .ZN(n710) );
  XOR2_X1 U787 ( .A(KEYINPUT100), .B(n710), .Z(n711) );
  NAND2_X1 U788 ( .A1(n712), .A2(n711), .ZN(n733) );
  NOR2_X1 U789 ( .A1(G2084), .A2(n726), .ZN(n723) );
  NOR2_X1 U790 ( .A1(n722), .A2(n723), .ZN(n713) );
  NAND2_X1 U791 ( .A1(G8), .A2(n713), .ZN(n714) );
  NOR2_X1 U792 ( .A1(n715), .A2(G168), .ZN(n718) );
  NOR2_X1 U793 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U794 ( .A1(n718), .A2(n717), .ZN(n720) );
  INV_X1 U795 ( .A(KEYINPUT31), .ZN(n719) );
  XNOR2_X1 U796 ( .A(n720), .B(n719), .ZN(n732) );
  NAND2_X1 U797 ( .A1(G8), .A2(n723), .ZN(n724) );
  NAND2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n741) );
  INV_X1 U799 ( .A(G8), .ZN(n731) );
  NOR2_X1 U800 ( .A1(G2090), .A2(n726), .ZN(n728) );
  NOR2_X1 U801 ( .A1(G1971), .A2(n761), .ZN(n727) );
  NOR2_X1 U802 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U803 ( .A1(G303), .A2(n729), .ZN(n730) );
  OR2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n735) );
  AND2_X1 U805 ( .A1(n732), .A2(n735), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n734), .A2(n733), .ZN(n738) );
  INV_X1 U807 ( .A(n735), .ZN(n736) );
  OR2_X1 U808 ( .A1(n736), .A2(G286), .ZN(n737) );
  NAND2_X1 U809 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U810 ( .A(n739), .B(KEYINPUT32), .ZN(n740) );
  NAND2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U812 ( .A(KEYINPUT104), .B(n742), .Z(n754) );
  NOR2_X1 U813 ( .A1(G303), .A2(G1971), .ZN(n743) );
  NOR2_X1 U814 ( .A1(G1976), .A2(G288), .ZN(n982) );
  OR2_X1 U815 ( .A1(n743), .A2(n982), .ZN(n744) );
  NOR2_X1 U816 ( .A1(n754), .A2(n744), .ZN(n747) );
  NAND2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n983) );
  INV_X1 U818 ( .A(n761), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n983), .A2(n745), .ZN(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U821 ( .A1(n748), .A2(KEYINPUT33), .ZN(n751) );
  NAND2_X1 U822 ( .A1(n982), .A2(KEYINPUT33), .ZN(n749) );
  XOR2_X1 U823 ( .A(G1981), .B(G305), .Z(n993) );
  NAND2_X1 U824 ( .A1(G8), .A2(G166), .ZN(n752) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n752), .ZN(n753) );
  NOR2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U827 ( .A(KEYINPUT105), .B(n755), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n756), .A2(n761), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n764) );
  NOR2_X1 U830 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U831 ( .A(n759), .B(KEYINPUT24), .Z(n760) );
  NOR2_X1 U832 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U833 ( .A(KEYINPUT99), .B(n762), .Z(n763) );
  NOR2_X1 U834 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U835 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U836 ( .A1(n768), .A2(n767), .ZN(n770) );
  XNOR2_X1 U837 ( .A(n770), .B(n769), .ZN(G329) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U839 ( .A(G57), .ZN(G237) );
  XOR2_X1 U840 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n772) );
  NAND2_X1 U841 ( .A1(G7), .A2(G661), .ZN(n771) );
  XOR2_X1 U842 ( .A(n772), .B(n771), .Z(n837) );
  NAND2_X1 U843 ( .A1(n837), .A2(G567), .ZN(n773) );
  XOR2_X1 U844 ( .A(KEYINPUT11), .B(n773), .Z(G234) );
  INV_X1 U845 ( .A(G860), .ZN(n779) );
  OR2_X1 U846 ( .A1(n1000), .A2(n779), .ZN(G153) );
  INV_X1 U847 ( .A(G171), .ZN(G301) );
  NAND2_X1 U848 ( .A1(G868), .A2(G301), .ZN(n776) );
  INV_X1 U849 ( .A(G868), .ZN(n817) );
  NAND2_X1 U850 ( .A1(n774), .A2(n817), .ZN(n775) );
  NAND2_X1 U851 ( .A1(n776), .A2(n775), .ZN(G284) );
  XOR2_X1 U852 ( .A(n979), .B(KEYINPUT74), .Z(G299) );
  NOR2_X1 U853 ( .A1(G299), .A2(G868), .ZN(n778) );
  NOR2_X1 U854 ( .A1(G286), .A2(n817), .ZN(n777) );
  NOR2_X1 U855 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U856 ( .A1(n779), .A2(G559), .ZN(n780) );
  NAND2_X1 U857 ( .A1(n780), .A2(n670), .ZN(n781) );
  XNOR2_X1 U858 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U859 ( .A1(G868), .A2(n1000), .ZN(n784) );
  NAND2_X1 U860 ( .A1(G868), .A2(n670), .ZN(n782) );
  NOR2_X1 U861 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U862 ( .A1(n784), .A2(n783), .ZN(G282) );
  NAND2_X1 U863 ( .A1(G123), .A2(n902), .ZN(n785) );
  XOR2_X1 U864 ( .A(KEYINPUT18), .B(n785), .Z(n786) );
  XNOR2_X1 U865 ( .A(n786), .B(KEYINPUT83), .ZN(n788) );
  NAND2_X1 U866 ( .A1(G135), .A2(n908), .ZN(n787) );
  NAND2_X1 U867 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U868 ( .A(KEYINPUT84), .B(n789), .ZN(n793) );
  NAND2_X1 U869 ( .A1(G99), .A2(n907), .ZN(n791) );
  NAND2_X1 U870 ( .A1(G111), .A2(n903), .ZN(n790) );
  NAND2_X1 U871 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U872 ( .A1(n793), .A2(n792), .ZN(n942) );
  XNOR2_X1 U873 ( .A(n942), .B(G2096), .ZN(n794) );
  INV_X1 U874 ( .A(G2100), .ZN(n854) );
  NAND2_X1 U875 ( .A1(n794), .A2(n854), .ZN(G156) );
  NAND2_X1 U876 ( .A1(G559), .A2(n670), .ZN(n795) );
  XNOR2_X1 U877 ( .A(n1000), .B(n795), .ZN(n815) );
  NOR2_X1 U878 ( .A1(n815), .A2(G860), .ZN(n806) );
  NAND2_X1 U879 ( .A1(G80), .A2(n645), .ZN(n798) );
  NAND2_X1 U880 ( .A1(G93), .A2(n796), .ZN(n797) );
  NAND2_X1 U881 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U882 ( .A1(G55), .A2(n799), .ZN(n800) );
  XNOR2_X1 U883 ( .A(KEYINPUT85), .B(n800), .ZN(n801) );
  NOR2_X1 U884 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U885 ( .A1(n520), .A2(G67), .ZN(n803) );
  NAND2_X1 U886 ( .A1(n804), .A2(n803), .ZN(n818) );
  XOR2_X1 U887 ( .A(n818), .B(KEYINPUT86), .Z(n805) );
  XNOR2_X1 U888 ( .A(n806), .B(n805), .ZN(G145) );
  XOR2_X1 U889 ( .A(G166), .B(G299), .Z(n814) );
  XOR2_X1 U890 ( .A(KEYINPUT19), .B(KEYINPUT89), .Z(n808) );
  XNOR2_X1 U891 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n807) );
  XNOR2_X1 U892 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U893 ( .A(n809), .B(G288), .ZN(n810) );
  XNOR2_X1 U894 ( .A(n810), .B(n818), .ZN(n811) );
  XNOR2_X1 U895 ( .A(n811), .B(G305), .ZN(n812) );
  XNOR2_X1 U896 ( .A(n812), .B(G290), .ZN(n813) );
  XNOR2_X1 U897 ( .A(n814), .B(n813), .ZN(n919) );
  XNOR2_X1 U898 ( .A(n919), .B(n815), .ZN(n816) );
  NOR2_X1 U899 ( .A1(n817), .A2(n816), .ZN(n820) );
  NOR2_X1 U900 ( .A1(G868), .A2(n818), .ZN(n819) );
  NOR2_X1 U901 ( .A1(n820), .A2(n819), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U903 ( .A(KEYINPUT92), .B(KEYINPUT20), .Z(n821) );
  XNOR2_X1 U904 ( .A(n822), .B(n821), .ZN(n823) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U906 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U907 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U908 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n827) );
  NAND2_X1 U910 ( .A1(G132), .A2(G82), .ZN(n826) );
  XNOR2_X1 U911 ( .A(n827), .B(n826), .ZN(n828) );
  NOR2_X1 U912 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U913 ( .A1(G96), .A2(n829), .ZN(n830) );
  XNOR2_X1 U914 ( .A(KEYINPUT94), .B(n830), .ZN(n843) );
  NAND2_X1 U915 ( .A1(n843), .A2(G2106), .ZN(n834) );
  NAND2_X1 U916 ( .A1(G69), .A2(G120), .ZN(n831) );
  NOR2_X1 U917 ( .A1(G237), .A2(n831), .ZN(n832) );
  NAND2_X1 U918 ( .A1(G108), .A2(n832), .ZN(n842) );
  NAND2_X1 U919 ( .A1(G567), .A2(n842), .ZN(n833) );
  NAND2_X1 U920 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U921 ( .A(n835), .B(KEYINPUT95), .Z(n841) );
  NAND2_X1 U922 ( .A1(G661), .A2(G483), .ZN(n836) );
  NOR2_X1 U923 ( .A1(n841), .A2(n836), .ZN(n840) );
  NAND2_X1 U924 ( .A1(n840), .A2(G36), .ZN(G176) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n837), .ZN(G217) );
  INV_X1 U926 ( .A(n837), .ZN(G223) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U928 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U931 ( .A(n841), .ZN(G319) );
  INV_X1 U933 ( .A(G132), .ZN(G219) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G82), .ZN(G220) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U940 ( .A(G1341), .B(G2454), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n844), .B(G2430), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n845), .B(G1348), .ZN(n851) );
  XOR2_X1 U943 ( .A(G2443), .B(G2427), .Z(n847) );
  XNOR2_X1 U944 ( .A(G2438), .B(G2446), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n849) );
  XOR2_X1 U946 ( .A(G2451), .B(G2435), .Z(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  NAND2_X1 U949 ( .A1(n852), .A2(G14), .ZN(n853) );
  XOR2_X1 U950 ( .A(KEYINPUT110), .B(n853), .Z(G401) );
  XNOR2_X1 U951 ( .A(n854), .B(G2096), .ZN(n856) );
  XNOR2_X1 U952 ( .A(KEYINPUT42), .B(G2678), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U954 ( .A(KEYINPUT43), .B(G2090), .Z(n858) );
  XNOR2_X1 U955 ( .A(G2072), .B(G2067), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2084), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(G227) );
  XNOR2_X1 U960 ( .A(n863), .B(G1956), .ZN(n865) );
  XNOR2_X1 U961 ( .A(G1971), .B(G1966), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U963 ( .A(n866), .B(G2474), .Z(n868) );
  XNOR2_X1 U964 ( .A(G1996), .B(G1991), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U966 ( .A(KEYINPUT41), .B(G1986), .Z(n870) );
  XNOR2_X1 U967 ( .A(G1981), .B(G1976), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(G229) );
  NAND2_X1 U970 ( .A1(G124), .A2(n902), .ZN(n873) );
  XOR2_X1 U971 ( .A(KEYINPUT44), .B(n873), .Z(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(KEYINPUT111), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G100), .A2(n907), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U975 ( .A1(n903), .A2(G112), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G136), .A2(n908), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(G162) );
  XOR2_X1 U979 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n883) );
  XOR2_X1 U980 ( .A(n881), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n888) );
  XOR2_X1 U983 ( .A(G164), .B(n886), .Z(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(G162), .Z(n901) );
  NAND2_X1 U986 ( .A1(G139), .A2(n908), .ZN(n890) );
  XNOR2_X1 U987 ( .A(KEYINPUT115), .B(n890), .ZN(n899) );
  XOR2_X1 U988 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n891) );
  XNOR2_X1 U989 ( .A(KEYINPUT47), .B(n891), .ZN(n895) );
  NAND2_X1 U990 ( .A1(G127), .A2(n902), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G115), .A2(n903), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G103), .A2(n907), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  NOR2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n935) );
  XNOR2_X1 U997 ( .A(G160), .B(n935), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n917) );
  NAND2_X1 U999 ( .A1(G130), .A2(n902), .ZN(n905) );
  NAND2_X1 U1000 ( .A1(G118), .A2(n903), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(KEYINPUT112), .B(n906), .ZN(n914) );
  NAND2_X1 U1003 ( .A1(G106), .A2(n907), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(G142), .A2(n908), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT113), .B(n911), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(KEYINPUT45), .B(n912), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n942), .B(n915), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n918), .ZN(G395) );
  XNOR2_X1 U1012 ( .A(G286), .B(n919), .ZN(n921) );
  XOR2_X1 U1013 ( .A(n670), .B(G171), .Z(n920) );
  XNOR2_X1 U1014 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1015 ( .A(n922), .B(n1000), .ZN(n923) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n923), .ZN(G397) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n924), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n925), .ZN(n926) );
  AND2_X1 U1020 ( .A1(G319), .A2(n926), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT120), .B(n931), .Z(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT51), .B(n932), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1030 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n950) );
  XNOR2_X1 U1035 ( .A(G160), .B(G2084), .ZN(n944) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT118), .B(n945), .ZN(n947) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1040 ( .A(KEYINPUT119), .B(n948), .Z(n949) );
  NAND2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1043 ( .A(KEYINPUT121), .B(n953), .Z(n954) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n954), .ZN(n955) );
  XOR2_X1 U1045 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n975) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n975), .ZN(n956) );
  NAND2_X1 U1047 ( .A1(n956), .A2(G29), .ZN(n1034) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n970) );
  XOR2_X1 U1049 ( .A(G2072), .B(G33), .Z(n957) );
  NAND2_X1 U1050 ( .A1(n957), .A2(G28), .ZN(n967) );
  XNOR2_X1 U1051 ( .A(n958), .B(G27), .ZN(n960) );
  XOR2_X1 U1052 ( .A(G1996), .B(G32), .Z(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT123), .B(n961), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(G2067), .B(G26), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G25), .B(G1991), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(KEYINPUT53), .B(n968), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1062 ( .A(G2084), .B(G34), .Z(n971) );
  XNOR2_X1 U1063 ( .A(KEYINPUT54), .B(n971), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n975), .B(n974), .ZN(n977) );
  INV_X1 U1066 ( .A(G29), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(G11), .A2(n978), .ZN(n1032) );
  INV_X1 U1069 ( .A(G16), .ZN(n1028) );
  XOR2_X1 U1070 ( .A(n1028), .B(KEYINPUT56), .Z(n1004) );
  XNOR2_X1 U1071 ( .A(n979), .B(G1956), .ZN(n989) );
  XOR2_X1 U1072 ( .A(G1971), .B(G303), .Z(n981) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n987) );
  INV_X1 U1074 ( .A(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1076 ( .A(KEYINPUT125), .B(n985), .Z(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n999) );
  XOR2_X1 U1079 ( .A(n670), .B(G1348), .Z(n991) );
  XOR2_X1 U1080 ( .A(G171), .B(G1961), .Z(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT124), .B(n992), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G168), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(KEYINPUT57), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1088 ( .A(G1341), .B(n1000), .Z(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1030) );
  XOR2_X1 U1091 ( .A(G1961), .B(KEYINPUT126), .Z(n1005) );
  XNOR2_X1 U1092 ( .A(n1005), .B(G5), .ZN(n1015) );
  XOR2_X1 U1093 ( .A(G1348), .B(KEYINPUT59), .Z(n1006) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1006), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G20), .B(G1956), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1981), .B(G6), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1013), .Z(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XNOR2_X1 U1103 ( .A(G1971), .B(G22), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G24), .B(G1986), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(G1976), .B(G23), .Z(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(G1966), .B(G21), .Z(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(n1025), .B(KEYINPUT127), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1035), .ZN(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

