

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740;

  XNOR2_X1 U365 ( .A(n582), .B(n581), .ZN(n740) );
  XNOR2_X2 U366 ( .A(n724), .B(G146), .ZN(n523) );
  BUF_X1 U367 ( .A(n664), .Z(n344) );
  NOR2_X2 U368 ( .A1(n542), .A2(n358), .ZN(n520) );
  XNOR2_X2 U369 ( .A(n406), .B(KEYINPUT0), .ZN(n542) );
  XNOR2_X2 U370 ( .A(n587), .B(n429), .ZN(n613) );
  XNOR2_X2 U371 ( .A(n397), .B(n522), .ZN(n473) );
  NOR2_X1 U372 ( .A1(G953), .A2(G237), .ZN(n505) );
  OR2_X1 U373 ( .A1(n565), .A2(n426), .ZN(n425) );
  AND2_X1 U374 ( .A1(n580), .A2(n646), .ZN(n582) );
  OR2_X1 U375 ( .A1(n618), .A2(n347), .ZN(n372) );
  AND2_X1 U376 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U377 ( .A(KEYINPUT45), .ZN(n423) );
  NOR2_X1 U378 ( .A1(n700), .A2(n712), .ZN(n398) );
  XNOR2_X1 U379 ( .A(n590), .B(n437), .ZN(n436) );
  NOR2_X1 U380 ( .A1(n612), .A2(n446), .ZN(n405) );
  NOR2_X1 U381 ( .A1(n541), .A2(n671), .ZN(n566) );
  AND2_X1 U382 ( .A1(n387), .A2(KEYINPUT84), .ZN(n386) );
  NOR2_X1 U383 ( .A1(n389), .A2(n445), .ZN(n385) );
  XNOR2_X1 U384 ( .A(n504), .B(n503), .ZN(n551) );
  NAND2_X1 U385 ( .A1(n421), .A2(n420), .ZN(n476) );
  XNOR2_X1 U386 ( .A(n471), .B(n470), .ZN(n397) );
  XNOR2_X1 U387 ( .A(n403), .B(n459), .ZN(n471) );
  XNOR2_X1 U388 ( .A(n349), .B(n472), .ZN(n522) );
  XNOR2_X1 U389 ( .A(n379), .B(G119), .ZN(n403) );
  XNOR2_X1 U390 ( .A(n469), .B(KEYINPUT16), .ZN(n470) );
  XNOR2_X1 U391 ( .A(G104), .B(KEYINPUT75), .ZN(n409) );
  INV_X1 U392 ( .A(KEYINPUT105), .ZN(n404) );
  XNOR2_X1 U393 ( .A(G116), .B(G113), .ZN(n379) );
  NOR2_X1 U394 ( .A1(n441), .A2(n440), .ZN(n439) );
  BUF_X1 U395 ( .A(n441), .Z(n345) );
  NAND2_X1 U396 ( .A1(n438), .A2(n362), .ZN(n441) );
  BUF_X1 U397 ( .A(n553), .Z(n346) );
  XNOR2_X1 U398 ( .A(n468), .B(n467), .ZN(n553) );
  XNOR2_X2 U399 ( .A(n430), .B(G469), .ZN(n587) );
  OR2_X2 U400 ( .A1(n378), .A2(G902), .ZN(n430) );
  XNOR2_X1 U401 ( .A(n508), .B(n456), .ZN(n411) );
  NAND2_X1 U402 ( .A1(n350), .A2(n479), .ZN(n390) );
  XNOR2_X1 U403 ( .A(KEYINPUT72), .B(G472), .ZN(n467) );
  NOR2_X1 U404 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X1 U405 ( .A1(n610), .A2(n434), .ZN(n376) );
  INV_X1 U406 ( .A(KEYINPUT46), .ZN(n437) );
  XNOR2_X1 U407 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n453) );
  XNOR2_X1 U408 ( .A(n512), .B(n474), .ZN(n454) );
  INV_X1 U409 ( .A(G143), .ZN(n464) );
  XNOR2_X1 U410 ( .A(n577), .B(KEYINPUT74), .ZN(n578) );
  XOR2_X1 U411 ( .A(G101), .B(KEYINPUT5), .Z(n461) );
  XNOR2_X1 U412 ( .A(n497), .B(n399), .ZN(n499) );
  INV_X1 U413 ( .A(KEYINPUT95), .ZN(n399) );
  XNOR2_X1 U414 ( .A(G107), .B(G116), .ZN(n495) );
  XNOR2_X1 U415 ( .A(n494), .B(n493), .ZN(n529) );
  XNOR2_X1 U416 ( .A(G110), .B(G101), .ZN(n472) );
  NOR2_X1 U417 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U418 ( .A(n518), .B(KEYINPUT100), .ZN(n358) );
  NOR2_X1 U419 ( .A1(G902), .A2(n708), .ZN(n504) );
  INV_X1 U420 ( .A(G478), .ZN(n502) );
  INV_X1 U421 ( .A(KEYINPUT6), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n535), .B(n534), .ZN(n664) );
  XNOR2_X1 U423 ( .A(n723), .B(n442), .ZN(n711) );
  XNOR2_X1 U424 ( .A(n444), .B(n443), .ZN(n442) );
  NAND2_X1 U425 ( .A1(n529), .A2(G221), .ZN(n443) );
  XNOR2_X1 U426 ( .A(n531), .B(n530), .ZN(n444) );
  XNOR2_X1 U427 ( .A(n514), .B(n513), .ZN(n703) );
  INV_X1 U428 ( .A(G469), .ZN(n414) );
  XNOR2_X1 U429 ( .A(n523), .B(n524), .ZN(n378) );
  XNOR2_X1 U430 ( .A(n522), .B(n521), .ZN(n524) );
  XNOR2_X1 U431 ( .A(n525), .B(n455), .ZN(n521) );
  AND2_X1 U432 ( .A1(G227), .A2(n727), .ZN(n455) );
  OR2_X1 U433 ( .A1(G902), .A2(G237), .ZN(n481) );
  INV_X1 U434 ( .A(n633), .ZN(n426) );
  XOR2_X1 U435 ( .A(KEYINPUT9), .B(G122), .Z(n496) );
  XNOR2_X1 U436 ( .A(KEYINPUT86), .B(G107), .ZN(n410) );
  AND2_X1 U437 ( .A1(n435), .A2(n611), .ZN(n432) );
  XOR2_X1 U438 ( .A(KEYINPUT99), .B(n517), .Z(n656) );
  INV_X1 U439 ( .A(KEYINPUT1), .ZN(n429) );
  XNOR2_X1 U440 ( .A(G128), .B(G110), .ZN(n527) );
  XOR2_X1 U441 ( .A(G137), .B(G119), .Z(n528) );
  XOR2_X1 U442 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n530) );
  XOR2_X1 U443 ( .A(G122), .B(G113), .Z(n510) );
  XNOR2_X1 U444 ( .A(G140), .B(G143), .ZN(n509) );
  XNOR2_X1 U445 ( .A(n360), .B(n359), .ZN(n511) );
  XNOR2_X1 U446 ( .A(n507), .B(n506), .ZN(n360) );
  XOR2_X1 U447 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n507) );
  XOR2_X1 U448 ( .A(KEYINPUT10), .B(n512), .Z(n526) );
  XOR2_X1 U449 ( .A(G140), .B(KEYINPUT69), .Z(n525) );
  XNOR2_X1 U450 ( .A(n454), .B(n452), .ZN(n477) );
  XNOR2_X1 U451 ( .A(n475), .B(n453), .ZN(n452) );
  NAND2_X1 U452 ( .A1(n396), .A2(n395), .ZN(n431) );
  INV_X1 U453 ( .A(n655), .ZN(n395) );
  XOR2_X1 U454 ( .A(KEYINPUT34), .B(KEYINPUT76), .Z(n548) );
  XNOR2_X1 U455 ( .A(n603), .B(KEYINPUT19), .ZN(n597) );
  XNOR2_X1 U456 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n415) );
  XNOR2_X1 U457 ( .A(n523), .B(n465), .ZN(n466) );
  NOR2_X1 U458 ( .A1(n441), .A2(n428), .ZN(n427) );
  INV_X1 U459 ( .A(G472), .ZN(n428) );
  XNOR2_X1 U460 ( .A(n501), .B(n500), .ZN(n708) );
  AND2_X1 U461 ( .A1(n375), .A2(n374), .ZN(n373) );
  AND2_X1 U462 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U463 ( .A1(n364), .A2(n363), .ZN(n556) );
  XNOR2_X1 U464 ( .A(KEYINPUT109), .B(n595), .ZN(n735) );
  NAND2_X1 U465 ( .A1(n555), .A2(n554), .ZN(n381) );
  XNOR2_X1 U466 ( .A(n393), .B(n451), .ZN(n450) );
  XNOR2_X1 U467 ( .A(n408), .B(n704), .ZN(n705) );
  NOR2_X1 U468 ( .A1(n345), .A2(n414), .ZN(n413) );
  INV_X2 U469 ( .A(G953), .ZN(n727) );
  OR2_X1 U470 ( .A1(n619), .A2(KEYINPUT107), .ZN(n347) );
  XOR2_X1 U471 ( .A(KEYINPUT78), .B(KEYINPUT88), .Z(n348) );
  XOR2_X1 U472 ( .A(n410), .B(n409), .Z(n349) );
  XOR2_X1 U473 ( .A(n480), .B(n348), .Z(n350) );
  AND2_X1 U474 ( .A1(n381), .A2(n380), .ZN(n351) );
  AND2_X1 U475 ( .A1(n436), .A2(n432), .ZN(n352) );
  NAND2_X1 U476 ( .A1(n384), .A2(n382), .ZN(n603) );
  AND2_X1 U477 ( .A1(n388), .A2(n383), .ZN(n353) );
  OR2_X1 U478 ( .A1(n350), .A2(n479), .ZN(n354) );
  INV_X1 U479 ( .A(n583), .ZN(n446) );
  INV_X1 U480 ( .A(n344), .ZN(n363) );
  INV_X1 U481 ( .A(KEYINPUT84), .ZN(n445) );
  INV_X1 U482 ( .A(n611), .ZN(n434) );
  XNOR2_X1 U483 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n355) );
  XOR2_X1 U484 ( .A(n699), .B(n698), .Z(n356) );
  XNOR2_X1 U485 ( .A(G902), .B(KEYINPUT15), .ZN(n628) );
  XNOR2_X1 U486 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n357) );
  NOR2_X1 U487 ( .A1(G952), .A2(n727), .ZN(n712) );
  INV_X1 U488 ( .A(n508), .ZN(n359) );
  INV_X1 U489 ( .A(n537), .ZN(n550) );
  XNOR2_X1 U490 ( .A(n516), .B(n515), .ZN(n537) );
  XNOR2_X2 U491 ( .A(n473), .B(n478), .ZN(n697) );
  NOR2_X1 U492 ( .A1(n591), .A2(n592), .ZN(n593) );
  NAND2_X1 U493 ( .A1(n575), .A2(n576), .ZN(n591) );
  NOR2_X1 U494 ( .A1(G902), .A2(n711), .ZN(n535) );
  NAND2_X1 U495 ( .A1(n622), .A2(n653), .ZN(n394) );
  INV_X1 U496 ( .A(n610), .ZN(n435) );
  NAND2_X1 U497 ( .A1(n361), .A2(n351), .ZN(n562) );
  XNOR2_X1 U498 ( .A(n561), .B(KEYINPUT66), .ZN(n361) );
  NAND2_X1 U499 ( .A1(n362), .A2(n627), .ZN(n692) );
  AND2_X1 U500 ( .A1(n362), .A2(G475), .ZN(n407) );
  AND2_X1 U501 ( .A1(n362), .A2(G217), .ZN(n392) );
  NAND2_X2 U502 ( .A1(n621), .A2(n620), .ZN(n362) );
  INV_X1 U503 ( .A(n365), .ZN(n364) );
  NAND2_X1 U504 ( .A1(n602), .A2(n365), .ZN(n400) );
  NAND2_X1 U505 ( .A1(n419), .A2(n365), .ZN(n418) );
  NOR2_X1 U506 ( .A1(n552), .A2(n365), .ZN(n536) );
  XNOR2_X2 U507 ( .A(n668), .B(n366), .ZN(n365) );
  NAND2_X1 U508 ( .A1(n373), .A2(n372), .ZN(n734) );
  NAND2_X1 U509 ( .A1(n369), .A2(n367), .ZN(n433) );
  NAND2_X1 U510 ( .A1(n368), .A2(n434), .ZN(n367) );
  INV_X1 U511 ( .A(n436), .ZN(n368) );
  NAND2_X1 U512 ( .A1(n372), .A2(n376), .ZN(n370) );
  INV_X1 U513 ( .A(n373), .ZN(n371) );
  NAND2_X1 U514 ( .A1(n619), .A2(KEYINPUT107), .ZN(n374) );
  NAND2_X1 U515 ( .A1(n618), .A2(KEYINPUT107), .ZN(n375) );
  NAND2_X1 U516 ( .A1(n377), .A2(n547), .ZN(n549) );
  NAND2_X1 U517 ( .A1(n377), .A2(n663), .ZN(n685) );
  NAND2_X1 U518 ( .A1(n682), .A2(n377), .ZN(n654) );
  XNOR2_X2 U519 ( .A(n418), .B(KEYINPUT33), .ZN(n377) );
  XNOR2_X1 U520 ( .A(n378), .B(n357), .ZN(n412) );
  INV_X1 U521 ( .A(n737), .ZN(n380) );
  XNOR2_X1 U522 ( .A(n381), .B(G110), .ZN(G12) );
  NAND2_X1 U523 ( .A1(n389), .A2(n388), .ZN(n592) );
  NAND2_X1 U524 ( .A1(n389), .A2(n353), .ZN(n382) );
  NOR2_X1 U525 ( .A1(n446), .A2(KEYINPUT84), .ZN(n383) );
  NAND2_X1 U526 ( .A1(n388), .A2(n583), .ZN(n387) );
  OR2_X2 U527 ( .A1(n697), .A2(n354), .ZN(n388) );
  NAND2_X1 U528 ( .A1(n697), .A2(n350), .ZN(n391) );
  NAND2_X1 U529 ( .A1(n392), .A2(n438), .ZN(n393) );
  INV_X1 U530 ( .A(n345), .ZN(n710) );
  XNOR2_X1 U531 ( .A(n492), .B(n457), .ZN(n501) );
  NOR2_X2 U532 ( .A1(n613), .A2(n671), .ZN(n546) );
  XNOR2_X1 U533 ( .A(n400), .B(KEYINPUT104), .ZN(n612) );
  XNOR2_X2 U534 ( .A(n394), .B(KEYINPUT81), .ZN(n725) );
  INV_X1 U535 ( .A(n591), .ZN(n396) );
  XNOR2_X1 U536 ( .A(n439), .B(n356), .ZN(n700) );
  XNOR2_X1 U537 ( .A(n398), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U538 ( .A1(n401), .A2(KEYINPUT44), .ZN(n563) );
  NAND2_X1 U539 ( .A1(n351), .A2(n560), .ZN(n401) );
  NAND2_X1 U540 ( .A1(n450), .A2(n630), .ZN(n449) );
  XNOR2_X2 U541 ( .A(n402), .B(KEYINPUT41), .ZN(n682) );
  NAND2_X1 U542 ( .A1(n660), .A2(n656), .ZN(n402) );
  XNOR2_X1 U543 ( .A(n405), .B(n404), .ZN(n614) );
  INV_X2 U544 ( .A(n553), .ZN(n668) );
  NAND2_X1 U545 ( .A1(n597), .A2(n488), .ZN(n406) );
  INV_X1 U546 ( .A(n473), .ZN(n713) );
  NAND2_X1 U547 ( .A1(n407), .A2(n438), .ZN(n408) );
  XNOR2_X2 U548 ( .A(n492), .B(n411), .ZN(n724) );
  XNOR2_X2 U549 ( .A(n476), .B(G134), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n413), .B(n412), .ZN(n701) );
  XNOR2_X1 U551 ( .A(n416), .B(n415), .ZN(n588) );
  NOR2_X1 U552 ( .A1(n346), .A2(n417), .ZN(n416) );
  INV_X1 U553 ( .A(n601), .ZN(n417) );
  XNOR2_X1 U554 ( .A(n546), .B(KEYINPUT102), .ZN(n419) );
  NAND2_X1 U555 ( .A1(n463), .A2(n464), .ZN(n420) );
  NAND2_X1 U556 ( .A1(n422), .A2(G143), .ZN(n421) );
  INV_X1 U557 ( .A(n463), .ZN(n422) );
  NAND2_X1 U558 ( .A1(n715), .A2(n626), .ZN(n627) );
  XNOR2_X2 U559 ( .A(n424), .B(n423), .ZN(n715) );
  NOR2_X2 U560 ( .A1(n564), .A2(n425), .ZN(n424) );
  XNOR2_X1 U561 ( .A(n427), .B(n629), .ZN(n631) );
  AND2_X2 U562 ( .A1(n627), .A2(n479), .ZN(n438) );
  XNOR2_X2 U563 ( .A(n431), .B(KEYINPUT39), .ZN(n580) );
  NOR2_X2 U564 ( .A1(n433), .A2(n352), .ZN(n622) );
  INV_X1 U565 ( .A(G210), .ZN(n440) );
  INV_X1 U566 ( .A(n592), .ZN(n619) );
  NOR2_X1 U567 ( .A1(n736), .A2(KEYINPUT44), .ZN(n561) );
  XNOR2_X2 U568 ( .A(n447), .B(n355), .ZN(n736) );
  NAND2_X1 U569 ( .A1(n448), .A2(n594), .ZN(n447) );
  XNOR2_X1 U570 ( .A(n549), .B(n548), .ZN(n448) );
  XNOR2_X1 U571 ( .A(n449), .B(KEYINPUT125), .ZN(G66) );
  INV_X1 U572 ( .A(n711), .ZN(n451) );
  INV_X1 U573 ( .A(n542), .ZN(n547) );
  XOR2_X1 U574 ( .A(G137), .B(KEYINPUT4), .Z(n456) );
  AND2_X1 U575 ( .A1(G217), .A2(n529), .ZN(n457) );
  XOR2_X1 U576 ( .A(n510), .B(n509), .Z(n458) );
  XNOR2_X1 U577 ( .A(n511), .B(n458), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n615), .B(KEYINPUT106), .ZN(n616) );
  XNOR2_X1 U579 ( .A(n502), .B(KEYINPUT97), .ZN(n503) );
  XNOR2_X1 U580 ( .A(n604), .B(KEYINPUT113), .ZN(n605) );
  INV_X1 U581 ( .A(n712), .ZN(n630) );
  XNOR2_X1 U582 ( .A(n606), .B(n605), .ZN(n608) );
  NAND2_X1 U583 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U584 ( .A(n632), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U585 ( .A(KEYINPUT71), .B(KEYINPUT3), .ZN(n459) );
  NAND2_X1 U586 ( .A1(n505), .A2(G210), .ZN(n460) );
  XNOR2_X1 U587 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U588 ( .A(n471), .B(n462), .ZN(n465) );
  XNOR2_X2 U589 ( .A(G128), .B(KEYINPUT77), .ZN(n463) );
  XOR2_X1 U590 ( .A(G131), .B(KEYINPUT68), .Z(n508) );
  XNOR2_X1 U591 ( .A(n466), .B(KEYINPUT62), .ZN(n629) );
  NOR2_X1 U592 ( .A1(G902), .A2(n466), .ZN(n468) );
  XOR2_X1 U593 ( .A(KEYINPUT73), .B(G122), .Z(n469) );
  XOR2_X2 U594 ( .A(G125), .B(G146), .Z(n512) );
  XNOR2_X1 U595 ( .A(KEYINPUT18), .B(KEYINPUT87), .ZN(n474) );
  NAND2_X1 U596 ( .A1(G224), .A2(n727), .ZN(n475) );
  XOR2_X1 U597 ( .A(n476), .B(n477), .Z(n478) );
  INV_X1 U598 ( .A(n628), .ZN(n479) );
  NAND2_X1 U599 ( .A1(G210), .A2(n481), .ZN(n480) );
  NAND2_X1 U600 ( .A1(G214), .A2(n481), .ZN(n583) );
  NOR2_X1 U601 ( .A1(G898), .A2(n727), .ZN(n482) );
  XNOR2_X1 U602 ( .A(KEYINPUT90), .B(n482), .ZN(n714) );
  NAND2_X1 U603 ( .A1(G237), .A2(G234), .ZN(n483) );
  XNOR2_X1 U604 ( .A(n483), .B(KEYINPUT14), .ZN(n485) );
  NAND2_X1 U605 ( .A1(n485), .A2(G902), .ZN(n484) );
  XNOR2_X1 U606 ( .A(n484), .B(KEYINPUT91), .ZN(n567) );
  NAND2_X1 U607 ( .A1(n714), .A2(n567), .ZN(n487) );
  NAND2_X1 U608 ( .A1(G952), .A2(n485), .ZN(n689) );
  NOR2_X1 U609 ( .A1(n689), .A2(G953), .ZN(n486) );
  XNOR2_X1 U610 ( .A(n486), .B(KEYINPUT89), .ZN(n570) );
  NAND2_X1 U611 ( .A1(n487), .A2(n570), .ZN(n488) );
  XOR2_X1 U612 ( .A(KEYINPUT21), .B(KEYINPUT92), .Z(n491) );
  NAND2_X1 U613 ( .A1(G234), .A2(n628), .ZN(n489) );
  XNOR2_X1 U614 ( .A(KEYINPUT20), .B(n489), .ZN(n532) );
  NAND2_X1 U615 ( .A1(n532), .A2(G221), .ZN(n490) );
  XNOR2_X1 U616 ( .A(n491), .B(n490), .ZN(n665) );
  XOR2_X1 U617 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n494) );
  NAND2_X1 U618 ( .A1(G234), .A2(n727), .ZN(n493) );
  XNOR2_X1 U619 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U620 ( .A(KEYINPUT96), .B(KEYINPUT7), .ZN(n498) );
  XNOR2_X1 U621 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U622 ( .A1(n505), .A2(G214), .ZN(n506) );
  XNOR2_X1 U623 ( .A(n526), .B(G104), .ZN(n513) );
  NOR2_X1 U624 ( .A1(G902), .A2(n703), .ZN(n516) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(G475), .ZN(n515) );
  AND2_X1 U626 ( .A1(n551), .A2(n550), .ZN(n517) );
  NAND2_X1 U627 ( .A1(n665), .A2(n656), .ZN(n518) );
  XNOR2_X1 U628 ( .A(KEYINPUT22), .B(KEYINPUT64), .ZN(n519) );
  XNOR2_X1 U629 ( .A(n520), .B(n519), .ZN(n558) );
  INV_X1 U630 ( .A(n613), .ZN(n607) );
  INV_X1 U631 ( .A(n607), .ZN(n672) );
  NAND2_X1 U632 ( .A1(n558), .A2(n672), .ZN(n552) );
  XNOR2_X1 U633 ( .A(n526), .B(n525), .ZN(n723) );
  XNOR2_X1 U634 ( .A(n528), .B(n527), .ZN(n531) );
  NAND2_X1 U635 ( .A1(n532), .A2(G217), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n533), .B(KEYINPUT25), .ZN(n534) );
  NAND2_X1 U637 ( .A1(n536), .A2(n344), .ZN(n633) );
  NOR2_X1 U638 ( .A1(n537), .A2(n551), .ZN(n648) );
  NAND2_X1 U639 ( .A1(n537), .A2(n551), .ZN(n538) );
  XOR2_X2 U640 ( .A(KEYINPUT98), .B(n538), .Z(n646) );
  NOR2_X1 U641 ( .A1(n648), .A2(n646), .ZN(n658) );
  NAND2_X1 U642 ( .A1(n665), .A2(n344), .ZN(n671) );
  NAND2_X1 U643 ( .A1(n546), .A2(n668), .ZN(n678) );
  NOR2_X1 U644 ( .A1(n542), .A2(n678), .ZN(n540) );
  XNOR2_X1 U645 ( .A(KEYINPUT31), .B(KEYINPUT93), .ZN(n539) );
  XNOR2_X1 U646 ( .A(n540), .B(n539), .ZN(n649) );
  INV_X1 U647 ( .A(n587), .ZN(n541) );
  NAND2_X1 U648 ( .A1(n566), .A2(n547), .ZN(n543) );
  NOR2_X1 U649 ( .A1(n668), .A2(n543), .ZN(n638) );
  NOR2_X1 U650 ( .A1(n649), .A2(n638), .ZN(n544) );
  XNOR2_X1 U651 ( .A(n544), .B(KEYINPUT94), .ZN(n545) );
  NOR2_X1 U652 ( .A1(n658), .A2(n545), .ZN(n565) );
  NOR2_X1 U653 ( .A1(n551), .A2(n550), .ZN(n594) );
  INV_X1 U654 ( .A(n736), .ZN(n560) );
  XNOR2_X1 U655 ( .A(n552), .B(KEYINPUT101), .ZN(n555) );
  AND2_X1 U656 ( .A1(n346), .A2(n363), .ZN(n554) );
  NOR2_X1 U657 ( .A1(n556), .A2(n672), .ZN(n557) );
  XNOR2_X1 U658 ( .A(n559), .B(KEYINPUT32), .ZN(n737) );
  NAND2_X1 U659 ( .A1(n562), .A2(n563), .ZN(n564) );
  XNOR2_X1 U660 ( .A(KEYINPUT108), .B(n566), .ZN(n576) );
  NAND2_X1 U661 ( .A1(G953), .A2(n567), .ZN(n568) );
  NOR2_X1 U662 ( .A1(G900), .A2(n568), .ZN(n569) );
  XNOR2_X1 U663 ( .A(n569), .B(KEYINPUT103), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n571), .A2(n570), .ZN(n585) );
  INV_X1 U665 ( .A(n585), .ZN(n574) );
  NAND2_X1 U666 ( .A1(n583), .A2(n668), .ZN(n572) );
  XNOR2_X1 U667 ( .A(KEYINPUT30), .B(n572), .ZN(n573) );
  NOR2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n575) );
  INV_X1 U669 ( .A(KEYINPUT38), .ZN(n577) );
  XNOR2_X1 U670 ( .A(n592), .B(n578), .ZN(n655) );
  NAND2_X1 U671 ( .A1(n580), .A2(n648), .ZN(n653) );
  XNOR2_X1 U672 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n579) );
  XNOR2_X1 U673 ( .A(n579), .B(KEYINPUT70), .ZN(n611) );
  XNOR2_X1 U674 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n581) );
  NOR2_X1 U675 ( .A1(n446), .A2(n655), .ZN(n584) );
  XNOR2_X1 U676 ( .A(KEYINPUT112), .B(n584), .ZN(n660) );
  NAND2_X1 U677 ( .A1(n665), .A2(n585), .ZN(n586) );
  NOR2_X1 U678 ( .A1(n344), .A2(n586), .ZN(n601) );
  AND2_X1 U679 ( .A1(n587), .A2(n588), .ZN(n596) );
  NAND2_X1 U680 ( .A1(n682), .A2(n596), .ZN(n589) );
  XNOR2_X1 U681 ( .A(KEYINPUT42), .B(n589), .ZN(n739) );
  NAND2_X1 U682 ( .A1(n740), .A2(n739), .ZN(n590) );
  NAND2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U684 ( .A1(KEYINPUT67), .A2(n658), .ZN(n598) );
  AND2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n644) );
  NAND2_X1 U686 ( .A1(n598), .A2(n644), .ZN(n599) );
  XNOR2_X1 U687 ( .A(KEYINPUT47), .B(n599), .ZN(n600) );
  NOR2_X1 U688 ( .A1(n735), .A2(n600), .ZN(n609) );
  AND2_X1 U689 ( .A1(n646), .A2(n601), .ZN(n602) );
  NOR2_X1 U690 ( .A1(n612), .A2(n603), .ZN(n606) );
  INV_X1 U691 ( .A(KEYINPUT36), .ZN(n604) );
  NAND2_X1 U692 ( .A1(n608), .A2(n607), .ZN(n652) );
  NAND2_X1 U693 ( .A1(n609), .A2(n652), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n614), .A2(n672), .ZN(n617) );
  INV_X1 U695 ( .A(KEYINPUT43), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n617), .B(n616), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n715), .A2(n725), .ZN(n621) );
  INV_X1 U698 ( .A(KEYINPUT2), .ZN(n620) );
  INV_X1 U699 ( .A(n622), .ZN(n625) );
  NAND2_X1 U700 ( .A1(KEYINPUT2), .A2(n653), .ZN(n623) );
  XOR2_X1 U701 ( .A(KEYINPUT79), .B(n623), .Z(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U703 ( .A(G101), .B(n633), .ZN(G3) );
  NAND2_X1 U704 ( .A1(n646), .A2(n638), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n634), .B(G104), .ZN(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n636) );
  XNOR2_X1 U707 ( .A(G107), .B(KEYINPUT26), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(n637) );
  XOR2_X1 U709 ( .A(KEYINPUT114), .B(n637), .Z(n640) );
  NAND2_X1 U710 ( .A1(n638), .A2(n648), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(G9) );
  XOR2_X1 U712 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n642) );
  NAND2_X1 U713 ( .A1(n648), .A2(n644), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(G128), .B(n643), .ZN(G30) );
  NAND2_X1 U716 ( .A1(n646), .A2(n644), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(G146), .ZN(G48) );
  NAND2_X1 U718 ( .A1(n646), .A2(n649), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(G113), .ZN(G15) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(G116), .ZN(G18) );
  XOR2_X1 U722 ( .A(G125), .B(KEYINPUT37), .Z(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(G27) );
  XNOR2_X1 U724 ( .A(G134), .B(n653), .ZN(G36) );
  XNOR2_X1 U725 ( .A(n654), .B(KEYINPUT123), .ZN(n691) );
  NAND2_X1 U726 ( .A1(n655), .A2(n446), .ZN(n657) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n662) );
  INV_X1 U728 ( .A(n658), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U731 ( .A1(n665), .A2(n344), .ZN(n667) );
  XNOR2_X1 U732 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n667), .B(n666), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U735 ( .A(KEYINPUT118), .B(n670), .ZN(n676) );
  XOR2_X1 U736 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n674) );
  NAND2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U738 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n677), .B(KEYINPUT120), .ZN(n679) );
  NAND2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U742 ( .A(KEYINPUT51), .B(n680), .Z(n681) );
  NAND2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U744 ( .A(KEYINPUT121), .B(n683), .Z(n684) );
  NAND2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U746 ( .A(n686), .B(KEYINPUT52), .ZN(n687) );
  XOR2_X1 U747 ( .A(KEYINPUT122), .B(n687), .Z(n688) );
  NOR2_X1 U748 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U751 ( .A(KEYINPUT124), .B(n694), .ZN(n695) );
  NOR2_X1 U752 ( .A1(n695), .A2(G953), .ZN(n696) );
  XNOR2_X1 U753 ( .A(n696), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U754 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n699) );
  XNOR2_X1 U755 ( .A(n697), .B(KEYINPUT85), .ZN(n698) );
  NOR2_X1 U756 ( .A1(n712), .A2(n701), .ZN(G54) );
  XOR2_X1 U757 ( .A(KEYINPUT59), .B(KEYINPUT65), .Z(n702) );
  XNOR2_X1 U758 ( .A(n703), .B(n702), .ZN(n704) );
  AND2_X1 U759 ( .A1(n630), .A2(n705), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n706), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U761 ( .A1(G478), .A2(n710), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U763 ( .A1(n712), .A2(n709), .ZN(G63) );
  NOR2_X1 U764 ( .A1(n714), .A2(n713), .ZN(n722) );
  NAND2_X1 U765 ( .A1(n727), .A2(n715), .ZN(n719) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n716) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n716), .ZN(n717) );
  NAND2_X1 U768 ( .A1(n717), .A2(G898), .ZN(n718) );
  NAND2_X1 U769 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n720), .B(KEYINPUT126), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(n729) );
  INV_X1 U773 ( .A(n729), .ZN(n726) );
  XOR2_X1 U774 ( .A(n726), .B(n725), .Z(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(n727), .ZN(n733) );
  XOR2_X1 U776 ( .A(G227), .B(n729), .Z(n730) );
  NAND2_X1 U777 ( .A1(n730), .A2(G900), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n731), .A2(G953), .ZN(n732) );
  NAND2_X1 U779 ( .A1(n733), .A2(n732), .ZN(G72) );
  XOR2_X1 U780 ( .A(n734), .B(G140), .Z(G42) );
  XOR2_X1 U781 ( .A(G143), .B(n735), .Z(G45) );
  XOR2_X1 U782 ( .A(n736), .B(G122), .Z(G24) );
  XNOR2_X1 U783 ( .A(G119), .B(KEYINPUT127), .ZN(n738) );
  XNOR2_X1 U784 ( .A(n738), .B(n737), .ZN(G21) );
  XNOR2_X1 U785 ( .A(n739), .B(G137), .ZN(G39) );
  XNOR2_X1 U786 ( .A(n740), .B(G131), .ZN(G33) );
endmodule

