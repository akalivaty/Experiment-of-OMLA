//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1388, new_n1389,
    new_n1390, new_n1391;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n213), .A2(G50), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n208), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(new_n205), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n216), .B(new_n224), .C1(KEYINPUT1), .C2(new_n222), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G97), .B(G107), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n242));
  INV_X1    g0042(.A(G226), .ZN(new_n243));
  INV_X1    g0043(.A(G1698), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G232), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G1698), .ZN(new_n249));
  NAND4_X1  g0049(.A1(new_n242), .A2(new_n245), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G97), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT13), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(new_n254), .A3(G274), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n254), .A2(G238), .A3(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n256), .A2(new_n257), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n254), .B1(new_n250), .B2(new_n251), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n264), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT13), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(G179), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT71), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n266), .A2(new_n272), .A3(new_n269), .ZN(new_n273));
  OAI211_X1 g0073(.A(KEYINPUT71), .B(KEYINPUT13), .C1(new_n267), .C2(new_n268), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G169), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT14), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n273), .A2(KEYINPUT14), .A3(G169), .A4(new_n274), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n271), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT67), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n282), .A2(KEYINPUT66), .A3(new_n209), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT66), .B1(new_n282), .B2(new_n209), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n209), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT66), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n282), .A2(KEYINPUT66), .A3(new_n209), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(KEYINPUT67), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G68), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G77), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n210), .A2(G33), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n291), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n283), .A2(new_n284), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n210), .A2(G1), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n293), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT12), .B1(new_n300), .B2(G68), .ZN(new_n305));
  OR3_X1    g0105(.A1(new_n300), .A2(KEYINPUT12), .A3(G68), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n302), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT11), .B1(new_n291), .B2(new_n297), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n280), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G244), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n255), .A2(new_n260), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n261), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT3), .B(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(G232), .A2(G1698), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n244), .A2(G238), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n255), .C1(G107), .C2(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G200), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  INV_X1    g0125(.A(new_n303), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n302), .A2(G77), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT15), .B(G87), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n296), .B1(new_n210), .B2(new_n295), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT69), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n330), .B(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n329), .B1(new_n332), .B2(new_n292), .ZN(new_n333));
  INV_X1    g0133(.A(new_n299), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n327), .B1(G77), .B2(new_n300), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n325), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n322), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n322), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n339), .A2(KEYINPUT70), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT70), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n335), .A2(new_n346), .A3(new_n338), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n336), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n273), .A2(G200), .A3(new_n274), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n266), .A2(G190), .A3(new_n269), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n310), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n312), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n255), .A2(new_n260), .A3(new_n243), .ZN(new_n354));
  NOR2_X1   g0154(.A1(G222), .A2(G1698), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n244), .A2(G223), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n317), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n242), .A2(new_n247), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n254), .B1(new_n358), .B2(new_n295), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n315), .B(new_n354), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n344), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G169), .B2(new_n360), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n285), .A2(new_n290), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n363), .A2(G50), .A3(new_n300), .A4(new_n326), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  INV_X1    g0166(.A(new_n292), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .C1(new_n296), .C2(new_n330), .ZN(new_n368));
  INV_X1    g0168(.A(G50), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(new_n291), .B1(new_n369), .B2(new_n301), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n360), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(G190), .B2(new_n360), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n371), .A2(KEYINPUT9), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n371), .A2(KEYINPUT9), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(KEYINPUT10), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(KEYINPUT10), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n373), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n330), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n301), .B1(new_n383), .B2(new_n326), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n285), .A2(new_n290), .A3(new_n300), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n383), .ZN(new_n386));
  INV_X1    g0186(.A(G58), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n293), .ZN(new_n388));
  OAI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n201), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n292), .A2(G159), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n358), .A2(new_n210), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n246), .A2(G33), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(KEYINPUT72), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n242), .A2(new_n247), .A3(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n393), .A2(new_n394), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n392), .B1(new_n400), .B2(new_n293), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n334), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n395), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n393), .A2(new_n394), .B1(new_n358), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT16), .B(new_n392), .C1(new_n405), .C2(new_n293), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n386), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n243), .A2(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n242), .A2(new_n408), .A3(new_n247), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n255), .ZN(new_n413));
  INV_X1    g0213(.A(new_n344), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n254), .A2(G232), .A3(new_n263), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n261), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n254), .B1(new_n410), .B2(new_n411), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n261), .A2(new_n415), .ZN(new_n419));
  OAI21_X1  g0219(.A(G169), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n417), .A2(KEYINPUT73), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT73), .B1(new_n417), .B2(new_n420), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT18), .B1(new_n407), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n413), .A2(new_n416), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n374), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n425), .B2(G190), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n397), .A2(new_n399), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n394), .B1(new_n317), .B2(G20), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n391), .B1(new_n430), .B2(G68), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n406), .B(new_n299), .C1(new_n431), .C2(KEYINPUT16), .ZN(new_n432));
  INV_X1    g0232(.A(new_n386), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n427), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n407), .A2(KEYINPUT17), .A3(new_n427), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n433), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT73), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n337), .B1(new_n413), .B2(new_n416), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n418), .A2(new_n419), .A3(new_n344), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n417), .A2(KEYINPUT73), .A3(new_n420), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n438), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n424), .A2(new_n436), .A3(new_n437), .A4(new_n446), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n447), .A2(KEYINPUT74), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(KEYINPUT74), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n353), .A2(new_n382), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n262), .B2(G33), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n300), .B(new_n452), .C1(new_n283), .C2(new_n284), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n301), .A2(new_n451), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n282), .A2(new_n209), .B1(G20), .B2(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n210), .C1(G33), .C2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT20), .B1(new_n455), .B2(new_n458), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n453), .B(new_n454), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT79), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n455), .A2(new_n458), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT20), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT79), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n453), .A4(new_n454), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n242), .A2(new_n247), .A3(G264), .A4(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT77), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT77), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n317), .A2(new_n473), .A3(G264), .A4(G1698), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT78), .B(G303), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n358), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n317), .A2(G257), .A3(new_n244), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n472), .A2(new_n474), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n255), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT5), .B(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n259), .A2(G1), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G270), .A3(new_n254), .ZN(new_n483));
  INV_X1    g0283(.A(G274), .ZN(new_n484));
  INV_X1    g0284(.A(new_n209), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n253), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n481), .A3(new_n480), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n337), .B1(new_n479), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n470), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT81), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(new_n495), .A3(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n470), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n479), .A2(new_n489), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G200), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(KEYINPUT82), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n488), .B1(new_n255), .B2(new_n478), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n374), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n504), .B2(new_n470), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(G190), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n490), .A2(KEYINPUT21), .B1(G179), .B2(new_n503), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT80), .B1(new_n508), .B2(new_n498), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n503), .A2(new_n492), .A3(new_n337), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n499), .A2(new_n341), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n510), .B(new_n470), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n497), .A2(new_n507), .A3(new_n509), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n242), .A2(new_n247), .A3(G244), .A4(new_n244), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT75), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n317), .A2(G250), .A3(G1698), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n456), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n517), .B1(new_n515), .B2(new_n516), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n255), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n482), .A2(G257), .A3(new_n254), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n523), .A2(new_n487), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n524), .A3(new_n344), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n300), .A2(G97), .ZN(new_n526));
  INV_X1    g0326(.A(G107), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n527), .A2(KEYINPUT6), .A3(G97), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  AND2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n400), .B2(new_n527), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n526), .B1(new_n536), .B2(new_n299), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n262), .A2(G33), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n363), .A2(G97), .A3(new_n300), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n522), .A2(new_n524), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n537), .A2(new_n539), .B1(new_n540), .B2(new_n337), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n527), .B1(new_n428), .B2(new_n429), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n528), .B1(new_n543), .B2(new_n530), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n544), .A2(new_n210), .B1(new_n295), .B2(new_n367), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n299), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n526), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n539), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n374), .B1(new_n522), .B2(new_n524), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n522), .A2(new_n524), .A3(G190), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n525), .A2(new_n541), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT23), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n527), .A3(G20), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT84), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT84), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n553), .A2(new_n555), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n242), .A2(new_n247), .A3(new_n210), .A4(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n317), .A2(new_n564), .A3(new_n210), .A4(G87), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT83), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n561), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n567), .B1(new_n561), .B2(new_n566), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT24), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n561), .A2(new_n566), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT83), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n574), .B2(new_n568), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n299), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n285), .A2(new_n290), .A3(new_n300), .A4(new_n538), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n527), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n301), .A2(new_n527), .ZN(new_n579));
  XNOR2_X1  g0379(.A(new_n579), .B(KEYINPUT25), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n482), .A2(G264), .A3(new_n254), .ZN(new_n582));
  MUX2_X1   g0382(.A(G250), .B(G257), .S(G1698), .Z(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n317), .B1(G33), .B2(G294), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n487), .C1(new_n584), .C2(new_n254), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(G190), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n374), .B2(new_n585), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n576), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n585), .A2(G179), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n337), .B2(new_n585), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT24), .B1(new_n569), .B2(new_n570), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n574), .A2(new_n572), .A3(new_n568), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n334), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n581), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G87), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n577), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g0398(.A1(KEYINPUT76), .A2(G87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(KEYINPUT76), .A2(G87), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n532), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n210), .B1(new_n251), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n317), .A2(new_n210), .A3(G68), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n602), .B1(new_n296), .B2(new_n457), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n299), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n328), .A2(new_n301), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G250), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n262), .B2(G45), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n486), .A2(new_n481), .B1(new_n254), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(G238), .A2(G1698), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n313), .B2(G1698), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(new_n317), .B1(G33), .B2(G116), .ZN(new_n616));
  OAI211_X1 g0416(.A(G190), .B(new_n613), .C1(new_n616), .C2(new_n254), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n613), .B1(new_n616), .B2(new_n254), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G200), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n598), .A2(new_n610), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n608), .B(new_n609), .C1(new_n577), .C2(new_n328), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n613), .B(new_n344), .C1(new_n616), .C2(new_n254), .ZN(new_n622));
  OR2_X1    g0422(.A1(G238), .A2(G1698), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n313), .A2(G1698), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n242), .A2(new_n623), .A3(new_n247), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(G33), .A2(G116), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n254), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n254), .A2(G274), .A3(new_n481), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n612), .A2(new_n254), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n337), .B1(new_n627), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n621), .A2(new_n622), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n620), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n552), .A2(new_n589), .A3(new_n596), .A4(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n450), .A2(new_n514), .A3(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n436), .A2(new_n437), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n345), .A2(new_n351), .A3(new_n347), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n312), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n417), .A2(new_n420), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n438), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(new_n439), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n380), .A2(new_n381), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n373), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n540), .A2(new_n337), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n647), .A2(new_n525), .A3(new_n548), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n631), .A2(KEYINPUT85), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT85), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n650), .B(new_n337), .C1(new_n627), .C2(new_n630), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n649), .A2(new_n622), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n619), .A2(new_n617), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n577), .A2(new_n597), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n608), .A2(new_n609), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n652), .A2(new_n621), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n648), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n647), .A2(new_n525), .A3(new_n548), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT26), .B1(new_n633), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n621), .A2(new_n622), .A3(new_n651), .A4(new_n649), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n470), .B1(new_n511), .B2(new_n512), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n497), .A2(new_n664), .A3(new_n596), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n594), .A2(new_n595), .A3(new_n587), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n540), .A2(G200), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(new_n539), .A3(new_n537), .A4(new_n551), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n660), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n620), .A2(new_n662), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n663), .B1(new_n665), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n646), .B1(new_n450), .B2(new_n672), .ZN(G369));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n495), .B1(new_n491), .B2(new_n492), .ZN(new_n675));
  AOI211_X1 g0475(.A(KEYINPUT81), .B(KEYINPUT21), .C1(new_n470), .C2(new_n490), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n509), .B(new_n513), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n507), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n262), .A2(new_n210), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n679), .B1(new_n498), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n664), .B1(new_n675), .B2(new_n676), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n498), .A2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n674), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n685), .B1(new_n594), .B2(new_n595), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n576), .A2(new_n581), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n692), .A2(new_n589), .B1(new_n693), .B2(new_n591), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n591), .B(new_n686), .C1(new_n594), .C2(new_n595), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n509), .A2(new_n513), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n685), .B1(new_n699), .B2(new_n497), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n696), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n206), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n599), .A2(new_n600), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(new_n451), .A3(new_n532), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n706), .A2(new_n708), .B1(new_n215), .B2(new_n705), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n585), .A2(new_n344), .A3(new_n618), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n540), .A3(new_n499), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT86), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n540), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n582), .B1(new_n584), .B2(new_n254), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n618), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n715), .A2(new_n512), .A3(KEYINPUT30), .A4(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n503), .A2(new_n717), .A3(G179), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n540), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n711), .A2(new_n540), .A3(KEYINPUT86), .A4(new_n499), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n714), .A2(new_n718), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n685), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n718), .A2(new_n721), .A3(new_n712), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n686), .A2(new_n725), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n666), .A2(new_n669), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n596), .A3(new_n634), .A4(new_n686), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n730), .B2(new_n514), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n634), .A2(new_n648), .A3(new_n658), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT26), .B1(new_n670), .B2(new_n660), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n662), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n699), .A2(new_n497), .A3(new_n596), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n671), .ZN(new_n737));
  OAI21_X1  g0537(.A(KEYINPUT29), .B1(new_n737), .B2(new_n685), .ZN(new_n738));
  INV_X1    g0538(.A(new_n663), .ZN(new_n739));
  INV_X1    g0539(.A(new_n596), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n688), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n552), .A2(new_n589), .A3(new_n657), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(new_n686), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n732), .A2(new_n738), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n710), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n514), .A2(new_n689), .ZN(new_n749));
  INV_X1    g0549(.A(new_n690), .ZN(new_n750));
  OAI21_X1  g0550(.A(G330), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n687), .A2(new_n674), .A3(new_n690), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n210), .A2(G13), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n262), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n751), .B(new_n752), .C1(new_n704), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n704), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n703), .A2(new_n358), .ZN(new_n758));
  NAND2_X1  g0558(.A1(G355), .A2(KEYINPUT87), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G355), .A2(KEYINPUT87), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(G116), .B2(new_n206), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n236), .A2(new_n259), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n703), .A2(new_n317), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n215), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(new_n259), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n762), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n209), .B1(G20), .B2(new_n337), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n757), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n210), .A2(G190), .A3(G200), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n414), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n358), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(new_n341), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(G329), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n341), .A2(G200), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT90), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(new_n210), .A3(G190), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n786), .A2(new_n210), .A3(new_n324), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G283), .A2(new_n787), .B1(new_n788), .B2(G303), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n344), .A2(new_n210), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(G326), .ZN(new_n792));
  INV_X1    g0592(.A(G294), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n324), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n210), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n783), .B(new_n789), .C1(new_n796), .C2(KEYINPUT91), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(KEYINPUT91), .B2(new_n796), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT88), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n324), .A2(G200), .ZN(new_n800));
  AND3_X1   g0600(.A1(new_n790), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n799), .B1(new_n790), .B2(new_n800), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n790), .A2(new_n324), .A3(G200), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT33), .B(G317), .Z(new_n806));
  OAI22_X1  g0606(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT92), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n798), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n317), .B1(new_n795), .B2(new_n457), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n777), .B2(G77), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n369), .B2(new_n791), .C1(new_n293), .C2(new_n805), .ZN(new_n812));
  INV_X1    g0612(.A(new_n787), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n527), .ZN(new_n814));
  INV_X1    g0614(.A(new_n788), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT32), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT89), .B(G159), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n781), .A2(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n815), .A2(new_n707), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n814), .B(new_n819), .C1(new_n816), .C2(new_n818), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n387), .B2(new_n803), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n809), .B1(new_n812), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n775), .B1(new_n822), .B2(new_n772), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n687), .A2(new_n690), .A3(new_n771), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n756), .A2(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n335), .A2(new_n685), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n348), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n827), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n345), .A2(new_n347), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n672), .B2(new_n685), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n348), .A2(new_n686), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n743), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n757), .B1(new_n836), .B2(new_n732), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n732), .B2(new_n836), .ZN(new_n838));
  INV_X1    g0638(.A(new_n772), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n770), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n757), .B1(G77), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n791), .ZN(new_n842));
  INV_X1    g0642(.A(new_n817), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n842), .A2(G137), .B1(new_n777), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(KEYINPUT93), .B(G143), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n366), .B2(new_n805), .C1(new_n803), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT34), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n317), .B1(new_n781), .B2(new_n848), .C1(new_n387), .C2(new_n795), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n813), .A2(new_n293), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n849), .B(new_n850), .C1(G50), .C2(new_n788), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n813), .A2(new_n597), .ZN(new_n853));
  INV_X1    g0653(.A(new_n795), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n317), .B1(new_n854), .B2(G97), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n855), .B1(new_n779), .B2(new_n781), .C1(new_n778), .C2(new_n451), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n853), .B(new_n856), .C1(G107), .C2(new_n788), .ZN(new_n857));
  INV_X1    g0657(.A(new_n805), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G283), .A2(new_n858), .B1(new_n842), .B2(G303), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(new_n793), .C2(new_n803), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n841), .B1(new_n861), .B2(new_n772), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n828), .A2(new_n830), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n770), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n838), .A2(new_n864), .ZN(G384));
  AOI211_X1 g0665(.A(new_n451), .B(new_n212), .C1(new_n534), .C2(KEYINPUT35), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(KEYINPUT35), .B2(new_n534), .ZN(new_n867));
  XNOR2_X1  g0667(.A(KEYINPUT94), .B(KEYINPUT36), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OR3_X1    g0669(.A1(new_n215), .A2(new_n295), .A3(new_n388), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n369), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n262), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n683), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n438), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n875), .A2(new_n434), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT37), .B1(new_n438), .B2(new_n445), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n392), .B1(new_n405), .B2(new_n293), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n402), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n291), .A3(new_n406), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n433), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n874), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n640), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n883), .A2(new_n884), .A3(new_n434), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n878), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT97), .ZN(new_n888));
  INV_X1    g0688(.A(new_n883), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n447), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n888), .B1(new_n447), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(KEYINPUT38), .B(new_n887), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n277), .A2(new_n278), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n270), .A3(new_n351), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n310), .A2(new_n686), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT96), .ZN(new_n901));
  INV_X1    g0701(.A(new_n899), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n351), .B(new_n902), .C1(new_n279), .C2(new_n310), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT96), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n898), .A2(new_n904), .A3(new_n899), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n514), .A2(new_n635), .A3(new_n685), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n724), .A2(new_n725), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n863), .B(new_n906), .C1(new_n907), .C2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n896), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n637), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n875), .B1(new_n642), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n641), .A2(new_n875), .A3(new_n434), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n876), .A2(new_n877), .B1(new_n918), .B2(KEYINPUT37), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n893), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n895), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n906), .A2(new_n863), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n910), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n635), .A2(new_n685), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n679), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n921), .A2(new_n923), .A3(KEYINPUT40), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n915), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n450), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n927), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n931), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(G330), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n905), .A2(new_n903), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n904), .B1(new_n898), .B2(new_n899), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n345), .A2(new_n347), .A3(new_n686), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT95), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n937), .B1(new_n835), .B2(new_n940), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n941), .A2(new_n896), .B1(new_n643), .B2(new_n683), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT39), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n921), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n280), .A2(new_n311), .A3(new_n686), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n738), .A2(new_n745), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n930), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n646), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n949), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n934), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n262), .B2(new_n753), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n934), .A2(new_n953), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n873), .B1(new_n955), .B2(new_n956), .ZN(G367));
  AOI21_X1  g0757(.A(new_n358), .B1(new_n777), .B2(G50), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n293), .B2(new_n795), .C1(new_n295), .C2(new_n813), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n805), .A2(new_n817), .B1(new_n791), .B2(new_n845), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n788), .A2(G58), .B1(G137), .B2(new_n782), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT104), .Z(new_n963));
  OAI211_X1 g0763(.A(new_n961), .B(new_n963), .C1(new_n366), .C2(new_n803), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G294), .A2(new_n858), .B1(new_n842), .B2(G311), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n787), .A2(G97), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n317), .B1(new_n777), .B2(G283), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G107), .A2(new_n854), .B1(new_n782), .B2(G317), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n803), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT103), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n815), .B2(new_n451), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n970), .A2(new_n475), .B1(new_n972), .B2(KEYINPUT46), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(KEYINPUT46), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n964), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n772), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n656), .A2(new_n686), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n657), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(KEYINPUT98), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(KEYINPUT98), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n979), .A2(new_n662), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n771), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n773), .B1(new_n206), .B2(new_n328), .C1(new_n232), .C2(new_n765), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n977), .A2(new_n757), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n648), .A2(KEYINPUT99), .A3(new_n685), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT99), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n660), .B2(new_n686), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n548), .A2(new_n685), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n552), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n677), .A2(new_n686), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n695), .C1(new_n995), .C2(new_n694), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n692), .A2(new_n589), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n999), .A2(new_n677), .A3(new_n596), .A4(new_n686), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n1000), .A2(KEYINPUT45), .A3(new_n695), .A4(new_n994), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n701), .B2(new_n994), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1000), .A2(new_n695), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n994), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n1007), .A3(new_n1003), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1002), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n698), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1009), .A2(KEYINPUT102), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n695), .B1(new_n999), .B2(new_n740), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n995), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n1000), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n691), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n751), .A2(new_n1000), .A3(new_n1013), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n746), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1010), .B1(new_n1009), .B2(KEYINPUT102), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n747), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n704), .B(KEYINPUT41), .Z(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n755), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT43), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n984), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n984), .A2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n994), .A2(new_n740), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n685), .B1(new_n1027), .B2(new_n660), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT100), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1007), .B2(new_n1000), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n697), .A2(new_n700), .A3(KEYINPUT100), .A4(new_n994), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1028), .B1(new_n1032), .B2(KEYINPUT42), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT42), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1025), .B(new_n1026), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1024), .A3(new_n984), .A4(new_n1035), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n1036), .A2(new_n1038), .B1(new_n698), .B2(new_n1007), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1026), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1025), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n698), .A2(new_n1007), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n1043), .A3(new_n1037), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n987), .B1(new_n1023), .B2(new_n1045), .ZN(G387));
  AOI22_X1  g0846(.A1(new_n708), .A2(new_n758), .B1(new_n527), .B2(new_n703), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n332), .A2(new_n369), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n259), .B1(new_n293), .B2(new_n295), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1050), .A2(new_n708), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n764), .B1(new_n229), .B2(new_n259), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1047), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n773), .ZN(new_n1055));
  INV_X1    g0855(.A(G159), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1056), .A2(new_n791), .B1(new_n805), .B2(new_n330), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n795), .A2(new_n328), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n777), .B2(G68), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n358), .B1(new_n782), .B2(G150), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n788), .A2(G77), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1059), .A2(new_n966), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1057), .B(new_n1062), .C1(G50), .C2(new_n970), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT106), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n358), .B1(new_n792), .B2(new_n781), .C1(new_n813), .C2(new_n451), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n777), .A2(new_n475), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n805), .B2(new_n779), .C1(new_n804), .C2(new_n791), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n970), .B2(G317), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT48), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT48), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n788), .A2(G294), .B1(new_n854), .B2(G283), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1065), .B1(new_n1072), .B2(KEYINPUT49), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1064), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n757), .B(new_n1055), .C1(new_n1077), .C2(new_n839), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1012), .B2(new_n771), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n755), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT107), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n747), .B2(new_n1080), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n747), .A2(new_n1080), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n746), .A2(KEYINPUT107), .A3(new_n1016), .A4(new_n1015), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1083), .A2(new_n704), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1081), .A2(new_n1086), .ZN(G393));
  NAND2_X1  g0887(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1004), .B(new_n994), .C1(new_n1000), .C2(new_n695), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n698), .A3(new_n1002), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1088), .A2(new_n755), .A3(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n803), .A2(new_n1056), .B1(new_n366), .B2(new_n791), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT51), .Z(new_n1095));
  AOI21_X1  g0895(.A(new_n853), .B1(new_n332), .B2(new_n777), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n293), .B2(new_n815), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n358), .B1(new_n854), .B2(G77), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n781), .B2(new_n845), .C1(new_n805), .C2(new_n369), .ZN(new_n1099));
  OR3_X1    g0899(.A1(new_n1095), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n858), .A2(new_n475), .B1(G116), .B2(new_n854), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT108), .Z(new_n1102));
  OAI221_X1 g0902(.A(new_n358), .B1(new_n804), .B2(new_n781), .C1(new_n778), .C2(new_n793), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n788), .A2(G283), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1103), .A2(new_n814), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n970), .A2(G311), .B1(G317), .B2(new_n842), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT52), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1102), .B(new_n1105), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT109), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1100), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n772), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1007), .A2(new_n771), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n773), .B1(new_n457), .B2(new_n206), .C1(new_n239), .C2(new_n765), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1115), .A2(new_n757), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1093), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n698), .B1(new_n1091), .B2(new_n1002), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1084), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n704), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(G390));
  OAI21_X1  g0925(.A(new_n940), .B1(new_n672), .B2(new_n833), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n947), .B1(new_n1126), .B2(new_n906), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT39), .B1(new_n895), .B2(new_n920), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n674), .B1(new_n926), .B2(new_n728), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n863), .A3(new_n906), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n947), .B1(new_n895), .B2(new_n920), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n677), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n742), .B1(new_n1135), .B2(new_n596), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n686), .B(new_n863), .C1(new_n1136), .C2(new_n735), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1137), .A2(new_n940), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT110), .B1(new_n935), .B2(new_n936), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT110), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n901), .A2(new_n1140), .A3(new_n903), .A4(new_n905), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1134), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1131), .A2(new_n1133), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n907), .A2(new_n910), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1146), .A2(new_n922), .A3(new_n674), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1127), .B1(new_n943), .B2(new_n945), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1137), .A2(new_n940), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n921), .A2(new_n946), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1147), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1145), .A2(new_n1152), .A3(new_n755), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT112), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n930), .A2(G330), .A3(new_n927), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n951), .A2(new_n646), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n906), .B1(new_n1132), .B2(new_n863), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1126), .B1(new_n1158), .B2(new_n1147), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1146), .A2(new_n674), .A3(new_n831), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1133), .B(new_n1138), .C1(new_n1160), .C2(new_n1142), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1157), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT111), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1145), .B(new_n1152), .C1(new_n1162), .C2(KEYINPUT111), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n704), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n769), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n757), .B1(new_n383), .B2(new_n840), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n317), .B1(new_n854), .B2(G77), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n793), .B2(new_n781), .C1(new_n778), .C2(new_n457), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n850), .B(new_n1172), .C1(G87), .C2(new_n788), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G107), .A2(new_n858), .B1(new_n842), .B2(G283), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n451), .C2(new_n803), .ZN(new_n1175));
  XOR2_X1   g0975(.A(KEYINPUT54), .B(G143), .Z(new_n1176));
  AOI22_X1  g0976(.A1(new_n777), .A2(new_n1176), .B1(new_n854), .B2(G159), .ZN(new_n1177));
  INV_X1    g0977(.A(G125), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n781), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n788), .A2(G150), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(KEYINPUT53), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT113), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n358), .B1(new_n787), .B2(G50), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n970), .A2(G132), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1181), .B(new_n1184), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n858), .A2(G137), .ZN(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n791), .C1(KEYINPUT53), .C2(new_n1180), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1175), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1170), .B1(new_n1189), .B2(new_n772), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1169), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1155), .A2(new_n1168), .A3(new_n1191), .ZN(G378));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n372), .A2(new_n683), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n382), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n382), .A2(new_n1195), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1193), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1198), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1193), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1200), .A2(new_n1196), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n915), .A2(G330), .A3(new_n1203), .A4(new_n928), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n949), .A2(KEYINPUT116), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n911), .B1(new_n895), .B2(new_n894), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G330), .B(new_n928), .C1(new_n1206), .C2(KEYINPUT40), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1203), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT116), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n942), .A2(new_n948), .A3(new_n1210), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n1204), .A2(new_n1205), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n949), .B1(new_n1209), .B2(new_n1204), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n755), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1203), .A2(new_n769), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n757), .B1(G50), .B2(new_n840), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n358), .A2(new_n258), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n369), .C1(G33), .C2(G41), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT114), .Z(new_n1219));
  OAI22_X1  g1019(.A1(new_n457), .A2(new_n805), .B1(new_n791), .B2(new_n451), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n813), .A2(new_n387), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1217), .B1(new_n854), .B2(G68), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n328), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n777), .A2(new_n1224), .B1(G283), .B2(new_n782), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1222), .A2(new_n1061), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1220), .B(new_n1226), .C1(G107), .C2(new_n970), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1219), .B1(new_n1227), .B2(KEYINPUT58), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n777), .A2(G137), .B1(new_n854), .B2(G150), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n788), .A2(new_n1176), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G132), .B2(new_n858), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n1178), .B2(new_n791), .C1(new_n1187), .C2(new_n803), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(KEYINPUT115), .B(G124), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n241), .B(new_n258), .C1(new_n781), .C2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n787), .B2(new_n843), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1228), .B1(KEYINPUT58), .B2(new_n1227), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1216), .B1(new_n1240), .B2(new_n772), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1215), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT117), .B1(new_n1214), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n949), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n674), .B1(new_n913), .B2(new_n914), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1203), .B1(new_n1245), .B2(new_n928), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1244), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1205), .A2(new_n1209), .A3(new_n1204), .A4(new_n1211), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n754), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT117), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1242), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1243), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1145), .A2(new_n1152), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1157), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1209), .A2(new_n1204), .A3(new_n949), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(KEYINPUT57), .C1(new_n1259), .C2(new_n1213), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1248), .A2(new_n1249), .B1(new_n1257), .B2(new_n1256), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n704), .C1(new_n1261), .C2(KEYINPUT57), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1254), .A2(new_n1262), .ZN(G375));
  NAND3_X1  g1063(.A1(new_n1157), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1163), .A2(new_n1022), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n757), .B1(G68), .B2(new_n840), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1142), .A2(new_n770), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n782), .A2(G303), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n778), .B2(new_n527), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1269), .A2(new_n317), .A3(new_n1058), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n970), .A2(G283), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G77), .A2(new_n787), .B1(new_n788), .B2(G97), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G116), .A2(new_n858), .B1(new_n842), .B2(G294), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n358), .B1(new_n782), .B2(G128), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n369), .B2(new_n795), .C1(new_n778), .C2(new_n366), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1221), .B(new_n1276), .C1(G159), .C2(new_n788), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n970), .A2(G137), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n858), .A2(new_n1176), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n791), .A2(new_n848), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT118), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1274), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1266), .B(new_n1267), .C1(new_n772), .C2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(new_n1255), .B2(new_n755), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1265), .A2(new_n1285), .ZN(G381));
  INV_X1    g1086(.A(G396), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1081), .A2(new_n1086), .A3(new_n1287), .ZN(new_n1288));
  OR4_X1    g1088(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1288), .ZN(new_n1289));
  OR4_X1    g1089(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1289), .ZN(G407));
  INV_X1    g1090(.A(G378), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n684), .A2(G213), .ZN(new_n1292));
  XOR2_X1   g1092(.A(new_n1292), .B(KEYINPUT119), .Z(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G407), .B(G213), .C1(G375), .C2(new_n1294), .ZN(G409));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1264), .B1(new_n1162), .B2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1159), .A2(new_n1157), .A3(new_n1161), .A4(KEYINPUT60), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n704), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n838), .A2(KEYINPUT120), .A3(new_n864), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1285), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT120), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G384), .A2(new_n1302), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1299), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(G2897), .A3(new_n1293), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1303), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1299), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT121), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(KEYINPUT121), .B(new_n1313), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1307), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT122), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G378), .B(new_n1262), .C1(new_n1243), .C2(new_n1253), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1261), .A2(new_n1022), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n755), .B1(new_n1259), .B2(new_n1213), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1242), .A3(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1291), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1292), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT122), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1326), .B(new_n1307), .C1(new_n1314), .C2(new_n1316), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1318), .A2(new_n1325), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1306), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1293), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT126), .B1(new_n1324), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  AOI211_X1 g1133(.A(new_n1333), .B(new_n1293), .C1(new_n1319), .C2(new_n1323), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1330), .B1(new_n1332), .B2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1324), .A2(new_n1292), .A3(new_n1312), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1329), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1288), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1287), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1339));
  OAI21_X1  g1139(.A(KEYINPUT123), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(G393), .A2(G396), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT123), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1288), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1340), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(G390), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G387), .A2(new_n1345), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n987), .B(G390), .C1(new_n1023), .C2(new_n1045), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1344), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1341), .A2(new_n1288), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1019), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1351), .A2(new_n1017), .A3(new_n1011), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1021), .B1(new_n1352), .B2(new_n747), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1044), .B(new_n1039), .C1(new_n1353), .C2(new_n755), .ZN(new_n1354));
  AOI21_X1  g1154(.A(G390), .B1(new_n1354), .B2(new_n987), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1350), .B1(new_n1355), .B2(KEYINPUT124), .ZN(new_n1356));
  AOI21_X1  g1156(.A(KEYINPUT124), .B1(G387), .B2(new_n1345), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1348), .B1(new_n1356), .B2(new_n1358), .ZN(new_n1359));
  OAI21_X1  g1159(.A(KEYINPUT125), .B1(new_n1359), .B2(KEYINPUT61), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT125), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT61), .ZN(new_n1362));
  AND3_X1   g1162(.A1(G387), .A2(KEYINPUT124), .A3(new_n1345), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1363), .A2(new_n1357), .A3(new_n1350), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1361), .B(new_n1362), .C1(new_n1364), .C2(new_n1348), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1360), .A2(new_n1365), .ZN(new_n1366));
  AND4_X1   g1166(.A1(new_n1328), .A2(new_n1335), .A3(new_n1337), .A4(new_n1366), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1359), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1324), .A2(new_n1331), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(new_n1333), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT62), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1317), .A2(new_n1371), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1324), .A2(KEYINPUT126), .A3(new_n1331), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1370), .A2(new_n1372), .A3(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(KEYINPUT61), .B1(new_n1306), .B2(KEYINPUT62), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1375), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1324), .A2(new_n1292), .A3(new_n1312), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1376), .B1(new_n1377), .B2(new_n1371), .ZN(new_n1378));
  AOI21_X1  g1178(.A(new_n1368), .B1(new_n1374), .B2(new_n1378), .ZN(new_n1379));
  OAI21_X1  g1179(.A(KEYINPUT127), .B1(new_n1367), .B2(new_n1379), .ZN(new_n1380));
  AND3_X1   g1180(.A1(new_n1370), .A2(new_n1372), .A3(new_n1373), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1375), .B1(new_n1336), .B2(KEYINPUT62), .ZN(new_n1382));
  OAI21_X1  g1182(.A(new_n1359), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT127), .ZN(new_n1384));
  NAND4_X1  g1184(.A1(new_n1328), .A2(new_n1335), .A3(new_n1366), .A4(new_n1337), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1383), .A2(new_n1384), .A3(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1380), .A2(new_n1386), .ZN(G405));
  AOI21_X1  g1187(.A(G378), .B1(new_n1254), .B2(new_n1262), .ZN(new_n1388));
  INV_X1    g1188(.A(new_n1319), .ZN(new_n1389));
  NOR2_X1   g1189(.A1(new_n1388), .A2(new_n1389), .ZN(new_n1390));
  XNOR2_X1  g1190(.A(new_n1390), .B(new_n1312), .ZN(new_n1391));
  XNOR2_X1  g1191(.A(new_n1391), .B(new_n1368), .ZN(G402));
endmodule


