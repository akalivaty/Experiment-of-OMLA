//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1263, new_n1264,
    new_n1265;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(new_n457), .B(KEYINPUT68), .Z(G261));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT70), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(G2106), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n454), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n453), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT69), .A3(G2106), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n465), .B2(new_n468), .ZN(G319));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n470), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n470), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(new_n478), .ZN(G160));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT71), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2105), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT72), .Z(new_n489));
  INV_X1    g064(.A(G2104), .ZN(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n489), .A2(new_n492), .B1(G136), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n473), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n495), .A2(KEYINPUT4), .A3(G138), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n472), .A2(G126), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  XOR2_X1   g082(.A(KEYINPUT5), .B(G543), .Z(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT75), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n521), .A2(new_n523), .A3(new_n511), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n515), .A2(new_n520), .B1(G88), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n522), .B2(G651), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT74), .A3(G50), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n521), .A2(new_n527), .ZN(new_n531));
  INV_X1    g106(.A(G50), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G166));
  NAND4_X1  g111(.A1(new_n521), .A2(G89), .A3(new_n523), .A4(new_n511), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n521), .A2(G51), .A3(new_n527), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n541), .A2(KEYINPUT76), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT76), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OR2_X1    g122(.A1(KEYINPUT5), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(KEYINPUT5), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(G77), .A2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n520), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n521), .A2(G52), .A3(new_n527), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n521), .A2(G90), .A3(new_n523), .A4(new_n511), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n548), .B2(new_n549), .ZN(new_n558));
  AND2_X1   g133(.A1(G68), .A2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n520), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n521), .A2(G43), .A3(new_n527), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n521), .A2(G81), .A3(new_n523), .A4(new_n511), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT77), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n560), .A2(new_n562), .A3(new_n565), .A4(new_n561), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  NAND3_X1  g148(.A1(new_n521), .A2(G53), .A3(new_n527), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n548), .B2(new_n549), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n521), .A2(KEYINPUT9), .A3(G53), .A4(new_n527), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n521), .A2(G91), .A3(new_n523), .A4(new_n511), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n576), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(G299));
  NAND2_X1  g160(.A1(new_n535), .A2(KEYINPUT79), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n525), .A2(new_n587), .A3(new_n534), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(G303));
  OAI21_X1  g164(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n590));
  INV_X1    g165(.A(G49), .ZN(new_n591));
  INV_X1    g166(.A(G87), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n521), .A2(new_n523), .A3(new_n511), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n590), .B1(new_n531), .B2(new_n591), .C1(new_n592), .C2(new_n593), .ZN(G288));
  AOI22_X1  g169(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n520), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n524), .A2(G86), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n528), .A2(G48), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n524), .A2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n508), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(new_n520), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n528), .A2(G47), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G54), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n609), .A2(new_n516), .B1(new_n531), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n593), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n511), .A2(new_n523), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n616), .A2(G92), .A3(new_n521), .A4(new_n612), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n611), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n608), .B1(new_n618), .B2(G868), .ZN(G321));
  XNOR2_X1  g194(.A(G321), .B(KEYINPUT81), .ZN(G284));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(G299), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G168), .B2(new_n621), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G168), .B2(new_n621), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n618), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g205(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT13), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n495), .A2(G135), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT82), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n486), .A2(G123), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(G2096), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n634), .A2(new_n641), .A3(new_n642), .ZN(G156));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(G14), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n654), .B2(new_n655), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(new_n662), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(new_n663), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n670), .B(new_n664), .C1(new_n660), .C2(new_n663), .ZN(new_n671));
  INV_X1    g246(.A(new_n664), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n660), .A3(new_n663), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g253(.A1(new_n668), .A2(new_n671), .A3(new_n674), .A4(new_n676), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(G227));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT19), .ZN(new_n682));
  NAND2_X1  g257(.A1(G1971), .A2(G1976), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(G1971), .A2(G1976), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G1971), .ZN(new_n687));
  INV_X1    g262(.A(G1976), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n689), .A2(KEYINPUT19), .A3(new_n683), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n695), .B1(new_n691), .B2(new_n694), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n681), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n686), .A2(new_n690), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n692), .A2(new_n693), .ZN(new_n701));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n702), .A2(KEYINPUT20), .A3(new_n696), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n692), .A2(new_n693), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n700), .B(KEYINPUT85), .C1(new_n705), .C2(new_n694), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n686), .A2(new_n690), .A3(KEYINPUT85), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n704), .B(new_n707), .C1(new_n701), .C2(new_n691), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n699), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n699), .A2(new_n703), .A3(new_n709), .A4(new_n711), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(G1991), .B(G1996), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(G1981), .B(G1986), .ZN(new_n718));
  INV_X1    g293(.A(new_n716), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n713), .A2(new_n719), .A3(new_n714), .ZN(new_n720));
  AND3_X1   g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(G229));
  NOR2_X1   g298(.A1(G29), .A2(G33), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT91), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n495), .A2(G139), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT92), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(new_n470), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT25), .Z(new_n731));
  NAND3_X1  g306(.A1(new_n727), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n725), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2072), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT100), .B(G1956), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G16), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT23), .ZN(new_n740));
  INV_X1    g315(.A(G299), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(new_n738), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n735), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n618), .A2(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G4), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n746), .A2(new_n747), .B1(new_n743), .B2(new_n737), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n747), .B2(new_n746), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n733), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT28), .Z(new_n751));
  NAND3_X1  g326(.A1(new_n483), .A2(G128), .A3(new_n485), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G116), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G140), .B2(new_n495), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(G28), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n733), .B1(new_n761), .B2(G28), .ZN(new_n763));
  AND2_X1   g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  NOR2_X1   g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n762), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT24), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n733), .B1(new_n767), .B2(G34), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n767), .B2(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G160), .B2(G29), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n766), .B1(new_n770), .B2(G2084), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n771), .B1(G2084), .B2(new_n770), .C1(new_n733), .C2(new_n640), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n744), .A2(new_n749), .A3(new_n760), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G168), .A2(new_n738), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n738), .B2(G21), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT95), .B(G1966), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n738), .A2(G19), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n568), .B2(new_n738), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT90), .B(G1341), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n733), .A2(G32), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n483), .A2(G129), .A3(new_n485), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT26), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(G141), .B(new_n470), .C1(new_n480), .C2(new_n481), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n783), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n782), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT93), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT94), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n775), .B2(new_n776), .ZN(new_n799));
  NOR2_X1   g374(.A1(G171), .A2(new_n738), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G5), .B2(new_n738), .ZN(new_n801));
  INV_X1    g376(.A(G1961), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2090), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n733), .A2(G35), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT98), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n497), .B2(G29), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n801), .A2(new_n802), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n804), .B2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n733), .A2(G27), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G164), .B2(new_n733), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT97), .B(G2078), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n801), .A2(new_n802), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n812), .A2(new_n814), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n796), .B2(new_n793), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n799), .A2(new_n809), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n773), .A2(new_n777), .A3(new_n781), .A4(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G305), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G16), .ZN(new_n821));
  OR2_X1    g396(.A1(G6), .A2(G16), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT32), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT32), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n821), .A2(new_n825), .A3(new_n822), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1981), .ZN(new_n828));
  NOR2_X1   g403(.A1(G16), .A2(G23), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT87), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G288), .B2(new_n738), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT33), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n688), .ZN(new_n833));
  NOR2_X1   g408(.A1(G16), .A2(G22), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G166), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n687), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n828), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT88), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n828), .A2(KEYINPUT88), .A3(new_n833), .A4(new_n836), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(KEYINPUT34), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n483), .A2(G119), .A3(new_n485), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(G107), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(G2105), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G131), .B2(new_n495), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G29), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(G25), .B2(G29), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G1991), .Z(new_n851));
  AOI21_X1  g426(.A(KEYINPUT89), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n738), .A2(G24), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT86), .Z(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G290), .B2(G16), .ZN(new_n856));
  INV_X1    g431(.A(G1986), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n841), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT34), .B1(new_n839), .B2(new_n840), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT36), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n839), .A2(new_n840), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT34), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n841), .A4(new_n859), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n819), .B1(new_n862), .B2(new_n867), .ZN(G311));
  NAND2_X1  g443(.A1(new_n862), .A2(new_n867), .ZN(new_n869));
  INV_X1    g444(.A(new_n819), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(G150));
  AOI22_X1  g446(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(new_n596), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n521), .A2(G93), .A3(new_n523), .A4(new_n511), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n521), .A2(G55), .A3(new_n527), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n874), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n567), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n875), .A2(new_n877), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT101), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n563), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n874), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT38), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n615), .A2(new_n617), .ZN(new_n890));
  INV_X1    g465(.A(new_n611), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(new_n625), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n889), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n895));
  AOI21_X1  g470(.A(G860), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n880), .A2(G860), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT37), .Z(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(G145));
  XNOR2_X1  g475(.A(G160), .B(KEYINPUT102), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(G162), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n903));
  XNOR2_X1  g478(.A(G160), .B(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(new_n497), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n640), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(G162), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n497), .ZN(new_n908));
  INV_X1    g483(.A(new_n640), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n842), .A2(KEYINPUT103), .A3(new_n846), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT103), .B1(new_n842), .B2(new_n846), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n632), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n847), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n632), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n842), .A2(new_n846), .A3(KEYINPUT103), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n486), .A2(G130), .ZN(new_n922));
  OAI21_X1  g497(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n923));
  INV_X1    g498(.A(G118), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(G2105), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(G142), .B2(new_n495), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n916), .A2(new_n921), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n916), .B2(new_n921), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n913), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n914), .A2(new_n915), .A3(new_n632), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n916), .A2(new_n921), .A3(new_n928), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(KEYINPUT104), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n792), .A2(new_n757), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n783), .A2(new_n752), .A3(new_n791), .A4(new_n756), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n937), .A2(new_n506), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n506), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n732), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n938), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n783), .A2(new_n791), .B1(new_n752), .B2(new_n756), .ZN(new_n943));
  OAI21_X1  g518(.A(G164), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n732), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n506), .A3(new_n938), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n931), .A2(new_n936), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n931), .B2(new_n936), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(new_n950), .B2(KEYINPUT105), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  AOI211_X1 g527(.A(new_n952), .B(new_n948), .C1(new_n936), .C2(new_n931), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n912), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n949), .A2(new_n911), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n929), .A2(new_n930), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n948), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n934), .A2(new_n935), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(KEYINPUT106), .A3(new_n947), .A4(new_n941), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g539(.A(new_n627), .B(KEYINPUT107), .Z(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(new_n888), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n890), .A2(G299), .A3(new_n891), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n618), .A2(KEYINPUT108), .A3(G299), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n892), .A2(KEYINPUT109), .A3(new_n741), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n618), .B2(G299), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n971), .A2(KEYINPUT41), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n972), .A3(new_n967), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT41), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n967), .A2(new_n968), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT108), .B1(new_n618), .B2(G299), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n974), .A2(new_n972), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n980), .B1(new_n966), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(KEYINPUT111), .A3(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g562(.A1(G166), .A2(new_n820), .ZN(new_n988));
  AND2_X1   g563(.A1(G290), .A2(G288), .ZN(new_n989));
  NOR2_X1   g564(.A1(G290), .A2(G288), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT110), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(G290), .A2(G288), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n993));
  NAND2_X1  g568(.A1(G290), .A2(G288), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n535), .A2(G305), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n988), .A2(new_n991), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n989), .A2(new_n990), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n820), .B1(new_n525), .B2(new_n534), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n535), .A2(G305), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n993), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI221_X1 g580(.A(new_n980), .B1(new_n1003), .B2(new_n1004), .C1(new_n966), .C2(new_n985), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n987), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1005), .B1(new_n987), .B2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g583(.A(G868), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n880), .A2(new_n621), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(G295));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1010), .ZN(G331));
  AOI22_X1  g587(.A1(new_n885), .A2(new_n874), .B1(new_n564), .B2(new_n566), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n873), .B(new_n563), .C1(new_n883), .C2(new_n884), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n541), .A2(new_n542), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT76), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n541), .A2(KEYINPUT76), .A3(new_n542), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(G301), .B1(new_n1019), .B2(new_n540), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n540), .B(G301), .C1(new_n543), .C2(new_n544), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n1013), .A2(new_n1014), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G286), .A2(G171), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n881), .A2(new_n887), .A3(new_n1024), .A4(new_n1021), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(KEYINPUT41), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n985), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1023), .A2(new_n976), .A3(new_n1025), .A4(KEYINPUT41), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1002), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1027), .A2(new_n1002), .A3(KEYINPUT112), .A4(new_n1028), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n974), .A2(new_n972), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1025), .A2(new_n1023), .B1(new_n1034), .B2(new_n971), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1035), .B1(new_n979), .B2(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n997), .A2(new_n1001), .ZN(new_n1039));
  AOI21_X1  g614(.A(G37), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1033), .A2(new_n1040), .A3(KEYINPUT113), .A4(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1033), .A2(new_n1041), .A3(new_n1040), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1036), .B1(new_n978), .B2(new_n975), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1002), .B1(new_n1045), .B2(new_n1035), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n979), .A2(new_n1037), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1036), .B1(new_n984), .B2(new_n983), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1039), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G37), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1044), .B1(new_n1051), .B2(KEYINPUT43), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1042), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1033), .A2(KEYINPUT43), .A3(new_n1040), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1041), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  MUX2_X1   g631(.A(new_n1053), .B(new_n1056), .S(KEYINPUT44), .Z(G397));
  INV_X1    g632(.A(G1384), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n506), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT114), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n506), .A2(new_n1062), .A3(new_n1058), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(G160), .A2(G40), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(KEYINPUT50), .B2(new_n1059), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1348), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1065), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1060), .A2(new_n1068), .A3(new_n1063), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G2067), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n618), .ZN(new_n1072));
  XOR2_X1   g647(.A(G299), .B(KEYINPUT57), .Z(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT119), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n1058), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1068), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT45), .B1(new_n506), .B2(new_n1058), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n506), .A2(new_n1062), .A3(new_n1058), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1062), .B1(new_n506), .B2(new_n1058), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT50), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n506), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n506), .A2(KEYINPUT117), .A3(new_n1061), .A4(new_n1058), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1083), .A2(new_n1088), .A3(new_n1068), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1080), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1074), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT118), .B(new_n1080), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1072), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1080), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1073), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1091), .A2(KEYINPUT61), .A3(new_n1073), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1071), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1081), .A2(new_n1082), .A3(new_n1065), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1106), .A2(new_n747), .B1(new_n759), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n892), .B1(new_n1108), .B2(KEYINPUT60), .ZN(new_n1109));
  NOR4_X1   g684(.A1(new_n1067), .A2(new_n1070), .A3(new_n1104), .A4(new_n618), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1103), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT45), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1059), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G1996), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n1068), .A4(new_n1075), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT58), .B(G1341), .Z(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT120), .B(new_n1116), .C1(new_n1107), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1069), .A2(new_n1117), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT120), .B1(new_n1121), .B2(new_n1116), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n568), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n568), .B(new_n1124), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n1091), .A2(new_n1073), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1099), .B1(new_n1112), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n1131));
  INV_X1    g706(.A(G2078), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1114), .A2(new_n1132), .A3(new_n1068), .A4(new_n1075), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1106), .A2(new_n802), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1113), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1068), .A2(new_n1075), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(KEYINPUT53), .A4(new_n1132), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(G301), .B(KEYINPUT54), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1132), .A2(KEYINPUT123), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1132), .A2(KEYINPUT123), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1131), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1138), .A2(new_n1139), .B1(new_n1134), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1106), .A2(G2084), .ZN(new_n1146));
  INV_X1    g721(.A(new_n776), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1148));
  OAI21_X1  g723(.A(G8), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT51), .ZN(new_n1150));
  NAND2_X1  g725(.A1(G286), .A2(G8), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT122), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1149), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1152), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT51), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1157), .A2(new_n1147), .B1(new_n1106), .B2(G2084), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1154), .B1(new_n1158), .B2(G8), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1145), .B(new_n1153), .C1(new_n1156), .C2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n687), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1106), .B2(G2090), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1162), .A2(G8), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n586), .A2(G8), .A3(new_n588), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT55), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n586), .A2(KEYINPUT55), .A3(G8), .A4(new_n588), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1166), .A2(KEYINPUT115), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT115), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(G288), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(G1976), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT52), .B1(G288), .B2(new_n688), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1069), .A2(G8), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1069), .A2(G8), .A3(new_n1172), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(KEYINPUT52), .ZN(new_n1176));
  NAND2_X1  g751(.A1(G305), .A2(G1981), .ZN(new_n1177));
  INV_X1    g752(.A(G1981), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n597), .A2(new_n598), .A3(new_n1178), .A4(new_n599), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(KEYINPUT49), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT49), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1181), .A2(KEYINPUT116), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT116), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1183), .B(KEYINPUT49), .C1(new_n1177), .C2(new_n1179), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1180), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1069), .A2(G8), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1174), .B(new_n1176), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1161), .B1(new_n1089), .B2(G2090), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(G8), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1170), .A2(new_n1188), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1160), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1130), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1149), .A2(G286), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1170), .A2(new_n1188), .A3(new_n1192), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1163), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n1191), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1149), .A2(new_n1198), .A3(G286), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1201), .A2(new_n1170), .A3(new_n1188), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1153), .B1(new_n1159), .B2(new_n1156), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AND3_X1   g782(.A1(new_n1170), .A2(new_n1192), .A3(new_n1188), .ZN(new_n1208));
  AOI21_X1  g783(.A(G301), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1209));
  OAI211_X1 g784(.A(KEYINPUT62), .B(new_n1153), .C1(new_n1159), .C2(new_n1156), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1170), .A2(new_n1187), .ZN(new_n1212));
  OAI211_X1 g787(.A(new_n688), .B(new_n1171), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1186), .B1(new_n1213), .B2(new_n1179), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1195), .A2(new_n1204), .A3(new_n1211), .A4(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n792), .B(new_n1115), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n757), .A2(G2067), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n752), .A2(new_n756), .A3(new_n759), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n847), .B(new_n851), .Z(new_n1221));
  NOR2_X1   g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(G290), .B(new_n857), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1114), .A2(new_n1065), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1216), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1225), .A2(new_n1115), .ZN(new_n1228));
  XNOR2_X1  g803(.A(new_n1228), .B(KEYINPUT46), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1225), .B1(new_n792), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1232), .B(KEYINPUT47), .ZN(new_n1233));
  XNOR2_X1  g808(.A(new_n1233), .B(KEYINPUT125), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n848), .A2(new_n851), .ZN(new_n1235));
  XOR2_X1   g810(.A(new_n1235), .B(KEYINPUT124), .Z(new_n1236));
  OAI21_X1  g811(.A(new_n1219), .B1(new_n1236), .B2(new_n1220), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1237), .A2(new_n1225), .ZN(new_n1238));
  INV_X1    g813(.A(new_n1225), .ZN(new_n1239));
  NOR2_X1   g814(.A1(new_n1222), .A2(new_n1239), .ZN(new_n1240));
  NOR3_X1   g815(.A1(new_n1239), .A2(G1986), .A3(G290), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1240), .B1(KEYINPUT48), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1242), .B1(KEYINPUT48), .B2(new_n1241), .ZN(new_n1243));
  AND3_X1   g818(.A1(new_n1234), .A2(new_n1238), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g819(.A1(new_n1227), .A2(new_n1244), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g820(.A(KEYINPUT127), .ZN(new_n1247));
  NAND3_X1  g821(.A1(new_n678), .A2(G319), .A3(new_n679), .ZN(new_n1248));
  AOI21_X1  g822(.A(new_n1248), .B1(new_n656), .B2(new_n658), .ZN(new_n1249));
  OAI21_X1  g823(.A(new_n1249), .B1(new_n721), .B2(new_n722), .ZN(new_n1250));
  NAND2_X1  g824(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1251));
  INV_X1    g825(.A(KEYINPUT126), .ZN(new_n1252));
  OAI211_X1 g826(.A(new_n1249), .B(new_n1252), .C1(new_n721), .C2(new_n722), .ZN(new_n1253));
  NAND2_X1  g827(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g828(.A1(new_n963), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g829(.A1(new_n1033), .A2(new_n1041), .A3(new_n1040), .ZN(new_n1256));
  AOI21_X1  g830(.A(new_n1041), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1257));
  OAI21_X1  g831(.A(new_n1256), .B1(new_n1257), .B2(new_n1044), .ZN(new_n1258));
  AOI211_X1 g832(.A(new_n1247), .B(new_n1255), .C1(new_n1258), .C2(new_n1042), .ZN(new_n1259));
  INV_X1    g833(.A(new_n1255), .ZN(new_n1260));
  AOI21_X1  g834(.A(KEYINPUT127), .B1(new_n1053), .B2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g835(.A1(new_n1259), .A2(new_n1261), .ZN(G308));
  NAND2_X1  g836(.A1(new_n1053), .A2(new_n1260), .ZN(new_n1263));
  NAND2_X1  g837(.A1(new_n1263), .A2(new_n1247), .ZN(new_n1264));
  NAND3_X1  g838(.A1(new_n1053), .A2(KEYINPUT127), .A3(new_n1260), .ZN(new_n1265));
  NAND2_X1  g839(.A1(new_n1264), .A2(new_n1265), .ZN(G225));
endmodule


