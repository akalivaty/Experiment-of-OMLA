

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582;

  INV_X1 U322 ( .A(n498), .ZN(n560) );
  XNOR2_X1 U323 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n504) );
  XNOR2_X1 U324 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n325) );
  OR2_X1 U325 ( .A1(n293), .A2(n360), .ZN(n294) );
  XNOR2_X1 U326 ( .A(n505), .B(n504), .ZN(n511) );
  XNOR2_X1 U327 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U328 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U329 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n447) );
  NOR2_X1 U330 ( .A1(n544), .A2(n543), .ZN(n568) );
  XOR2_X1 U331 ( .A(n572), .B(KEYINPUT41), .Z(n529) );
  XNOR2_X1 U332 ( .A(n448), .B(n447), .ZN(n490) );
  XNOR2_X1 U333 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n449) );
  XNOR2_X1 U334 ( .A(n306), .B(n305), .ZN(n572) );
  AND2_X1 U335 ( .A1(n560), .A2(n562), .ZN(n556) );
  XNOR2_X1 U336 ( .A(n450), .B(n449), .ZN(n477) );
  XNOR2_X1 U337 ( .A(n455), .B(G50GAT), .ZN(n456) );
  XNOR2_X1 U338 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U339 ( .A(n457), .B(n456), .ZN(G1331GAT) );
  XNOR2_X1 U340 ( .A(G99GAT), .B(G71GAT), .ZN(n290) );
  XNOR2_X1 U341 ( .A(n290), .B(G120GAT), .ZN(n329) );
  XOR2_X1 U342 ( .A(G57GAT), .B(KEYINPUT13), .Z(n411) );
  XNOR2_X1 U343 ( .A(n329), .B(n411), .ZN(n292) );
  NAND2_X1 U344 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U346 ( .A(G148GAT), .B(G78GAT), .Z(n360) );
  NAND2_X1 U347 ( .A1(n293), .A2(n360), .ZN(n295) );
  NAND2_X1 U348 ( .A1(n295), .A2(n294), .ZN(n297) );
  XNOR2_X1 U349 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n296) );
  XOR2_X1 U350 ( .A(n297), .B(n296), .Z(n301) );
  XOR2_X1 U351 ( .A(KEYINPUT70), .B(KEYINPUT72), .Z(n299) );
  XNOR2_X1 U352 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n306) );
  XNOR2_X1 U355 ( .A(G85GAT), .B(KEYINPUT69), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n302), .B(G106GAT), .ZN(n436) );
  XOR2_X1 U357 ( .A(G204GAT), .B(G64GAT), .Z(n304) );
  XNOR2_X1 U358 ( .A(G176GAT), .B(G92GAT), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n347) );
  XNOR2_X1 U360 ( .A(n436), .B(n347), .ZN(n305) );
  XOR2_X1 U361 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n308) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(KEYINPUT29), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n316) );
  XOR2_X1 U364 ( .A(G36GAT), .B(G8GAT), .Z(n352) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(G15GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n309), .B(G113GAT), .ZN(n324) );
  XOR2_X1 U367 ( .A(n352), .B(n324), .Z(n311) );
  NAND2_X1 U368 ( .A1(G229GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U370 ( .A(G22GAT), .B(G141GAT), .Z(n361) );
  XOR2_X1 U371 ( .A(n312), .B(n361), .Z(n314) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(G197GAT), .ZN(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U375 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n318) );
  XNOR2_X1 U376 ( .A(G50GAT), .B(G29GAT), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U378 ( .A(KEYINPUT66), .B(n319), .Z(n441) );
  XNOR2_X1 U379 ( .A(n320), .B(n441), .ZN(n569) );
  XOR2_X1 U380 ( .A(KEYINPUT68), .B(n569), .Z(n547) );
  NAND2_X1 U381 ( .A1(n572), .A2(n547), .ZN(n321) );
  XOR2_X1 U382 ( .A(KEYINPUT73), .B(n321), .Z(n465) );
  XOR2_X1 U383 ( .A(KEYINPUT0), .B(KEYINPUT80), .Z(n323) );
  XNOR2_X1 U384 ( .A(G134GAT), .B(G127GAT), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n323), .B(n322), .ZN(n383) );
  XNOR2_X1 U386 ( .A(n324), .B(n383), .ZN(n341) );
  XNOR2_X1 U387 ( .A(n325), .B(KEYINPUT17), .ZN(n326) );
  XOR2_X1 U388 ( .A(KEYINPUT84), .B(n326), .Z(n328) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(G183GAT), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n328), .B(n327), .ZN(n351) );
  XNOR2_X1 U391 ( .A(n351), .B(n329), .ZN(n337) );
  XOR2_X1 U392 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n331) );
  XNOR2_X1 U393 ( .A(KEYINPUT83), .B(KEYINPUT81), .ZN(n330) );
  XNOR2_X1 U394 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U395 ( .A(G190GAT), .B(G176GAT), .Z(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n335) );
  XOR2_X1 U397 ( .A(KEYINPUT64), .B(KEYINPUT82), .Z(n334) );
  NAND2_X1 U398 ( .A1(G227GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n498) );
  XOR2_X1 U401 ( .A(KEYINPUT93), .B(KEYINPUT95), .Z(n343) );
  NAND2_X1 U402 ( .A1(G226GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U404 ( .A(n344), .B(KEYINPUT94), .Z(n349) );
  XOR2_X1 U405 ( .A(KEYINPUT21), .B(G211GAT), .Z(n346) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(G218GAT), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n369) );
  XNOR2_X1 U408 ( .A(n347), .B(n369), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U410 ( .A(G190GAT), .B(KEYINPUT76), .Z(n437) );
  XOR2_X1 U411 ( .A(n350), .B(n437), .Z(n354) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n538) );
  NAND2_X1 U414 ( .A1(n560), .A2(n538), .ZN(n373) );
  XOR2_X1 U415 ( .A(G155GAT), .B(G162GAT), .Z(n356) );
  XNOR2_X1 U416 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U418 ( .A(KEYINPUT2), .B(n357), .Z(n382) );
  XOR2_X1 U419 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n359) );
  XNOR2_X1 U420 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n365) );
  XOR2_X1 U422 ( .A(n360), .B(G106GAT), .Z(n363) );
  XNOR2_X1 U423 ( .A(G50GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U425 ( .A(n365), .B(n364), .Z(n367) );
  NAND2_X1 U426 ( .A1(G228GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U428 ( .A(n368), .B(KEYINPUT87), .Z(n371) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT89), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n382), .B(n372), .ZN(n545) );
  NAND2_X1 U432 ( .A1(n373), .A2(n545), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n374), .B(KEYINPUT25), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n375), .B(KEYINPUT97), .ZN(n379) );
  NOR2_X1 U435 ( .A1(n560), .A2(n545), .ZN(n377) );
  XNOR2_X1 U436 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n567) );
  XNOR2_X1 U438 ( .A(n538), .B(KEYINPUT27), .ZN(n402) );
  NAND2_X1 U439 ( .A1(n567), .A2(n402), .ZN(n378) );
  NAND2_X1 U440 ( .A1(n379), .A2(n378), .ZN(n401) );
  XOR2_X1 U441 ( .A(KEYINPUT90), .B(G148GAT), .Z(n381) );
  XNOR2_X1 U442 ( .A(G141GAT), .B(G113GAT), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n387) );
  XOR2_X1 U444 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n385) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n399) );
  NAND2_X1 U448 ( .A1(G225GAT), .A2(G233GAT), .ZN(n393) );
  XOR2_X1 U449 ( .A(G57GAT), .B(KEYINPUT75), .Z(n389) );
  XNOR2_X1 U450 ( .A(G1GAT), .B(G120GAT), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U452 ( .A(G29GAT), .B(G85GAT), .Z(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U455 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n395) );
  XNOR2_X1 U456 ( .A(KEYINPUT5), .B(KEYINPUT92), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n544) );
  INV_X1 U460 ( .A(n544), .ZN(n400) );
  NAND2_X1 U461 ( .A1(n401), .A2(n400), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n498), .B(KEYINPUT86), .ZN(n405) );
  NAND2_X1 U463 ( .A1(n544), .A2(n402), .ZN(n513) );
  XNOR2_X1 U464 ( .A(KEYINPUT65), .B(KEYINPUT28), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n403), .B(n545), .ZN(n497) );
  NOR2_X1 U466 ( .A1(n513), .A2(n497), .ZN(n404) );
  NAND2_X1 U467 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U468 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n408), .B(KEYINPUT98), .ZN(n463) );
  XOR2_X1 U470 ( .A(G64GAT), .B(G211GAT), .Z(n410) );
  XNOR2_X1 U471 ( .A(G8GAT), .B(G183GAT), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n412) );
  XOR2_X1 U473 ( .A(n412), .B(n411), .Z(n414) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(G15GAT), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n427) );
  XOR2_X1 U476 ( .A(KEYINPUT14), .B(G78GAT), .Z(n416) );
  NAND2_X1 U477 ( .A1(G231GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U479 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n418) );
  XNOR2_X1 U480 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U482 ( .A(n420), .B(n419), .Z(n425) );
  XOR2_X1 U483 ( .A(KEYINPUT78), .B(G155GAT), .Z(n422) );
  XNOR2_X1 U484 ( .A(G22GAT), .B(G127GAT), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U486 ( .A(G71GAT), .B(n423), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n557) );
  XOR2_X1 U489 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n429) );
  XNOR2_X1 U490 ( .A(G162GAT), .B(KEYINPUT75), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n445) );
  XOR2_X1 U492 ( .A(KEYINPUT10), .B(G218GAT), .Z(n431) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(G134GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U495 ( .A(KEYINPUT9), .B(G92GAT), .Z(n433) );
  XNOR2_X1 U496 ( .A(G36GAT), .B(G99GAT), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U498 ( .A(n435), .B(n434), .Z(n443) );
  XOR2_X1 U499 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U500 ( .A1(G232GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n559) );
  INV_X1 U505 ( .A(n559), .ZN(n536) );
  XNOR2_X1 U506 ( .A(n536), .B(KEYINPUT36), .ZN(n580) );
  NOR2_X1 U507 ( .A1(n557), .A2(n580), .ZN(n446) );
  NAND2_X1 U508 ( .A1(n463), .A2(n446), .ZN(n448) );
  NOR2_X1 U509 ( .A1(n465), .A2(n490), .ZN(n450) );
  NAND2_X1 U510 ( .A1(n477), .A2(n560), .ZN(n454) );
  XOR2_X1 U511 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n452) );
  INV_X1 U512 ( .A(G43GAT), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  NAND2_X1 U514 ( .A1(n477), .A2(n497), .ZN(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n455) );
  INV_X1 U516 ( .A(G29GAT), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n477), .A2(n544), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(G1328GAT) );
  XOR2_X1 U521 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n467) );
  INV_X1 U522 ( .A(n557), .ZN(n575) );
  NOR2_X1 U523 ( .A1(n575), .A2(n559), .ZN(n462) );
  XNOR2_X1 U524 ( .A(KEYINPUT16), .B(n462), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n464), .A2(n463), .ZN(n479) );
  NOR2_X1 U526 ( .A1(n465), .A2(n479), .ZN(n473) );
  NAND2_X1 U527 ( .A1(n473), .A2(n544), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n468), .ZN(G1324GAT) );
  NAND2_X1 U530 ( .A1(n473), .A2(n538), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n469), .B(KEYINPUT100), .ZN(n470) );
  XNOR2_X1 U532 ( .A(G8GAT), .B(n470), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .Z(n472) );
  NAND2_X1 U534 ( .A1(n473), .A2(n560), .ZN(n471) );
  XNOR2_X1 U535 ( .A(n472), .B(n471), .ZN(G1326GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n475) );
  NAND2_X1 U537 ( .A1(n473), .A2(n497), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n476), .ZN(G1327GAT) );
  NAND2_X1 U540 ( .A1(n477), .A2(n538), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n478), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U542 ( .A(n529), .B(KEYINPUT109), .ZN(n553) );
  NAND2_X1 U543 ( .A1(n569), .A2(n553), .ZN(n489) );
  NOR2_X1 U544 ( .A1(n479), .A2(n489), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n480), .B(KEYINPUT110), .ZN(n485) );
  NAND2_X1 U546 ( .A1(n544), .A2(n485), .ZN(n481) );
  XNOR2_X1 U547 ( .A(KEYINPUT42), .B(n481), .ZN(n482) );
  XNOR2_X1 U548 ( .A(G57GAT), .B(n482), .ZN(G1332GAT) );
  NAND2_X1 U549 ( .A1(n485), .A2(n538), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n483), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U551 ( .A1(n485), .A2(n560), .ZN(n484) );
  XNOR2_X1 U552 ( .A(n484), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n487) );
  NAND2_X1 U554 ( .A1(n485), .A2(n497), .ZN(n486) );
  XNOR2_X1 U555 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U556 ( .A(G78GAT), .B(n488), .Z(G1335GAT) );
  NOR2_X1 U557 ( .A1(n490), .A2(n489), .ZN(n494) );
  NAND2_X1 U558 ( .A1(n544), .A2(n494), .ZN(n491) );
  XNOR2_X1 U559 ( .A(G85GAT), .B(n491), .ZN(G1336GAT) );
  NAND2_X1 U560 ( .A1(n494), .A2(n538), .ZN(n492) );
  XNOR2_X1 U561 ( .A(n492), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U562 ( .A1(n560), .A2(n494), .ZN(n493) );
  XNOR2_X1 U563 ( .A(n493), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U564 ( .A1(n497), .A2(n494), .ZN(n495) );
  XNOR2_X1 U565 ( .A(n495), .B(KEYINPUT44), .ZN(n496) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(n496), .ZN(G1339GAT) );
  NOR2_X1 U567 ( .A1(n498), .A2(n497), .ZN(n514) );
  INV_X1 U568 ( .A(KEYINPUT112), .ZN(n502) );
  NOR2_X1 U569 ( .A1(n569), .A2(n529), .ZN(n499) );
  XNOR2_X1 U570 ( .A(n499), .B(KEYINPUT46), .ZN(n500) );
  NOR2_X1 U571 ( .A1(n500), .A2(n557), .ZN(n501) );
  XNOR2_X1 U572 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U573 ( .A1(n503), .A2(n559), .ZN(n505) );
  NOR2_X1 U574 ( .A1(n575), .A2(n580), .ZN(n507) );
  XNOR2_X1 U575 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n506) );
  XNOR2_X1 U576 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U577 ( .A1(n572), .A2(n508), .ZN(n509) );
  NOR2_X1 U578 ( .A1(n547), .A2(n509), .ZN(n510) );
  NOR2_X1 U579 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U580 ( .A(KEYINPUT48), .B(n512), .ZN(n540) );
  NOR2_X1 U581 ( .A1(n540), .A2(n513), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n514), .A2(n526), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(KEYINPUT115), .ZN(n522) );
  NAND2_X1 U584 ( .A1(n522), .A2(n547), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n516), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n518) );
  NAND2_X1 U587 ( .A1(n522), .A2(n553), .ZN(n517) );
  XNOR2_X1 U588 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U589 ( .A(G120GAT), .B(n519), .ZN(G1341GAT) );
  NAND2_X1 U590 ( .A1(n557), .A2(n522), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n520), .B(KEYINPUT50), .ZN(n521) );
  XNOR2_X1 U592 ( .A(G127GAT), .B(n521), .ZN(G1342GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n524) );
  NAND2_X1 U594 ( .A1(n522), .A2(n559), .ZN(n523) );
  XNOR2_X1 U595 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U596 ( .A(G134GAT), .B(n525), .Z(G1343GAT) );
  NAND2_X1 U597 ( .A1(n567), .A2(n526), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n569), .A2(n535), .ZN(n527) );
  XOR2_X1 U599 ( .A(G141GAT), .B(n527), .Z(n528) );
  XNOR2_X1 U600 ( .A(KEYINPUT118), .B(n528), .ZN(G1344GAT) );
  NOR2_X1 U601 ( .A1(n529), .A2(n535), .ZN(n531) );
  XNOR2_X1 U602 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n530) );
  XNOR2_X1 U603 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U604 ( .A(G148GAT), .B(n532), .ZN(G1345GAT) );
  NOR2_X1 U605 ( .A1(n575), .A2(n535), .ZN(n534) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n533) );
  XNOR2_X1 U607 ( .A(n534), .B(n533), .ZN(G1346GAT) );
  NOR2_X1 U608 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U609 ( .A(G162GAT), .B(n537), .Z(G1347GAT) );
  XOR2_X1 U610 ( .A(G169GAT), .B(KEYINPUT121), .Z(n549) );
  INV_X1 U611 ( .A(KEYINPUT54), .ZN(n542) );
  XOR2_X1 U612 ( .A(KEYINPUT120), .B(n538), .Z(n539) );
  NOR2_X1 U613 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U614 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U615 ( .A1(n568), .A2(n545), .ZN(n546) );
  XNOR2_X1 U616 ( .A(KEYINPUT55), .B(n546), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n556), .A2(n547), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n551) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n550) );
  XNOR2_X1 U621 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(n552), .Z(n555) );
  NAND2_X1 U623 ( .A1(n556), .A2(n553), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT58), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n579) );
  NOR2_X1 U635 ( .A1(n569), .A2(n579), .ZN(n570) );
  XOR2_X1 U636 ( .A(n571), .B(n570), .Z(G1352GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n579), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n579), .ZN(n576) );
  XOR2_X1 U641 ( .A(G211GAT), .B(n576), .Z(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

