

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NOR2_X1 U559 ( .A1(G651), .A2(n658), .ZN(n667) );
  NOR2_X2 U560 ( .A1(n989), .A2(n719), .ZN(n705) );
  XNOR2_X2 U561 ( .A(n703), .B(n702), .ZN(n719) );
  AND2_X1 U562 ( .A1(n753), .A2(n752), .ZN(n755) );
  AND2_X2 U563 ( .A1(n526), .A2(G2105), .ZN(n910) );
  XNOR2_X1 U564 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n525) );
  INV_X1 U565 ( .A(KEYINPUT64), .ZN(n533) );
  INV_X1 U566 ( .A(KEYINPUT98), .ZN(n702) );
  NAND2_X1 U567 ( .A1(n697), .A2(n804), .ZN(n734) );
  INV_X1 U568 ( .A(KEYINPUT13), .ZN(n604) );
  AND2_X2 U569 ( .A1(n538), .A2(n537), .ZN(G160) );
  OR2_X1 U570 ( .A1(n791), .A2(n790), .ZN(n523) );
  INV_X2 U571 ( .A(G2104), .ZN(n526) );
  INV_X1 U572 ( .A(KEYINPUT27), .ZN(n698) );
  INV_X1 U573 ( .A(n734), .ZN(n706) );
  INV_X1 U574 ( .A(KEYINPUT101), .ZN(n732) );
  BUF_X1 U575 ( .A(n734), .Z(n746) );
  XNOR2_X1 U576 ( .A(KEYINPUT32), .B(KEYINPUT104), .ZN(n754) );
  XNOR2_X1 U577 ( .A(n599), .B(KEYINPUT73), .ZN(n600) );
  INV_X1 U578 ( .A(KEYINPUT106), .ZN(n828) );
  INV_X1 U579 ( .A(KEYINPUT77), .ZN(n618) );
  XNOR2_X1 U580 ( .A(n601), .B(n600), .ZN(n603) );
  XNOR2_X1 U581 ( .A(n618), .B(KEYINPUT15), .ZN(n619) );
  INV_X2 U582 ( .A(G2105), .ZN(n531) );
  XNOR2_X1 U583 ( .A(n620), .B(n619), .ZN(n714) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n662) );
  XNOR2_X1 U585 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U586 ( .A(n534), .B(n533), .ZN(n535) );
  INV_X1 U587 ( .A(KEYINPUT66), .ZN(n529) );
  NOR2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n564) );
  NAND2_X1 U590 ( .A1(n564), .A2(G137), .ZN(n528) );
  NOR2_X4 U591 ( .A1(n526), .A2(n531), .ZN(n909) );
  NAND2_X1 U592 ( .A1(G113), .A2(n909), .ZN(n527) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n538) );
  AND2_X4 U595 ( .A1(n531), .A2(G2104), .ZN(n915) );
  NAND2_X1 U596 ( .A1(G101), .A2(n915), .ZN(n532) );
  XNOR2_X1 U597 ( .A(KEYINPUT23), .B(n532), .ZN(n536) );
  NAND2_X1 U598 ( .A1(G125), .A2(n910), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n915), .A2(G102), .ZN(n539) );
  XNOR2_X1 U600 ( .A(n539), .B(KEYINPUT84), .ZN(n541) );
  NAND2_X1 U601 ( .A1(G138), .A2(n564), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n542), .B(KEYINPUT85), .ZN(n546) );
  NAND2_X1 U604 ( .A1(G114), .A2(n909), .ZN(n544) );
  NAND2_X1 U605 ( .A1(G126), .A2(n910), .ZN(n543) );
  AND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n545) );
  AND2_X2 U607 ( .A1(n546), .A2(n545), .ZN(G164) );
  NAND2_X1 U608 ( .A1(G85), .A2(n662), .ZN(n548) );
  XOR2_X1 U609 ( .A(KEYINPUT0), .B(G543), .Z(n658) );
  INV_X1 U610 ( .A(G651), .ZN(n549) );
  NOR2_X2 U611 ( .A1(n658), .A2(n549), .ZN(n661) );
  NAND2_X1 U612 ( .A1(G72), .A2(n661), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n554) );
  NOR2_X1 U614 ( .A1(G543), .A2(n549), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT1), .B(n550), .Z(n666) );
  NAND2_X1 U616 ( .A1(G60), .A2(n666), .ZN(n552) );
  NAND2_X1 U617 ( .A1(G47), .A2(n667), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  OR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(G290) );
  XOR2_X1 U620 ( .A(G2443), .B(G2446), .Z(n556) );
  XNOR2_X1 U621 ( .A(G2427), .B(G2451), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n562) );
  XOR2_X1 U623 ( .A(G2430), .B(G2454), .Z(n558) );
  XNOR2_X1 U624 ( .A(G1341), .B(G1348), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n560) );
  XOR2_X1 U626 ( .A(G2435), .B(G2438), .Z(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(n562), .B(n561), .Z(n563) );
  AND2_X1 U629 ( .A1(G14), .A2(n563), .ZN(G401) );
  BUF_X1 U630 ( .A(n564), .Z(n913) );
  NAND2_X1 U631 ( .A1(G135), .A2(n913), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G111), .A2(n909), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n910), .A2(G123), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT18), .B(n567), .Z(n568) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n915), .A2(G99), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n935) );
  XNOR2_X1 U639 ( .A(G2096), .B(n935), .ZN(n572) );
  OR2_X1 U640 ( .A1(G2100), .A2(n572), .ZN(G156) );
  INV_X1 U641 ( .A(G132), .ZN(G219) );
  INV_X1 U642 ( .A(G82), .ZN(G220) );
  INV_X1 U643 ( .A(G120), .ZN(G236) );
  INV_X1 U644 ( .A(G69), .ZN(G235) );
  INV_X1 U645 ( .A(G108), .ZN(G238) );
  NAND2_X1 U646 ( .A1(n667), .A2(G52), .ZN(n573) );
  XNOR2_X1 U647 ( .A(KEYINPUT67), .B(n573), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G90), .A2(n662), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G77), .A2(n661), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U651 ( .A(n576), .B(KEYINPUT68), .ZN(n577) );
  XNOR2_X1 U652 ( .A(n577), .B(KEYINPUT9), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n666), .A2(G64), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U655 ( .A1(n581), .A2(n580), .ZN(G171) );
  NAND2_X1 U656 ( .A1(n662), .A2(G89), .ZN(n582) );
  XNOR2_X1 U657 ( .A(n582), .B(KEYINPUT4), .ZN(n584) );
  NAND2_X1 U658 ( .A1(G76), .A2(n661), .ZN(n583) );
  NAND2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U660 ( .A(n585), .B(KEYINPUT5), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n667), .A2(G51), .ZN(n586) );
  XNOR2_X1 U662 ( .A(n586), .B(KEYINPUT78), .ZN(n588) );
  NAND2_X1 U663 ( .A1(G63), .A2(n666), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U665 ( .A(KEYINPUT6), .B(n589), .Z(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U668 ( .A(G168), .B(KEYINPUT8), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT79), .ZN(G286) );
  NAND2_X1 U670 ( .A1(G94), .A2(G452), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n594), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U672 ( .A1(G7), .A2(G661), .ZN(n595) );
  XNOR2_X1 U673 ( .A(n595), .B(KEYINPUT72), .ZN(n596) );
  XNOR2_X1 U674 ( .A(KEYINPUT10), .B(n596), .ZN(G223) );
  INV_X1 U675 ( .A(G223), .ZN(n850) );
  NAND2_X1 U676 ( .A1(n850), .A2(G567), .ZN(n597) );
  XOR2_X1 U677 ( .A(KEYINPUT11), .B(n597), .Z(G234) );
  NAND2_X1 U678 ( .A1(G56), .A2(n666), .ZN(n598) );
  XOR2_X1 U679 ( .A(KEYINPUT14), .B(n598), .Z(n607) );
  NAND2_X1 U680 ( .A1(G81), .A2(n662), .ZN(n601) );
  XOR2_X1 U681 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n599) );
  NAND2_X1 U682 ( .A1(n661), .A2(G68), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n605) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n667), .A2(G43), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n986) );
  INV_X1 U687 ( .A(G860), .ZN(n639) );
  OR2_X1 U688 ( .A1(n986), .A2(n639), .ZN(G153) );
  INV_X1 U689 ( .A(G171), .ZN(G301) );
  NAND2_X1 U690 ( .A1(G868), .A2(G301), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n661), .A2(G79), .ZN(n610) );
  XOR2_X1 U692 ( .A(KEYINPUT75), .B(n610), .Z(n612) );
  NAND2_X1 U693 ( .A1(n667), .A2(G54), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT76), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G66), .A2(n666), .ZN(n615) );
  NAND2_X1 U697 ( .A1(G92), .A2(n662), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n620) );
  BUF_X1 U700 ( .A(n714), .Z(n999) );
  INV_X1 U701 ( .A(G868), .ZN(n681) );
  NAND2_X1 U702 ( .A1(n999), .A2(n681), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(G284) );
  NAND2_X1 U704 ( .A1(G91), .A2(n662), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G78), .A2(n661), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G53), .A2(n667), .ZN(n625) );
  XNOR2_X1 U708 ( .A(n625), .B(KEYINPUT70), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n666), .A2(G65), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n989) );
  XNOR2_X1 U712 ( .A(n989), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U713 ( .A1(G286), .A2(G868), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G299), .A2(n681), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(G297) );
  NAND2_X1 U716 ( .A1(n639), .A2(G559), .ZN(n632) );
  INV_X1 U717 ( .A(n999), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n632), .A2(n637), .ZN(n633) );
  XNOR2_X1 U719 ( .A(n633), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U720 ( .A1(G868), .A2(n986), .ZN(n636) );
  NAND2_X1 U721 ( .A1(G868), .A2(n637), .ZN(n634) );
  NOR2_X1 U722 ( .A1(G559), .A2(n634), .ZN(n635) );
  NOR2_X1 U723 ( .A1(n636), .A2(n635), .ZN(G282) );
  NAND2_X1 U724 ( .A1(G559), .A2(n637), .ZN(n638) );
  XOR2_X1 U725 ( .A(n986), .B(n638), .Z(n678) );
  NAND2_X1 U726 ( .A1(n639), .A2(n678), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G80), .A2(n661), .ZN(n640) );
  XNOR2_X1 U728 ( .A(n640), .B(KEYINPUT80), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n666), .A2(G67), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U731 ( .A1(G93), .A2(n662), .ZN(n644) );
  NAND2_X1 U732 ( .A1(G55), .A2(n667), .ZN(n643) );
  NAND2_X1 U733 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U734 ( .A1(n646), .A2(n645), .ZN(n680) );
  XOR2_X1 U735 ( .A(n647), .B(n680), .Z(G145) );
  NAND2_X1 U736 ( .A1(G61), .A2(n666), .ZN(n649) );
  NAND2_X1 U737 ( .A1(G86), .A2(n662), .ZN(n648) );
  NAND2_X1 U738 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U739 ( .A1(n661), .A2(G73), .ZN(n650) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(n650), .Z(n651) );
  NOR2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U742 ( .A1(n667), .A2(G48), .ZN(n653) );
  NAND2_X1 U743 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U744 ( .A1(G49), .A2(n667), .ZN(n656) );
  NAND2_X1 U745 ( .A1(G74), .A2(G651), .ZN(n655) );
  NAND2_X1 U746 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U747 ( .A1(n666), .A2(n657), .ZN(n660) );
  NAND2_X1 U748 ( .A1(n658), .A2(G87), .ZN(n659) );
  NAND2_X1 U749 ( .A1(n660), .A2(n659), .ZN(G288) );
  NAND2_X1 U750 ( .A1(n661), .A2(G75), .ZN(n665) );
  NAND2_X1 U751 ( .A1(G88), .A2(n662), .ZN(n663) );
  XOR2_X1 U752 ( .A(KEYINPUT81), .B(n663), .Z(n664) );
  NAND2_X1 U753 ( .A1(n665), .A2(n664), .ZN(n671) );
  NAND2_X1 U754 ( .A1(G62), .A2(n666), .ZN(n669) );
  NAND2_X1 U755 ( .A1(G50), .A2(n667), .ZN(n668) );
  NAND2_X1 U756 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U757 ( .A1(n671), .A2(n670), .ZN(G166) );
  INV_X1 U758 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U759 ( .A(n680), .B(G305), .ZN(n672) );
  XNOR2_X1 U760 ( .A(n672), .B(G299), .ZN(n673) );
  XNOR2_X1 U761 ( .A(KEYINPUT82), .B(n673), .ZN(n675) );
  XNOR2_X1 U762 ( .A(G288), .B(KEYINPUT19), .ZN(n674) );
  XNOR2_X1 U763 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U764 ( .A(n676), .B(G290), .ZN(n677) );
  XNOR2_X1 U765 ( .A(n677), .B(G303), .ZN(n857) );
  XOR2_X1 U766 ( .A(n857), .B(n678), .Z(n679) );
  NOR2_X1 U767 ( .A1(n681), .A2(n679), .ZN(n683) );
  AND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U769 ( .A1(n683), .A2(n682), .ZN(G295) );
  NAND2_X1 U770 ( .A1(G2078), .A2(G2084), .ZN(n684) );
  XOR2_X1 U771 ( .A(KEYINPUT20), .B(n684), .Z(n685) );
  NAND2_X1 U772 ( .A1(G2090), .A2(n685), .ZN(n686) );
  XNOR2_X1 U773 ( .A(KEYINPUT21), .B(n686), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n687), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U775 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U776 ( .A1(G235), .A2(G236), .ZN(n688) );
  XNOR2_X1 U777 ( .A(n688), .B(KEYINPUT83), .ZN(n689) );
  NOR2_X1 U778 ( .A1(G238), .A2(n689), .ZN(n690) );
  NAND2_X1 U779 ( .A1(G57), .A2(n690), .ZN(n854) );
  NAND2_X1 U780 ( .A1(G567), .A2(n854), .ZN(n695) );
  NOR2_X1 U781 ( .A1(G220), .A2(G219), .ZN(n691) );
  XOR2_X1 U782 ( .A(KEYINPUT22), .B(n691), .Z(n692) );
  NOR2_X1 U783 ( .A1(G218), .A2(n692), .ZN(n693) );
  NAND2_X1 U784 ( .A1(G96), .A2(n693), .ZN(n855) );
  NAND2_X1 U785 ( .A1(G2106), .A2(n855), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n856) );
  NAND2_X1 U787 ( .A1(G483), .A2(G661), .ZN(n696) );
  NOR2_X1 U788 ( .A1(n856), .A2(n696), .ZN(n853) );
  NAND2_X1 U789 ( .A1(n853), .A2(G36), .ZN(G176) );
  NAND2_X1 U790 ( .A1(G160), .A2(G40), .ZN(n805) );
  INV_X1 U791 ( .A(n805), .ZN(n697) );
  NOR2_X2 U792 ( .A1(G164), .A2(G1384), .ZN(n804) );
  NAND2_X1 U793 ( .A1(n706), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U794 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U795 ( .A1(G1956), .A2(n746), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n703) );
  XNOR2_X1 U797 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n704) );
  XNOR2_X1 U798 ( .A(n705), .B(n704), .ZN(n723) );
  NAND2_X1 U799 ( .A1(G1348), .A2(n746), .ZN(n708) );
  BUF_X2 U800 ( .A(n706), .Z(n726) );
  NAND2_X1 U801 ( .A1(G2067), .A2(n726), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n999), .A2(n713), .ZN(n718) );
  XNOR2_X1 U804 ( .A(G1996), .B(KEYINPUT100), .ZN(n963) );
  NAND2_X1 U805 ( .A1(n963), .A2(n726), .ZN(n709) );
  XNOR2_X1 U806 ( .A(n709), .B(KEYINPUT26), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n746), .A2(G1341), .ZN(n710) );
  NAND2_X1 U808 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U809 ( .A1(n986), .A2(n712), .ZN(n716) );
  NOR2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X2 U811 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n989), .A2(n719), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U816 ( .A(n724), .B(KEYINPUT29), .ZN(n731) );
  XOR2_X1 U817 ( .A(KEYINPUT25), .B(G2078), .Z(n964) );
  NOR2_X1 U818 ( .A1(n964), .A2(n746), .ZN(n725) );
  XOR2_X1 U819 ( .A(KEYINPUT97), .B(n725), .Z(n729) );
  XOR2_X1 U820 ( .A(G1961), .B(KEYINPUT95), .Z(n1019) );
  NOR2_X1 U821 ( .A1(n726), .A2(n1019), .ZN(n727) );
  XNOR2_X1 U822 ( .A(KEYINPUT96), .B(n727), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n739) );
  NOR2_X1 U824 ( .A1(G301), .A2(n739), .ZN(n730) );
  NOR2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n733) );
  XNOR2_X1 U826 ( .A(n733), .B(n732), .ZN(n744) );
  NAND2_X1 U827 ( .A1(G8), .A2(n734), .ZN(n791) );
  NOR2_X1 U828 ( .A1(G1966), .A2(n791), .ZN(n757) );
  NOR2_X1 U829 ( .A1(G2084), .A2(n746), .ZN(n756) );
  NOR2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n735) );
  NAND2_X1 U831 ( .A1(G8), .A2(n735), .ZN(n736) );
  XNOR2_X1 U832 ( .A(KEYINPUT30), .B(n736), .ZN(n737) );
  NOR2_X1 U833 ( .A1(G168), .A2(n737), .ZN(n738) );
  XNOR2_X1 U834 ( .A(n738), .B(KEYINPUT102), .ZN(n741) );
  AND2_X1 U835 ( .A1(n739), .A2(G301), .ZN(n740) );
  NOR2_X1 U836 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U837 ( .A(KEYINPUT31), .B(n742), .ZN(n743) );
  NOR2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U839 ( .A(n745), .B(KEYINPUT103), .ZN(n758) );
  NAND2_X1 U840 ( .A1(n758), .A2(G286), .ZN(n753) );
  INV_X1 U841 ( .A(G8), .ZN(n751) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n791), .ZN(n748) );
  NOR2_X1 U843 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U844 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U845 ( .A1(n749), .A2(G303), .ZN(n750) );
  OR2_X1 U846 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X2 U847 ( .A(n755), .B(n754), .ZN(n776) );
  NAND2_X1 U848 ( .A1(G8), .A2(n756), .ZN(n761) );
  INV_X1 U849 ( .A(n757), .ZN(n759) );
  AND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n774) );
  AND2_X1 U852 ( .A1(n774), .A2(n791), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n776), .A2(n762), .ZN(n766) );
  INV_X1 U854 ( .A(n791), .ZN(n767) );
  NOR2_X1 U855 ( .A1(G2090), .A2(G303), .ZN(n763) );
  NAND2_X1 U856 ( .A1(G8), .A2(n763), .ZN(n764) );
  OR2_X1 U857 ( .A1(n767), .A2(n764), .ZN(n765) );
  AND2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n786) );
  NAND2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n988) );
  AND2_X1 U860 ( .A1(n767), .A2(n988), .ZN(n768) );
  NOR2_X1 U861 ( .A1(KEYINPUT33), .A2(n768), .ZN(n773) );
  XOR2_X1 U862 ( .A(G1981), .B(G305), .Z(n983) );
  INV_X1 U863 ( .A(n983), .ZN(n771) );
  NOR2_X1 U864 ( .A1(G1976), .A2(G288), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n779), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U866 ( .A1(n791), .A2(n769), .ZN(n770) );
  OR2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n777) );
  AND2_X1 U869 ( .A1(n774), .A2(n777), .ZN(n775) );
  NAND2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n784) );
  INV_X1 U871 ( .A(n777), .ZN(n782) );
  NOR2_X1 U872 ( .A1(G1971), .A2(G303), .ZN(n778) );
  NOR2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n990) );
  INV_X1 U874 ( .A(KEYINPUT33), .ZN(n780) );
  AND2_X1 U875 ( .A1(n990), .A2(n780), .ZN(n781) );
  OR2_X1 U876 ( .A1(n782), .A2(n781), .ZN(n783) );
  AND2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U879 ( .A(n787), .B(KEYINPUT105), .ZN(n792) );
  NOR2_X1 U880 ( .A1(G1981), .A2(G305), .ZN(n788) );
  XOR2_X1 U881 ( .A(n788), .B(KEYINPUT24), .Z(n789) );
  XNOR2_X1 U882 ( .A(KEYINPUT94), .B(n789), .ZN(n790) );
  AND2_X1 U883 ( .A1(n792), .A2(n523), .ZN(n827) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n843) );
  XNOR2_X1 U885 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G116), .A2(n909), .ZN(n794) );
  NAND2_X1 U887 ( .A1(G128), .A2(n910), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U889 ( .A(n796), .B(n795), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n915), .A2(G104), .ZN(n797) );
  XNOR2_X1 U891 ( .A(n797), .B(KEYINPUT88), .ZN(n799) );
  NAND2_X1 U892 ( .A1(G140), .A2(n913), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U894 ( .A(KEYINPUT34), .B(n800), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U896 ( .A(KEYINPUT36), .B(n803), .ZN(n923) );
  NOR2_X1 U897 ( .A1(n843), .A2(n923), .ZN(n944) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U899 ( .A(n806), .B(KEYINPUT86), .ZN(n845) );
  NAND2_X1 U900 ( .A1(n944), .A2(n845), .ZN(n807) );
  XNOR2_X1 U901 ( .A(KEYINPUT90), .B(n807), .ZN(n841) );
  NAND2_X1 U902 ( .A1(G105), .A2(n915), .ZN(n808) );
  XNOR2_X1 U903 ( .A(n808), .B(KEYINPUT38), .ZN(n815) );
  NAND2_X1 U904 ( .A1(G141), .A2(n913), .ZN(n810) );
  NAND2_X1 U905 ( .A1(G117), .A2(n909), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n910), .A2(G129), .ZN(n811) );
  XOR2_X1 U908 ( .A(KEYINPUT92), .B(n811), .Z(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n905) );
  NAND2_X1 U911 ( .A1(G1996), .A2(n905), .ZN(n816) );
  XOR2_X1 U912 ( .A(KEYINPUT93), .B(n816), .Z(n825) );
  NAND2_X1 U913 ( .A1(G131), .A2(n913), .ZN(n818) );
  NAND2_X1 U914 ( .A1(G107), .A2(n909), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n821) );
  NAND2_X1 U916 ( .A1(G95), .A2(n915), .ZN(n819) );
  XNOR2_X1 U917 ( .A(KEYINPUT91), .B(n819), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n910), .A2(G119), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n891) );
  NAND2_X1 U921 ( .A1(G1991), .A2(n891), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n943) );
  NAND2_X1 U923 ( .A1(n845), .A2(n943), .ZN(n835) );
  NAND2_X1 U924 ( .A1(n841), .A2(n835), .ZN(n826) );
  NOR2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n829) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n833) );
  INV_X1 U927 ( .A(n845), .ZN(n830) );
  XOR2_X1 U928 ( .A(G1986), .B(G290), .Z(n995) );
  NOR2_X1 U929 ( .A1(n830), .A2(n995), .ZN(n831) );
  XOR2_X1 U930 ( .A(KEYINPUT87), .B(n831), .Z(n832) );
  NOR2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n834), .B(KEYINPUT107), .ZN(n848) );
  NOR2_X1 U933 ( .A1(G1996), .A2(n905), .ZN(n938) );
  INV_X1 U934 ( .A(n835), .ZN(n838) );
  NOR2_X1 U935 ( .A1(G1986), .A2(G290), .ZN(n836) );
  NOR2_X1 U936 ( .A1(G1991), .A2(n891), .ZN(n934) );
  NOR2_X1 U937 ( .A1(n836), .A2(n934), .ZN(n837) );
  NOR2_X1 U938 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U939 ( .A1(n938), .A2(n839), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n840), .B(KEYINPUT39), .ZN(n842) );
  NAND2_X1 U941 ( .A1(n842), .A2(n841), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n843), .A2(n923), .ZN(n948) );
  NAND2_X1 U943 ( .A1(n844), .A2(n948), .ZN(n846) );
  NAND2_X1 U944 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U947 ( .A1(G2106), .A2(n850), .ZN(G217) );
  AND2_X1 U948 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U949 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U950 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(G188) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  NOR2_X1 U954 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U955 ( .A(G325), .ZN(G261) );
  XOR2_X1 U956 ( .A(KEYINPUT108), .B(n856), .Z(G319) );
  XNOR2_X1 U957 ( .A(n986), .B(n857), .ZN(n859) );
  XNOR2_X1 U958 ( .A(G286), .B(G171), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(n999), .ZN(n861) );
  NOR2_X1 U961 ( .A1(G37), .A2(n861), .ZN(G397) );
  XOR2_X1 U962 ( .A(KEYINPUT41), .B(G1981), .Z(n863) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(n864), .B(KEYINPUT113), .Z(n866) );
  XNOR2_X1 U966 ( .A(G1956), .B(G1976), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U968 ( .A(G1966), .B(G1961), .Z(n868) );
  XNOR2_X1 U969 ( .A(G1986), .B(G1971), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U971 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U972 ( .A(G2474), .B(KEYINPUT112), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(G229) );
  XNOR2_X1 U974 ( .A(G2067), .B(G2078), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n873), .B(KEYINPUT42), .ZN(n883) );
  XOR2_X1 U976 ( .A(KEYINPUT111), .B(G2678), .Z(n875) );
  XNOR2_X1 U977 ( .A(KEYINPUT110), .B(G2096), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U979 ( .A(G2100), .B(G2084), .Z(n877) );
  XNOR2_X1 U980 ( .A(G2090), .B(G2072), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U982 ( .A(n879), .B(n878), .Z(n881) );
  XNOR2_X1 U983 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n880) );
  XNOR2_X1 U984 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(G227) );
  NAND2_X1 U986 ( .A1(G124), .A2(n910), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n884), .B(KEYINPUT44), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n909), .A2(G112), .ZN(n885) );
  NAND2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G100), .A2(n915), .ZN(n888) );
  NAND2_X1 U991 ( .A1(G136), .A2(n913), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U993 ( .A1(n890), .A2(n889), .ZN(G162) );
  XNOR2_X1 U994 ( .A(G164), .B(n891), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n892), .B(n935), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n894) );
  XNOR2_X1 U997 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n893) );
  XNOR2_X1 U998 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U999 ( .A(n896), .B(n895), .Z(n908) );
  NAND2_X1 U1000 ( .A1(G103), .A2(n915), .ZN(n898) );
  NAND2_X1 U1001 ( .A1(G139), .A2(n913), .ZN(n897) );
  NAND2_X1 U1002 ( .A1(n898), .A2(n897), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(G115), .A2(n909), .ZN(n900) );
  NAND2_X1 U1004 ( .A1(G127), .A2(n910), .ZN(n899) );
  NAND2_X1 U1005 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1006 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U1007 ( .A1(n903), .A2(n902), .ZN(n950) );
  XOR2_X1 U1008 ( .A(G160), .B(n950), .Z(n904) );
  XNOR2_X1 U1009 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1010 ( .A(G162), .B(n906), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(n908), .B(n907), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(G118), .A2(n909), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(G130), .A2(n910), .ZN(n911) );
  NAND2_X1 U1014 ( .A1(n912), .A2(n911), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(n913), .A2(G142), .ZN(n914) );
  XNOR2_X1 U1016 ( .A(n914), .B(KEYINPUT114), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(G106), .A2(n915), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1019 ( .A(n918), .B(KEYINPUT45), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(n922), .B(n921), .Z(n924) );
  XNOR2_X1 U1022 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n925), .ZN(G395) );
  INV_X1 U1024 ( .A(G319), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n926), .A2(G401), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(G229), .A2(G227), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(G397), .A2(n928), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n931), .A2(G395), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(KEYINPUT117), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1034 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1041) );
  XOR2_X1 U1035 ( .A(G160), .B(G2084), .Z(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1040 ( .A(KEYINPUT118), .B(n939), .Z(n940) );
  XOR2_X1 U1041 ( .A(KEYINPUT51), .B(n940), .Z(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(n947), .B(KEYINPUT119), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n955) );
  XOR2_X1 U1047 ( .A(G2072), .B(n950), .Z(n952) );
  XOR2_X1 U1048 ( .A(G164), .B(G2078), .Z(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1050 ( .A(KEYINPUT50), .B(n953), .Z(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT52), .B(n956), .ZN(n958) );
  INV_X1 U1053 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n959), .A2(G29), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT120), .B(n960), .ZN(n1039) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(G2072), .B(G33), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n963), .B(G32), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G27), .B(n964), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n972) );
  XOR2_X1 U1064 ( .A(G1991), .B(G25), .Z(n969) );
  NAND2_X1 U1065 ( .A1(n969), .A2(G28), .ZN(n970) );
  XOR2_X1 U1066 ( .A(KEYINPUT121), .B(n970), .Z(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1068 ( .A(KEYINPUT53), .B(n973), .Z(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT54), .B(G34), .Z(n974) );
  XNOR2_X1 U1070 ( .A(G2084), .B(n974), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G35), .B(G2090), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1074 ( .A(KEYINPUT55), .B(n979), .Z(n980) );
  NOR2_X1 U1075 ( .A1(G29), .A2(n980), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT122), .B(n981), .Z(n982) );
  NAND2_X1 U1077 ( .A1(G11), .A2(n982), .ZN(n1037) );
  XNOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .ZN(n1009) );
  XNOR2_X1 U1079 ( .A(G168), .B(G1966), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(n985), .B(KEYINPUT57), .ZN(n1007) );
  XNOR2_X1 U1082 ( .A(n986), .B(G1341), .ZN(n1005) );
  XNOR2_X1 U1083 ( .A(G171), .B(G1961), .ZN(n998) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n987) );
  NAND2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n989), .B(G1956), .ZN(n991) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1090 ( .A(KEYINPUT124), .B(n996), .Z(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XOR2_X1 U1092 ( .A(G1348), .B(n999), .Z(n1000) );
  XNOR2_X1 U1093 ( .A(KEYINPUT123), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(KEYINPUT125), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1035) );
  INV_X1 U1099 ( .A(G16), .ZN(n1033) );
  XOR2_X1 U1100 ( .A(G1341), .B(G19), .Z(n1013) );
  XNOR2_X1 U1101 ( .A(G1981), .B(G6), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(G20), .B(G1956), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1105 ( .A(KEYINPUT126), .B(n1014), .ZN(n1017) );
  XOR2_X1 U1106 ( .A(KEYINPUT59), .B(G1348), .Z(n1015) );
  XNOR2_X1 U1107 ( .A(G4), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1109 ( .A(KEYINPUT60), .B(n1018), .ZN(n1028) );
  XNOR2_X1 U1110 ( .A(n1019), .B(G5), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(G1971), .B(G22), .ZN(n1021) );
  XNOR2_X1 U1112 ( .A(G23), .B(G1976), .ZN(n1020) );
  NOR2_X1 U1113 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XOR2_X1 U1114 ( .A(G1986), .B(G24), .Z(n1022) );
  NAND2_X1 U1115 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1116 ( .A(KEYINPUT58), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1117 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1118 ( .A1(n1028), .A2(n1027), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(G21), .B(G1966), .ZN(n1029) );
  NOR2_X1 U1120 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1122 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1123 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1124 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1125 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1126 ( .A(n1041), .B(n1040), .ZN(G311) );
  INV_X1 U1127 ( .A(G311), .ZN(G150) );
endmodule

