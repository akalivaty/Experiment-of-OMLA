//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NAND2_X1  g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT83), .ZN(new_n207));
  NOR4_X1   g006(.A1(new_n207), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT83), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n206), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n206), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n210), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n207), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n209), .A2(KEYINPUT83), .A3(new_n210), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT84), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n203), .B1(new_n214), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT15), .B1(new_n202), .B2(KEYINPUT85), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n204), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n218), .A2(KEYINPUT86), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT86), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n227), .A3(new_n210), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n215), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n202), .A2(KEYINPUT85), .A3(KEYINPUT15), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n225), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n233), .A2(G1gat), .ZN(new_n234));
  INV_X1    g033(.A(G8gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT16), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n236), .B2(G1gat), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n235), .B1(new_n234), .B2(new_n237), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n203), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n204), .B1(new_n221), .B2(KEYINPUT84), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n212), .A2(new_n213), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OR3_X1    g044(.A1(new_n225), .A2(new_n229), .A3(new_n230), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n240), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT13), .Z(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n249), .A2(new_n251), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT17), .B1(new_n223), .B2(new_n231), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT17), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n245), .A2(new_n257), .A3(new_n246), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT87), .B1(new_n259), .B2(new_n240), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT87), .ZN(new_n261));
  AOI211_X1 g060(.A(new_n261), .B(new_n248), .C1(new_n256), .C2(new_n258), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n255), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT18), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT88), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n223), .A2(new_n231), .A3(KEYINPUT17), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n257), .B1(new_n245), .B2(new_n246), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n240), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n261), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n259), .A2(KEYINPUT87), .A3(new_n240), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n249), .A2(KEYINPUT18), .A3(new_n251), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n266), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI211_X1 g074(.A(KEYINPUT88), .B(new_n273), .C1(new_n270), .C2(new_n271), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n265), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G141gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(G197gat), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT11), .B(G169gat), .Z(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT12), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n274), .B1(new_n260), .B2(new_n262), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT88), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n272), .A2(new_n266), .A3(new_n274), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n253), .A2(new_n282), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n263), .B2(new_n264), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n277), .A2(new_n283), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n291));
  XNOR2_X1  g090(.A(G1gat), .B(G29gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT0), .ZN(new_n293));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n296), .B(new_n299), .C1(new_n300), .C2(KEYINPUT2), .ZN(new_n301));
  INV_X1    g100(.A(G141gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G148gat), .ZN(new_n303));
  INV_X1    g102(.A(G148gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G141gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n299), .A2(new_n296), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G134gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G127gat), .ZN(new_n312));
  INV_X1    g111(.A(G127gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G134gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(KEYINPUT1), .ZN(new_n317));
  INV_X1    g116(.A(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G113gat), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G120gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n301), .A2(new_n317), .A3(new_n309), .A4(new_n325), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT73), .B(KEYINPUT5), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n327), .B2(new_n328), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT5), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n328), .A2(KEYINPUT4), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT71), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT72), .B1(new_n328), .B2(KEYINPUT4), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n301), .A2(new_n309), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n317), .A2(new_n325), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT71), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n345), .A3(KEYINPUT4), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n338), .A2(new_n339), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n330), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n341), .B1(KEYINPUT3), .B2(new_n310), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n301), .A2(new_n350), .A3(new_n309), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n343), .A3(new_n341), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n357), .B(new_n355), .C1(new_n328), .C2(KEYINPUT4), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n337), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n328), .B2(KEYINPUT4), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT75), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n328), .A4(new_n359), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT5), .B(new_n348), .C1(new_n349), .C2(new_n351), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI211_X1 g165(.A(new_n291), .B(new_n295), .C1(new_n354), .C2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G211gat), .B(G218gat), .Z(new_n371));
  AOI21_X1  g170(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n372));
  AND2_X1   g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(G197gat), .A2(G204gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n371), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n372), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n377), .B(new_n378), .C1(new_n374), .C2(new_n373), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n379), .A3(KEYINPUT68), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT68), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n371), .B(new_n381), .C1(new_n372), .C2(new_n375), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n388));
  NOR4_X1   g187(.A1(KEYINPUT64), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT64), .ZN(new_n390));
  NOR2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT26), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n387), .B(new_n388), .C1(new_n389), .C2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395));
  INV_X1    g194(.A(G183gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT27), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G183gat), .ZN(new_n399));
  INV_X1    g198(.A(G190gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n395), .B1(new_n401), .B2(KEYINPUT28), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n397), .A2(new_n399), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n400), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G183gat), .A2(G190gat), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n387), .B1(new_n407), .B2(KEYINPUT24), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n400), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(KEYINPUT24), .A3(new_n407), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT25), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n409), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT24), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n395), .A2(new_n417), .B1(G169gat), .B2(G176gat), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n416), .A2(new_n418), .A3(new_n414), .A4(KEYINPUT25), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n406), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n386), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n416), .A2(new_n418), .A3(new_n414), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT25), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n419), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n385), .B1(new_n427), .B2(new_n406), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n384), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n386), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n427), .B2(new_n406), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n430), .B(new_n383), .C1(new_n386), .C2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(KEYINPUT37), .A3(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G8gat), .B(G36gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT69), .ZN(new_n435));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT37), .B1(new_n429), .B2(new_n432), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n438), .A2(KEYINPUT38), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n429), .B2(new_n432), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n354), .A2(new_n366), .ZN(new_n443));
  INV_X1    g242(.A(new_n295), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT6), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n354), .A2(new_n366), .A3(new_n295), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n367), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n370), .B(new_n442), .C1(new_n447), .C2(new_n369), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n444), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n291), .A3(new_n446), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n368), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT79), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n454), .A2(KEYINPUT80), .A3(new_n370), .A4(new_n442), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n439), .B1(new_n438), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n456), .B2(new_n438), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT38), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n450), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n349), .A2(new_n351), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n361), .A2(new_n461), .A3(new_n364), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n348), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n329), .A2(new_n330), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(KEYINPUT39), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n462), .A2(new_n466), .A3(new_n348), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n295), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT30), .ZN(new_n471));
  AOI211_X1 g270(.A(new_n471), .B(new_n437), .C1(new_n429), .C2(new_n432), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n429), .A2(new_n437), .A3(new_n432), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n441), .A2(KEYINPUT30), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n465), .A2(KEYINPUT40), .A3(new_n295), .A4(new_n467), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n470), .A2(new_n451), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n380), .A2(new_n422), .A3(new_n382), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n350), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n310), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n351), .A2(new_n422), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n383), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT77), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n382), .A2(new_n380), .B1(new_n351), .B2(new_n422), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT77), .ZN(new_n488));
  INV_X1    g287(.A(G228gat), .ZN(new_n489));
  INV_X1    g288(.A(G233gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n482), .A2(new_n486), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G22gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n376), .A2(new_n379), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n422), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n340), .B1(new_n495), .B2(new_n350), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n496), .A2(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n493), .B1(new_n492), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g298(.A(G78gat), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n491), .B1(new_n487), .B2(KEYINPUT77), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n340), .B1(new_n480), .B2(new_n350), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n383), .A2(new_n483), .A3(KEYINPUT77), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n497), .ZN(new_n505));
  OAI21_X1  g304(.A(G22gat), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G78gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n497), .A3(new_n493), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT31), .B(G50gat), .ZN(new_n510));
  INV_X1    g309(.A(G106gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n500), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n500), .B2(new_n509), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n479), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n460), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G43gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(G71gat), .B(G99gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n427), .A2(new_n341), .A3(new_n406), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n341), .B1(new_n427), .B2(new_n406), .ZN(new_n523));
  OAI211_X1 g322(.A(G227gat), .B(G233gat), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G227gat), .A2(G233gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n421), .A2(new_n326), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n427), .A2(new_n341), .A3(new_n406), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT65), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT65), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n524), .A2(new_n533), .A3(KEYINPUT32), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n526), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n524), .B(KEYINPUT32), .C1(new_n525), .C2(new_n521), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT67), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n528), .A2(new_n527), .A3(new_n529), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT34), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT66), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n527), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n541), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n538), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n548));
  AND4_X1   g347(.A1(new_n539), .A2(new_n535), .A3(new_n536), .A4(new_n545), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n547), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n441), .A2(KEYINPUT30), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT70), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n473), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n556), .A2(new_n476), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT70), .B1(new_n472), .B2(new_n474), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n453), .A2(new_n557), .A3(KEYINPUT76), .A4(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT76), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n556), .A3(new_n476), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n447), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n515), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT78), .B1(new_n553), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n512), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n498), .A2(new_n499), .A3(G78gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n507), .B1(new_n506), .B2(new_n508), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n500), .A2(new_n509), .A3(new_n512), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n561), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT76), .B1(new_n571), .B2(new_n453), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n447), .A2(new_n561), .A3(new_n560), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n547), .A2(new_n550), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT36), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n545), .B1(new_n537), .B2(KEYINPUT67), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n549), .B1(new_n577), .B2(new_n540), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n548), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n574), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n518), .A2(new_n564), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n454), .A2(new_n370), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n584), .A2(new_n575), .A3(new_n515), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n559), .A2(new_n562), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT82), .B1(new_n578), .B2(new_n570), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT82), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n575), .A2(new_n589), .A3(new_n515), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n290), .B1(new_n583), .B2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G190gat), .B(G218gat), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT95), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT8), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n603), .A2(new_n606), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT92), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G99gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n511), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n602), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n611), .A2(new_n615), .A3(new_n619), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n612), .A2(KEYINPUT93), .A3(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n259), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT94), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT94), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n259), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n247), .A2(new_n626), .B1(KEYINPUT41), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n599), .B(new_n601), .C1(new_n632), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n596), .A2(new_n597), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(KEYINPUT41), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT91), .Z(new_n640));
  XOR2_X1   g439(.A(new_n638), .B(new_n640), .Z(new_n641));
  AOI21_X1  g440(.A(new_n636), .B1(new_n629), .B2(new_n631), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n600), .B1(new_n642), .B2(new_n598), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n637), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n637), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G57gat), .B(G64gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G71gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n507), .ZN(new_n650));
  NAND2_X1  g449(.A1(G71gat), .A2(G78gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT9), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n648), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n651), .B(new_n650), .C1(new_n647), .C2(new_n653), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT21), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT89), .ZN(new_n660));
  XOR2_X1   g459(.A(G127gat), .B(G155gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT20), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G183gat), .B(G211gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n240), .B1(new_n658), .B2(new_n657), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n667));
  NAND2_X1  g466(.A1(G231gat), .A2(G233gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n666), .B(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n665), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT99), .Z(new_n675));
  XOR2_X1   g474(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n611), .B1(new_n615), .B2(new_n619), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n623), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n611), .A2(KEYINPUT97), .A3(new_n615), .A4(new_n619), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n657), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n657), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n624), .B2(new_n625), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n677), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n683), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n675), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n675), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n682), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(G120gat), .B(G148gat), .Z(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n693), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n646), .A2(new_n673), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n594), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n453), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(G1gat), .Z(G1324gat));
  INV_X1    g501(.A(new_n700), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n235), .B1(new_n703), .B2(new_n477), .ZN(new_n704));
  INV_X1    g503(.A(new_n477), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT16), .B(G8gat), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n700), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT42), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(KEYINPUT42), .B2(new_n707), .ZN(G1325gat));
  XNOR2_X1  g508(.A(new_n580), .B(KEYINPUT100), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G15gat), .B1(new_n700), .B2(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n578), .A2(G15gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n700), .B2(new_n713), .ZN(G1326gat));
  AND2_X1   g513(.A1(new_n594), .A2(new_n570), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n699), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT43), .B(G22gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n583), .A2(new_n593), .ZN(new_n720));
  INV_X1    g519(.A(new_n645), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n637), .A2(new_n641), .A3(new_n643), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n719), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n590), .A2(new_n588), .ZN(new_n725));
  INV_X1    g524(.A(new_n587), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n592), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n586), .ZN(new_n728));
  INV_X1    g527(.A(new_n459), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n448), .B2(new_n449), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n516), .B1(new_n730), .B2(new_n455), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n574), .A2(new_n580), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n727), .A2(new_n728), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n733), .A2(new_n723), .A3(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n724), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n290), .A2(new_n673), .A3(new_n696), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G29gat), .B1(new_n738), .B2(new_n453), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n720), .A2(new_n723), .A3(new_n737), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n217), .A3(new_n447), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(G1328gat));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n210), .A3(new_n477), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT46), .Z(new_n745));
  OAI21_X1  g544(.A(G36gat), .B1(new_n738), .B2(new_n705), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(G1329gat));
  INV_X1    g546(.A(G43gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n740), .A2(new_n748), .A3(new_n575), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT102), .Z(new_n750));
  OAI21_X1  g549(.A(G43gat), .B1(new_n738), .B2(new_n580), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G43gat), .B1(new_n738), .B2(new_n711), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n754), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g554(.A(G50gat), .B1(new_n738), .B2(new_n515), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT48), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n673), .A2(G50gat), .A3(new_n696), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n715), .A2(new_n723), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n756), .B(new_n760), .C1(new_n757), .C2(KEYINPUT48), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1331gat));
  INV_X1    g563(.A(new_n290), .ZN(new_n765));
  INV_X1    g564(.A(new_n673), .ZN(new_n766));
  NOR4_X1   g565(.A1(new_n723), .A2(new_n765), .A3(new_n766), .A4(new_n697), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n733), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n447), .B(KEYINPUT104), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g570(.A(new_n705), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT105), .Z(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1333gat));
  NAND3_X1  g575(.A1(new_n768), .A2(new_n649), .A3(new_n575), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n768), .A2(new_n710), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n649), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g579(.A1(new_n768), .A2(new_n570), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT106), .B(G78gat), .Z(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n765), .A2(new_n673), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n733), .A2(new_n723), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n723), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(KEYINPUT107), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(KEYINPUT107), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n790), .A2(new_n791), .A3(new_n697), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(new_n607), .A3(new_n447), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n765), .A2(new_n673), .A3(new_n697), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n736), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G85gat), .B1(new_n795), .B2(new_n453), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(G1336gat));
  NAND3_X1  g596(.A1(new_n736), .A2(new_n477), .A3(new_n794), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n786), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n800), .A3(KEYINPUT51), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n697), .A2(new_n705), .A3(G92gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n805), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n807), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n806), .A2(new_n807), .B1(new_n799), .B2(new_n809), .ZN(G1337gat));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n616), .A3(new_n575), .ZN(new_n811));
  OAI21_X1  g610(.A(G99gat), .B1(new_n795), .B2(new_n711), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1338gat));
  OAI211_X1 g612(.A(new_n570), .B(new_n794), .C1(new_n724), .C2(new_n735), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n515), .A2(G106gat), .A3(new_n697), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n802), .A2(new_n803), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT53), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT53), .B1(new_n789), .B2(new_n816), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n815), .A2(new_n820), .A3(KEYINPUT109), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT109), .B1(new_n815), .B2(new_n820), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT110), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n819), .B(new_n825), .C1(new_n821), .C2(new_n822), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(G1339gat));
  INV_X1    g626(.A(new_n249), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n270), .B2(new_n271), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n829), .A2(new_n251), .B1(new_n250), .B2(new_n252), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n287), .A2(new_n289), .B1(new_n830), .B2(new_n281), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n696), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n626), .A2(new_n657), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n679), .B1(new_n612), .B2(new_n620), .ZN(new_n834));
  INV_X1    g633(.A(new_n623), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n681), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n683), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n676), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n686), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n688), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n685), .A2(new_n675), .A3(new_n686), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n693), .B1(new_n687), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT111), .A4(KEYINPUT55), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n695), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT55), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n843), .A2(new_n845), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g653(.A(KEYINPUT112), .B(KEYINPUT55), .C1(new_n843), .C2(new_n845), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n847), .B(new_n850), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n832), .B1(new_n856), .B2(new_n290), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n646), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n850), .A2(new_n695), .A3(new_n846), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n852), .A2(new_n853), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT112), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n852), .A2(new_n851), .A3(new_n853), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n723), .A2(new_n859), .A3(new_n863), .A4(new_n831), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n673), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n698), .A2(new_n765), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n865), .A2(KEYINPUT113), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n289), .B1(new_n275), .B2(new_n276), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n282), .B1(new_n287), .B2(new_n265), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n859), .B(new_n863), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n723), .B1(new_n872), .B2(new_n832), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n251), .B1(new_n272), .B2(new_n249), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n250), .A2(new_n252), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n281), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n646), .A2(new_n856), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n766), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n866), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n867), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n725), .A3(new_n769), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n477), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n765), .A2(new_n320), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT115), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT113), .B1(new_n865), .B2(new_n866), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n879), .A2(new_n880), .A3(new_n868), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n570), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n453), .A2(new_n477), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n575), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n290), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n320), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT114), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n895), .A2(KEYINPUT114), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n887), .B1(new_n897), .B2(new_n898), .ZN(G1340gat));
  AOI21_X1  g698(.A(G120gat), .B1(new_n884), .B2(new_n696), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n893), .A2(new_n318), .A3(new_n697), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(G1341gat));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n313), .A3(new_n673), .ZN(new_n903));
  OAI21_X1  g702(.A(G127gat), .B1(new_n893), .B2(new_n766), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1342gat));
  NOR4_X1   g704(.A1(new_n883), .A2(G134gat), .A3(new_n477), .A4(new_n646), .ZN(new_n906));
  XOR2_X1   g705(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n907));
  OR2_X1    g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G134gat), .B1(new_n893), .B2(new_n646), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(new_n907), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G1343gat));
  NAND2_X1  g710(.A1(new_n580), .A2(new_n892), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n888), .A2(new_n570), .A3(new_n889), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n515), .A2(new_n915), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT117), .B1(new_n831), .B2(new_n696), .ZN(new_n919));
  AND4_X1   g718(.A1(KEYINPUT117), .A2(new_n869), .A3(new_n696), .A4(new_n876), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n847), .A2(new_n850), .A3(new_n860), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n919), .A2(new_n920), .B1(new_n290), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI221_X1 g723(.A(KEYINPUT118), .B1(new_n290), .B2(new_n921), .C1(new_n919), .C2(new_n920), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n646), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n673), .B1(new_n926), .B2(new_n864), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n917), .B(new_n918), .C1(new_n927), .C2(new_n866), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n916), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n723), .B1(new_n922), .B2(new_n923), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n878), .B1(new_n930), .B2(new_n925), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n880), .B1(new_n931), .B2(new_n673), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n917), .B1(new_n932), .B2(new_n918), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n765), .B(new_n913), .C1(new_n929), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G141gat), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n710), .A2(new_n515), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n888), .A2(new_n889), .A3(new_n769), .A4(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n290), .A2(G141gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n705), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT58), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n882), .A2(KEYINPUT120), .A3(new_n769), .A4(new_n936), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n943), .A2(new_n705), .A3(new_n939), .A4(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT58), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n935), .A2(new_n948), .A3(KEYINPUT121), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT121), .B1(new_n935), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(G1344gat));
  NAND2_X1  g750(.A1(new_n943), .A2(new_n945), .ZN(new_n952));
  OR4_X1    g751(.A1(G148gat), .A2(new_n952), .A3(new_n477), .A4(new_n697), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n304), .A2(KEYINPUT59), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n929), .A2(new_n933), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n955), .A2(new_n912), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n956), .B2(new_n696), .ZN(new_n957));
  XOR2_X1   g756(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n958));
  NAND2_X1  g757(.A1(new_n932), .A2(new_n570), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n915), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n915), .B2(new_n914), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n696), .A3(new_n913), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n958), .B1(new_n962), .B2(G148gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n953), .B1(new_n957), .B2(new_n963), .ZN(G1345gat));
  NAND2_X1  g763(.A1(new_n673), .A2(G155gat), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT123), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n943), .A2(new_n705), .A3(new_n673), .A4(new_n945), .ZN(new_n967));
  AOI22_X1  g766(.A1(new_n956), .A2(new_n966), .B1(new_n297), .B2(new_n967), .ZN(G1346gat));
  NOR3_X1   g767(.A1(new_n955), .A2(new_n646), .A3(new_n912), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n723), .A2(new_n298), .A3(new_n705), .ZN(new_n970));
  OAI22_X1  g769(.A1(new_n969), .A2(new_n298), .B1(new_n952), .B2(new_n970), .ZN(G1347gat));
  NOR2_X1   g770(.A1(new_n769), .A2(new_n705), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT125), .Z(new_n973));
  NAND3_X1  g772(.A1(new_n891), .A2(new_n575), .A3(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(G169gat), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n974), .A2(new_n975), .A3(new_n290), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n882), .A2(new_n453), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n705), .B1(new_n977), .B2(KEYINPUT124), .ZN(new_n978));
  OR3_X1    g777(.A1(new_n890), .A2(KEYINPUT124), .A3(new_n447), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n978), .A2(new_n725), .A3(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n765), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n976), .B1(new_n982), .B2(new_n975), .ZN(G1348gat));
  OAI21_X1  g782(.A(G176gat), .B1(new_n974), .B2(new_n697), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n697), .A2(G176gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n980), .B2(new_n985), .ZN(G1349gat));
  OAI21_X1  g785(.A(G183gat), .B1(new_n974), .B2(new_n766), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n673), .A2(new_n403), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g789(.A(G190gat), .B1(new_n974), .B2(new_n646), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT61), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n646), .A2(G190gat), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n993), .B1(new_n981), .B2(new_n994), .ZN(new_n995));
  NOR4_X1   g794(.A1(new_n980), .A2(KEYINPUT126), .A3(G190gat), .A4(new_n646), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G1351gat));
  AND2_X1   g796(.A1(new_n973), .A2(new_n711), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n961), .A2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(G197gat), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n999), .A2(new_n1000), .A3(new_n290), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n978), .A2(new_n979), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1002), .A2(new_n765), .A3(new_n936), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1001), .B1(new_n1000), .B2(new_n1003), .ZN(G1352gat));
  NOR2_X1   g803(.A1(new_n697), .A2(G204gat), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n978), .A2(new_n936), .A3(new_n979), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n961), .A2(new_n696), .A3(new_n998), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(G204gat), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1008), .B1(new_n1012), .B2(new_n1013), .ZN(G1353gat));
  NAND3_X1  g813(.A1(new_n961), .A2(new_n673), .A3(new_n998), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n1015), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT63), .B1(new_n1015), .B2(G211gat), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n936), .ZN(new_n1018));
  OR2_X1    g817(.A1(new_n766), .A2(G211gat), .ZN(new_n1019));
  OAI22_X1  g818(.A1(new_n1016), .A2(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(G1354gat));
  OAI21_X1  g819(.A(G218gat), .B1(new_n999), .B2(new_n646), .ZN(new_n1021));
  OR2_X1    g820(.A1(new_n646), .A2(G218gat), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1021), .B1(new_n1018), .B2(new_n1022), .ZN(G1355gat));
endmodule


