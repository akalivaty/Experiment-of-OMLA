//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT2), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G141gat), .B(G148gat), .Z(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(KEYINPUT75), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n211), .B(KEYINPUT2), .C1(new_n204), .C2(new_n205), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n207), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(new_n202), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT76), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n216), .A3(new_n202), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n209), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT29), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G197gat), .B(G204gat), .ZN(new_n221));
  AND2_X1   g020(.A1(G211gat), .A2(G218gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(KEYINPUT22), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G211gat), .B(G218gat), .Z(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT71), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n226), .A2(new_n227), .B1(new_n228), .B2(new_n224), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n220), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT29), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT3), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(G228gat), .B(G233gat), .C1(new_n232), .C2(new_n218), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n220), .A2(KEYINPUT81), .A3(new_n229), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n218), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n226), .A2(KEYINPUT29), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n223), .A2(new_n225), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n219), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT81), .B1(new_n220), .B2(new_n229), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G228gat), .A2(G233gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n234), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G22gat), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT82), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G78gat), .B(G106gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT80), .B(G50gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n251));
  XOR2_X1   g050(.A(new_n250), .B(new_n251), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n243), .A2(new_n244), .ZN(new_n254));
  INV_X1    g053(.A(new_n234), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n246), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI211_X1 g055(.A(G22gat), .B(new_n234), .C1(new_n243), .C2(new_n244), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n247), .A2(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n255), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G22gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n246), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT82), .A4(new_n252), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G15gat), .B(G43gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G71gat), .B(G99gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT67), .B(G190gat), .Z(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT27), .B(G183gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT26), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT66), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n274), .A2(new_n276), .B1(G183gat), .B2(G190gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT25), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n273), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n276), .ZN(new_n282));
  NOR2_X1   g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT24), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT24), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(G183gat), .A3(G190gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n283), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n279), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n287), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT67), .B(G190gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(G183gat), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n276), .A4(new_n281), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n297));
  AND2_X1   g096(.A1(KEYINPUT68), .A2(G127gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n299), .A2(KEYINPUT69), .ZN(new_n300));
  INV_X1    g099(.A(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G113gat), .ZN(new_n302));
  INV_X1    g101(.A(G113gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G120gat), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT1), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(new_n299), .B2(KEYINPUT69), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n296), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n267), .B1(new_n295), .B2(new_n309), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n272), .A2(new_n277), .B1(new_n289), .B2(new_n293), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n300), .A2(new_n306), .B1(new_n305), .B2(new_n296), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT70), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n309), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G227gat), .A2(G233gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT64), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT65), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT33), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n266), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(KEYINPUT32), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n315), .A2(new_n317), .ZN(new_n324));
  INV_X1    g123(.A(new_n315), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n318), .A2(KEYINPUT34), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n324), .A2(KEYINPUT34), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n319), .B(KEYINPUT32), .C1(new_n320), .C2(new_n266), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n323), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n263), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n295), .A2(new_n231), .ZN(new_n334));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n295), .A2(G226gat), .A3(G233gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n229), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n295), .A2(KEYINPUT72), .A3(G226gat), .A4(G233gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n311), .B2(new_n335), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n339), .A2(new_n341), .B1(new_n334), .B2(new_n335), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n338), .B1(new_n342), .B2(new_n229), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(KEYINPUT73), .ZN(new_n346));
  XOR2_X1   g145(.A(G64gat), .B(G92gat), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(KEYINPUT30), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n338), .B(new_n348), .C1(new_n342), .C2(new_n229), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n348), .B(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n349), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT5), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n312), .A2(new_n218), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT77), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n312), .A2(new_n360), .A3(new_n218), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n237), .A2(new_n309), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n357), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(new_n367), .A3(new_n361), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n218), .A2(new_n219), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n218), .A2(new_n219), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n309), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n358), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT4), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n368), .A2(new_n372), .A3(new_n364), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n367), .B1(new_n359), .B2(new_n361), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n373), .A2(KEYINPUT4), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(new_n309), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n357), .B(new_n364), .C1(new_n380), .C2(new_n369), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT0), .ZN(new_n386));
  XNOR2_X1  g185(.A(G57gat), .B(G85gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT6), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n375), .A2(new_n366), .B1(new_n379), .B2(new_n382), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n388), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(KEYINPUT78), .A3(new_n392), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n391), .A2(new_n397), .A3(new_n388), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n333), .A2(KEYINPUT35), .A3(new_n356), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT35), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n258), .A2(new_n262), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n356), .A3(new_n331), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n398), .B1(new_n392), .B2(new_n390), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n348), .B1(new_n343), .B2(KEYINPUT37), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n339), .A2(new_n341), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n336), .ZN(new_n412));
  INV_X1    g211(.A(new_n229), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n338), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n416), .B1(new_n407), .B2(new_n408), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT38), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT38), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n353), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n336), .A2(new_n337), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n421), .B2(new_n413), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n412), .A2(new_n229), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n424), .A2(new_n416), .B1(new_n344), .B2(new_n348), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n418), .A2(new_n393), .A3(new_n399), .A4(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n363), .A2(new_n365), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT39), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n372), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n430), .A2(new_n377), .A3(new_n378), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n431), .B2(new_n364), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n379), .A2(new_n372), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n428), .A3(new_n365), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n434), .A3(new_n388), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT40), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n384), .A2(new_n389), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n432), .A2(new_n434), .A3(KEYINPUT40), .A4(new_n388), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n355), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n426), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n258), .A2(new_n262), .A3(new_n356), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n441), .A2(new_n403), .B1(new_n400), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n331), .A2(KEYINPUT36), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n329), .B2(new_n330), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n401), .B(new_n406), .C1(new_n443), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n450));
  NAND2_X1  g249(.A1(G229gat), .A2(G233gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT13), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G15gat), .B(G22gat), .ZN(new_n454));
  INV_X1    g253(.A(G1gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT16), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(G1gat), .B2(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G8gat), .ZN(new_n459));
  INV_X1    g258(.A(G8gat), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n457), .B(new_n460), .C1(G1gat), .C2(new_n454), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT88), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT88), .ZN(new_n464));
  NAND2_X1  g263(.A1(G29gat), .A2(G36gat), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NOR3_X1   g266(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(KEYINPUT15), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n472));
  INV_X1    g271(.A(G29gat), .ZN(new_n473));
  INV_X1    g272(.A(G36gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n468), .A2(KEYINPUT86), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n480));
  XOR2_X1   g279(.A(G43gat), .B(G50gat), .Z(new_n481));
  INV_X1    g280(.A(KEYINPUT15), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n479), .A2(new_n465), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n463), .A2(new_n464), .A3(new_n471), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n465), .A3(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n475), .A2(new_n476), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n468), .A2(KEYINPUT86), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n467), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n471), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n464), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n462), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n453), .B1(new_n485), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n484), .A2(KEYINPUT87), .A3(new_n494), .A4(new_n471), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n459), .A3(new_n461), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n451), .A3(new_n492), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n493), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n500), .A2(KEYINPUT18), .A3(new_n451), .A4(new_n492), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n503), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n503), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n450), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n503), .A2(new_n511), .ZN(new_n515));
  INV_X1    g314(.A(new_n510), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n503), .A2(new_n510), .A3(new_n511), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT89), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n449), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n449), .A2(KEYINPUT90), .A3(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n400), .ZN(new_n526));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT8), .ZN(new_n528));
  INV_X1    g327(.A(G85gat), .ZN(new_n529));
  INV_X1    g328(.A(G92gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(KEYINPUT95), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n537));
  NOR2_X1   g336(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n538));
  OAI22_X1  g337(.A1(new_n537), .A2(new_n538), .B1(new_n529), .B2(new_n530), .ZN(new_n539));
  OR2_X1    g338(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n540));
  AND2_X1   g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT96), .ZN(new_n545));
  XOR2_X1   g344(.A(G99gat), .B(G106gat), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n536), .A2(new_n544), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n528), .A2(KEYINPUT95), .A3(new_n531), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT95), .B1(new_n528), .B2(new_n531), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n539), .A2(new_n543), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n547), .A3(new_n544), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(KEYINPUT96), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n499), .A2(new_n548), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n548), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n490), .ZN(new_n558));
  NAND3_X1  g357(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G190gat), .B(G218gat), .Z(new_n561));
  AND2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n567), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G57gat), .B(G64gat), .Z(new_n571));
  NAND2_X1  g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(KEYINPUT9), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(KEYINPUT91), .ZN(new_n575));
  NOR2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT91), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n572), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G57gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G64gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n576), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT9), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n572), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G127gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n587), .ZN(new_n594));
  AOI211_X1 g393(.A(new_n462), .B(new_n491), .C1(KEYINPUT21), .C2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n593), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT93), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G155gat), .ZN(new_n599));
  XOR2_X1   g398(.A(G183gat), .B(G211gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n593), .A2(new_n595), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n593), .A2(new_n595), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n605), .A3(new_n601), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n555), .A2(new_n587), .A3(new_n548), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n553), .A3(new_n554), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT97), .A4(new_n611), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n609), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n608), .B1(new_n610), .B2(new_n612), .ZN(new_n620));
  XOR2_X1   g419(.A(G120gat), .B(G148gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT98), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n608), .B(KEYINPUT99), .Z(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n617), .B2(new_n618), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n625), .B1(new_n630), .B2(new_n620), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n570), .A2(new_n607), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n525), .A2(new_n526), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g434(.A1(new_n449), .A2(KEYINPUT90), .A3(new_n520), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT90), .B1(new_n449), .B2(new_n520), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n355), .B(new_n633), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT100), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n525), .A2(new_n640), .A3(new_n355), .A4(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n641), .A3(G8gat), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT16), .B(G8gat), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT42), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n638), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n633), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n523), .B2(new_n524), .ZN(new_n648));
  INV_X1    g447(.A(new_n645), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n648), .A2(KEYINPUT101), .A3(new_n355), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n644), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n639), .B2(new_n641), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n642), .B(new_n651), .C1(new_n653), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g453(.A(new_n648), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n655), .B2(new_n447), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n332), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n655), .B2(new_n657), .ZN(G1326gat));
  NAND3_X1  g457(.A1(new_n525), .A2(new_n263), .A3(new_n633), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  INV_X1    g460(.A(new_n570), .ZN(new_n662));
  INV_X1    g461(.A(new_n607), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n662), .A2(new_n663), .A3(new_n632), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n525), .A2(new_n473), .A3(new_n526), .A4(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT45), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n449), .A2(new_n570), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n449), .A2(KEYINPUT44), .A3(new_n570), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n607), .B(KEYINPUT102), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n632), .B(KEYINPUT103), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n512), .A2(new_n513), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678), .B2(new_n400), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n665), .A2(new_n666), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n667), .A2(new_n679), .A3(new_n680), .ZN(G1328gat));
  NOR2_X1   g480(.A1(new_n356), .A2(G36gat), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n664), .B(new_n682), .C1(new_n636), .C2(new_n637), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT104), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n525), .A2(new_n685), .A3(new_n664), .A4(new_n682), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G36gat), .B1(new_n678), .B2(new_n356), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n686), .A3(KEYINPUT46), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(G1329gat));
  NAND4_X1  g491(.A1(new_n670), .A2(new_n448), .A3(new_n671), .A4(new_n677), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n332), .A2(G43gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n525), .A2(new_n664), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(new_n694), .B2(new_n696), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(G1330gat));
  NAND4_X1  g499(.A1(new_n670), .A2(new_n263), .A3(new_n671), .A4(new_n677), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G50gat), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT48), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n403), .A2(G50gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n525), .A2(new_n664), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n702), .B(new_n706), .C1(new_n703), .C2(KEYINPUT48), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1331gat));
  NAND4_X1  g509(.A1(new_n675), .A2(new_n676), .A3(new_n663), .A4(new_n662), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n400), .A2(KEYINPUT35), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n404), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n400), .A2(new_n442), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n424), .A2(new_n416), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n350), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n407), .A2(new_n408), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n409), .A3(new_n416), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n718), .B2(KEYINPUT38), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n439), .A2(new_n438), .A3(new_n355), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n719), .A2(new_n405), .B1(new_n720), .B2(new_n437), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n714), .B1(new_n721), .B2(new_n263), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n713), .B1(new_n722), .B2(new_n447), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n711), .B1(new_n723), .B2(new_n406), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n526), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g525(.A(new_n356), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1333gat));
  XNOR2_X1  g529(.A(new_n331), .B(KEYINPUT108), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n724), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(G71gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n724), .A2(G71gat), .A3(new_n448), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(KEYINPUT107), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(KEYINPUT107), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n735), .B(new_n740), .C1(new_n737), .C2(new_n738), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n724), .A2(new_n263), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  INV_X1    g545(.A(new_n676), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n663), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n632), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n672), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n400), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n662), .B1(new_n723), .B2(new_n406), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT51), .B1(new_n754), .B2(new_n748), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n668), .A2(new_n756), .A3(new_n749), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n632), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n526), .A2(new_n529), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n753), .B1(new_n758), .B2(new_n759), .ZN(G1336gat));
  NOR2_X1   g559(.A1(new_n356), .A2(G92gat), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n675), .B(new_n761), .C1(new_n755), .C2(new_n757), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n670), .A2(new_n355), .A3(new_n671), .A4(new_n751), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G92gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n764), .A3(KEYINPUT110), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT52), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n762), .A2(new_n764), .A3(KEYINPUT110), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n752), .B2(new_n447), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n332), .A2(G99gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n758), .B2(new_n771), .ZN(G1338gat));
  NOR2_X1   g571(.A1(new_n403), .A2(G106gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n675), .B(new_n773), .C1(new_n755), .C2(new_n757), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n670), .A2(new_n263), .A3(new_n671), .A4(new_n751), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n617), .A2(new_n618), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n608), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n618), .A2(new_n629), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n615), .B2(new_n616), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n782), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n624), .B1(new_n630), .B2(new_n787), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n627), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n629), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n783), .A2(new_n787), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n625), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n619), .A2(new_n787), .A3(new_n786), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n782), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n791), .A2(new_n796), .A3(new_n747), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n451), .B1(new_n500), .B2(new_n492), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n485), .A2(new_n492), .A3(new_n453), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n508), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n518), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n632), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n570), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  AND4_X1   g603(.A1(new_n570), .A2(new_n802), .A3(new_n791), .A4(new_n796), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n673), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n633), .A2(new_n676), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n806), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n404), .A2(new_n400), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n520), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n813), .A2(new_n303), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n813), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n747), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n303), .B2(new_n817), .ZN(G1340gat));
  OAI21_X1  g617(.A(new_n301), .B1(new_n813), .B2(new_n750), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n675), .A2(G120gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT112), .Z(G1341gat));
  OAI21_X1  g621(.A(G127gat), .B1(new_n813), .B2(new_n673), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n663), .A2(new_n592), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n813), .B2(new_n824), .ZN(G1342gat));
  NAND2_X1  g624(.A1(new_n816), .A2(new_n570), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n826), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT56), .B1(new_n826), .B2(G134gat), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT113), .B1(new_n826), .B2(G134gat), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n826), .A2(KEYINPUT113), .A3(G134gat), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n520), .A2(new_n791), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n784), .A2(new_n788), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n790), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n835));
  XNOR2_X1  g634(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n834), .B2(KEYINPUT114), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n832), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n803), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n662), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n805), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n663), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n676), .B2(new_n633), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT57), .B1(new_n843), .B2(new_n403), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n809), .A2(new_n810), .A3(new_n403), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n448), .A2(new_n355), .A3(new_n400), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G141gat), .B1(new_n849), .B2(new_n814), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n845), .A2(new_n848), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(G141gat), .A3(new_n814), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(KEYINPUT58), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n844), .A2(new_n847), .A3(new_n747), .A4(new_n848), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n852), .B1(new_n856), .B2(G141gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(G1344gat));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(G148gat), .C1(new_n849), .C2(new_n750), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n647), .A2(new_n520), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n846), .B(new_n263), .C1(new_n842), .C2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n848), .A2(new_n632), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n863), .B(new_n864), .C1(new_n845), .C2(new_n846), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G148gat), .ZN(new_n866));
  XOR2_X1   g665(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n861), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  AOI211_X1 g668(.A(KEYINPUT117), .B(new_n867), .C1(new_n865), .C2(G148gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n851), .A2(G148gat), .A3(new_n750), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1345gat));
  NOR3_X1   g672(.A1(new_n849), .A2(new_n204), .A3(new_n673), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n851), .A2(new_n607), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n876));
  AOI21_X1  g675(.A(G155gat), .B1(new_n875), .B2(KEYINPUT118), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(G1346gat));
  NOR3_X1   g677(.A1(new_n849), .A2(new_n205), .A3(new_n662), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n845), .A2(new_n570), .A3(new_n848), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n205), .B2(new_n880), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n333), .A2(new_n355), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n811), .A2(new_n400), .A3(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(G169gat), .A3(new_n676), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT119), .Z(new_n886));
  NAND2_X1  g685(.A1(new_n806), .A2(new_n808), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT111), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n400), .A2(new_n355), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(new_n731), .A3(new_n263), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n888), .A2(new_n889), .A3(new_n891), .A4(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n814), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n886), .A2(new_n897), .ZN(G1348gat));
  INV_X1    g697(.A(new_n675), .ZN(new_n899));
  OAI21_X1  g698(.A(G176gat), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n750), .A2(G176gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n884), .B2(new_n901), .ZN(G1349gat));
  NAND2_X1  g701(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n663), .A2(new_n269), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n884), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n894), .A2(new_n674), .A3(new_n895), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(G183gat), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n907), .B(new_n908), .ZN(G1350gat));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n570), .A3(new_n895), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT123), .B1(new_n911), .B2(G190gat), .ZN(new_n913));
  OAI211_X1 g712(.A(KEYINPUT124), .B(new_n910), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(G190gat), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n911), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n918));
  XNOR2_X1  g717(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n884), .A2(new_n291), .A3(new_n662), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT122), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n920), .A3(new_n922), .ZN(G1351gat));
  AOI21_X1  g722(.A(new_n356), .B1(new_n444), .B2(new_n446), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n263), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT125), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n811), .A2(new_n400), .A3(new_n926), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(G197gat), .A3(new_n676), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n888), .A2(new_n889), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT57), .B1(new_n929), .B2(new_n403), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n448), .A2(new_n890), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n930), .A2(new_n520), .A3(new_n863), .A4(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n928), .B1(new_n932), .B2(G197gat), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT126), .ZN(G1352gat));
  INV_X1    g733(.A(G204gat), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n930), .A2(new_n863), .A3(new_n931), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n675), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n632), .A2(new_n935), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n927), .A2(KEYINPUT62), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT62), .B1(new_n927), .B2(new_n938), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT127), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n930), .A2(new_n863), .A3(new_n931), .ZN(new_n943));
  OAI21_X1  g742(.A(G204gat), .B1(new_n943), .B2(new_n899), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n944), .A2(new_n945), .A3(new_n940), .A4(new_n939), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n942), .A2(new_n946), .ZN(G1353gat));
  OR3_X1    g746(.A1(new_n927), .A2(G211gat), .A3(new_n607), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n930), .A2(new_n663), .A3(new_n863), .A4(new_n931), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n943), .B2(new_n662), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n662), .A2(G218gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n953), .B1(new_n927), .B2(new_n954), .ZN(G1355gat));
endmodule


