

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U548 ( .A1(n777), .A2(n696), .ZN(n737) );
  AND2_X1 U549 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U550 ( .A1(KEYINPUT33), .A2(n763), .ZN(n515) );
  AND2_X1 U551 ( .A1(n742), .A2(n741), .ZN(n516) );
  OR2_X1 U552 ( .A1(KEYINPUT33), .A2(n762), .ZN(n517) );
  OR2_X1 U553 ( .A1(n775), .A2(n774), .ZN(n518) );
  AND2_X1 U554 ( .A1(n931), .A2(n820), .ZN(n519) );
  NAND2_X1 U555 ( .A1(n737), .A2(G1341), .ZN(n520) );
  XOR2_X1 U556 ( .A(n730), .B(KEYINPUT28), .Z(n521) );
  OR2_X1 U557 ( .A1(n737), .A2(n722), .ZN(n723) );
  INV_X1 U558 ( .A(KEYINPUT97), .ZN(n732) );
  XNOR2_X1 U559 ( .A(n732), .B(KEYINPUT29), .ZN(n733) );
  XNOR2_X1 U560 ( .A(n734), .B(n733), .ZN(n746) );
  INV_X1 U561 ( .A(n934), .ZN(n759) );
  NOR2_X1 U562 ( .A1(n756), .A2(n755), .ZN(n767) );
  NOR2_X1 U563 ( .A1(n945), .A2(n515), .ZN(n764) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n777) );
  NOR2_X1 U565 ( .A1(n807), .A2(n519), .ZN(n808) );
  AND2_X1 U566 ( .A1(n526), .A2(G2104), .ZN(n882) );
  XOR2_X1 U567 ( .A(KEYINPUT64), .B(n527), .Z(n878) );
  NOR2_X1 U568 ( .A1(G651), .A2(n653), .ZN(n657) );
  NOR2_X1 U569 ( .A1(n538), .A2(n537), .ZN(G160) );
  XNOR2_X1 U570 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X1 U572 ( .A(n523), .B(n522), .ZN(n881) );
  NAND2_X1 U573 ( .A1(G138), .A2(n881), .ZN(n525) );
  INV_X1 U574 ( .A(G2105), .ZN(n526) );
  NAND2_X1 U575 ( .A1(G102), .A2(n882), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n526), .ZN(n877) );
  NAND2_X1 U578 ( .A1(n877), .A2(G126), .ZN(n529) );
  NAND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  NAND2_X1 U580 ( .A1(G114), .A2(n878), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U582 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U583 ( .A1(n881), .A2(G137), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G101), .A2(n882), .ZN(n532) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n532), .Z(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U587 ( .A1(n877), .A2(G125), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G113), .A2(n878), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n537) );
  INV_X1 U590 ( .A(G651), .ZN(n541) );
  NOR2_X1 U591 ( .A1(G543), .A2(n541), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n539), .Z(n656) );
  NAND2_X1 U593 ( .A1(n656), .A2(G64), .ZN(n540) );
  XNOR2_X1 U594 ( .A(KEYINPUT67), .B(n540), .ZN(n550) );
  XOR2_X1 U595 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  NOR2_X1 U596 ( .A1(n653), .A2(n541), .ZN(n664) );
  NAND2_X1 U597 ( .A1(n664), .A2(G77), .ZN(n542) );
  XNOR2_X1 U598 ( .A(n542), .B(KEYINPUT68), .ZN(n544) );
  NOR2_X1 U599 ( .A1(G651), .A2(G543), .ZN(n660) );
  NAND2_X1 U600 ( .A1(G90), .A2(n660), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U602 ( .A(KEYINPUT69), .B(n545), .Z(n546) );
  XNOR2_X1 U603 ( .A(n546), .B(KEYINPUT9), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G52), .A2(n657), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U607 ( .A(KEYINPUT70), .B(n551), .ZN(G171) );
  INV_X1 U608 ( .A(G171), .ZN(G301) );
  XOR2_X1 U609 ( .A(G2435), .B(G2454), .Z(n553) );
  XNOR2_X1 U610 ( .A(KEYINPUT101), .B(G2438), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n553), .B(n552), .ZN(n560) );
  XOR2_X1 U612 ( .A(G2446), .B(G2430), .Z(n555) );
  XNOR2_X1 U613 ( .A(G2451), .B(G2443), .ZN(n554) );
  XNOR2_X1 U614 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U615 ( .A(n556), .B(G2427), .Z(n558) );
  XNOR2_X1 U616 ( .A(G1341), .B(G1348), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n560), .B(n559), .ZN(n561) );
  AND2_X1 U619 ( .A1(n561), .A2(G14), .ZN(G401) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  INV_X1 U621 ( .A(G132), .ZN(G219) );
  INV_X1 U622 ( .A(G82), .ZN(G220) );
  NAND2_X1 U623 ( .A1(G88), .A2(n660), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G75), .A2(n664), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G62), .A2(n656), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G50), .A2(n657), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U629 ( .A1(n567), .A2(n566), .ZN(G166) );
  NAND2_X1 U630 ( .A1(n657), .A2(G53), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G91), .A2(n660), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G65), .A2(n656), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n664), .A2(G78), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT72), .B(n570), .Z(n571) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT73), .B(n575), .Z(G299) );
  NAND2_X1 U639 ( .A1(n660), .A2(G89), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT4), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G76), .A2(n664), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT5), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G63), .A2(n656), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G51), .A2(n657), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(KEYINPUT6), .B(n582), .Z(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(G94), .A2(G452), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n586), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n587), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n825) );
  NAND2_X1 U656 ( .A1(n825), .A2(G567), .ZN(n588) );
  XOR2_X1 U657 ( .A(KEYINPUT11), .B(n588), .Z(G234) );
  XOR2_X1 U658 ( .A(G860), .B(KEYINPUT74), .Z(n610) );
  NAND2_X1 U659 ( .A1(G56), .A2(n656), .ZN(n589) );
  XOR2_X1 U660 ( .A(KEYINPUT14), .B(n589), .Z(n595) );
  NAND2_X1 U661 ( .A1(n660), .A2(G81), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G68), .A2(n664), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U665 ( .A(KEYINPUT13), .B(n593), .Z(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n657), .A2(G43), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n929) );
  OR2_X1 U669 ( .A1(n610), .A2(n929), .ZN(G153) );
  NAND2_X1 U670 ( .A1(G301), .A2(G868), .ZN(n607) );
  NAND2_X1 U671 ( .A1(n657), .A2(G54), .ZN(n604) );
  NAND2_X1 U672 ( .A1(G66), .A2(n656), .ZN(n599) );
  NAND2_X1 U673 ( .A1(G79), .A2(n664), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U675 ( .A1(G92), .A2(n660), .ZN(n600) );
  XNOR2_X1 U676 ( .A(KEYINPUT75), .B(n600), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U679 ( .A(KEYINPUT15), .B(n605), .Z(n719) );
  INV_X1 U680 ( .A(G868), .ZN(n676) );
  NAND2_X1 U681 ( .A1(n719), .A2(n676), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(G284) );
  NAND2_X1 U683 ( .A1(G286), .A2(G868), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G299), .A2(n676), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n610), .A2(G559), .ZN(n611) );
  INV_X1 U687 ( .A(n719), .ZN(n928) );
  NAND2_X1 U688 ( .A1(n611), .A2(n928), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n929), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G868), .A2(n928), .ZN(n613) );
  NOR2_X1 U692 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G282) );
  XNOR2_X1 U694 ( .A(G2100), .B(KEYINPUT77), .ZN(n625) );
  NAND2_X1 U695 ( .A1(G135), .A2(n881), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G111), .A2(n878), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n877), .A2(G123), .ZN(n618) );
  XOR2_X1 U699 ( .A(KEYINPUT18), .B(n618), .Z(n619) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n882), .A2(G99), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n985) );
  XOR2_X1 U703 ( .A(G2096), .B(KEYINPUT76), .Z(n623) );
  XNOR2_X1 U704 ( .A(n985), .B(n623), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U706 ( .A(n626), .B(KEYINPUT78), .ZN(G156) );
  NAND2_X1 U707 ( .A1(n928), .A2(G559), .ZN(n674) );
  XOR2_X1 U708 ( .A(KEYINPUT79), .B(n929), .Z(n627) );
  XNOR2_X1 U709 ( .A(n674), .B(n627), .ZN(n628) );
  NOR2_X1 U710 ( .A1(G860), .A2(n628), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G67), .A2(n656), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT80), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G93), .A2(n660), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G80), .A2(n664), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U716 ( .A1(G55), .A2(n657), .ZN(n632) );
  XNOR2_X1 U717 ( .A(KEYINPUT81), .B(n632), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n677) );
  XOR2_X1 U720 ( .A(n637), .B(n677), .Z(G145) );
  NAND2_X1 U721 ( .A1(n656), .A2(G61), .ZN(n638) );
  XNOR2_X1 U722 ( .A(KEYINPUT83), .B(n638), .ZN(n645) );
  NAND2_X1 U723 ( .A1(G86), .A2(n660), .ZN(n639) );
  XNOR2_X1 U724 ( .A(n639), .B(KEYINPUT84), .ZN(n643) );
  XOR2_X1 U725 ( .A(KEYINPUT85), .B(KEYINPUT2), .Z(n641) );
  NAND2_X1 U726 ( .A1(G73), .A2(n664), .ZN(n640) );
  XNOR2_X1 U727 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U730 ( .A(n646), .B(KEYINPUT86), .ZN(n648) );
  NAND2_X1 U731 ( .A1(G48), .A2(n657), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G49), .A2(n657), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U736 ( .A(KEYINPUT82), .B(n651), .ZN(n652) );
  NOR2_X1 U737 ( .A1(n656), .A2(n652), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(G288) );
  NAND2_X1 U740 ( .A1(G60), .A2(n656), .ZN(n659) );
  NAND2_X1 U741 ( .A1(G47), .A2(n657), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U743 ( .A1(G85), .A2(n660), .ZN(n661) );
  XOR2_X1 U744 ( .A(KEYINPUT66), .B(n661), .Z(n662) );
  NOR2_X1 U745 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n664), .A2(G72), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n666), .A2(n665), .ZN(G290) );
  XNOR2_X1 U748 ( .A(G166), .B(G305), .ZN(n669) );
  XNOR2_X1 U749 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n667), .B(G288), .ZN(n668) );
  XNOR2_X1 U751 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(n929), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n671), .B(G299), .ZN(n672) );
  XNOR2_X1 U754 ( .A(n672), .B(G290), .ZN(n673) );
  XNOR2_X1 U755 ( .A(n673), .B(n677), .ZN(n895) );
  XOR2_X1 U756 ( .A(n895), .B(n674), .Z(n675) );
  NAND2_X1 U757 ( .A1(G868), .A2(n675), .ZN(n679) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n679), .A2(n678), .ZN(G295) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n681) );
  NAND2_X1 U761 ( .A1(G2084), .A2(G2078), .ZN(n680) );
  XNOR2_X1 U762 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U766 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U769 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G96), .A2(n687), .ZN(n830) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n830), .ZN(n691) );
  NAND2_X1 U772 ( .A1(G69), .A2(G120), .ZN(n688) );
  NOR2_X1 U773 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U774 ( .A1(G108), .A2(n689), .ZN(n831) );
  NAND2_X1 U775 ( .A1(G567), .A2(n831), .ZN(n690) );
  NAND2_X1 U776 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U777 ( .A(KEYINPUT89), .B(n692), .ZN(G319) );
  INV_X1 U778 ( .A(G319), .ZN(n694) );
  NAND2_X1 U779 ( .A1(G661), .A2(G483), .ZN(n693) );
  NOR2_X1 U780 ( .A1(n694), .A2(n693), .ZN(n827) );
  NAND2_X1 U781 ( .A1(n827), .A2(G36), .ZN(n695) );
  XNOR2_X1 U782 ( .A(KEYINPUT90), .B(n695), .ZN(G176) );
  INV_X1 U783 ( .A(G166), .ZN(G303) );
  AND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n696) );
  NAND2_X1 U785 ( .A1(G8), .A2(n737), .ZN(n770) );
  NOR2_X1 U786 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XOR2_X1 U787 ( .A(n697), .B(KEYINPUT24), .Z(n698) );
  NOR2_X1 U788 ( .A1(n770), .A2(n698), .ZN(n775) );
  NOR2_X1 U789 ( .A1(G1976), .A2(G288), .ZN(n699) );
  XOR2_X1 U790 ( .A(KEYINPUT98), .B(n699), .Z(n939) );
  NOR2_X1 U791 ( .A1(G1971), .A2(G303), .ZN(n757) );
  INV_X1 U792 ( .A(G286), .ZN(n709) );
  NOR2_X1 U793 ( .A1(G1966), .A2(n770), .ZN(n754) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n737), .ZN(n750) );
  NOR2_X1 U795 ( .A1(n754), .A2(n750), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n700), .A2(G8), .ZN(n701) );
  XNOR2_X1 U797 ( .A(n701), .B(KEYINPUT30), .ZN(n702) );
  NOR2_X1 U798 ( .A1(G168), .A2(n702), .ZN(n707) );
  INV_X1 U799 ( .A(n737), .ZN(n712) );
  XOR2_X1 U800 ( .A(KEYINPUT25), .B(G2078), .Z(n912) );
  NAND2_X1 U801 ( .A1(n712), .A2(n912), .ZN(n704) );
  NAND2_X1 U802 ( .A1(G1961), .A2(n737), .ZN(n703) );
  NAND2_X1 U803 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U804 ( .A(KEYINPUT94), .B(n705), .Z(n735) );
  NOR2_X1 U805 ( .A1(n735), .A2(G171), .ZN(n706) );
  NOR2_X1 U806 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U807 ( .A(KEYINPUT31), .B(n708), .Z(n748) );
  OR2_X1 U808 ( .A1(n709), .A2(n748), .ZN(n743) );
  NAND2_X1 U809 ( .A1(G1348), .A2(n737), .ZN(n711) );
  NAND2_X1 U810 ( .A1(G2067), .A2(n712), .ZN(n710) );
  NAND2_X1 U811 ( .A1(n711), .A2(n710), .ZN(n718) );
  NOR2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n717) );
  XOR2_X1 U813 ( .A(G1996), .B(KEYINPUT95), .Z(n911) );
  NAND2_X1 U814 ( .A1(n712), .A2(n911), .ZN(n713) );
  XNOR2_X1 U815 ( .A(KEYINPUT26), .B(n713), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n714), .A2(n520), .ZN(n715) );
  NOR2_X1 U817 ( .A1(n715), .A2(n929), .ZN(n716) );
  NOR2_X1 U818 ( .A1(n717), .A2(n716), .ZN(n721) );
  AND2_X1 U819 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U820 ( .A1(n721), .A2(n720), .ZN(n728) );
  INV_X1 U821 ( .A(G2072), .ZN(n722) );
  XOR2_X1 U822 ( .A(KEYINPUT27), .B(n723), .Z(n725) );
  NAND2_X1 U823 ( .A1(G1956), .A2(n737), .ZN(n724) );
  NAND2_X1 U824 ( .A1(n725), .A2(n724), .ZN(n729) );
  NOR2_X1 U825 ( .A1(G299), .A2(n729), .ZN(n726) );
  XNOR2_X1 U826 ( .A(n726), .B(KEYINPUT96), .ZN(n727) );
  NOR2_X1 U827 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U828 ( .A1(G299), .A2(n729), .ZN(n730) );
  NOR2_X1 U829 ( .A1(n731), .A2(n521), .ZN(n734) );
  NAND2_X1 U830 ( .A1(n735), .A2(G171), .ZN(n747) );
  AND2_X1 U831 ( .A1(n747), .A2(G286), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n746), .A2(n736), .ZN(n742) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n770), .ZN(n739) );
  NOR2_X1 U834 ( .A1(G2090), .A2(n737), .ZN(n738) );
  NOR2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U836 ( .A1(n740), .A2(G303), .ZN(n741) );
  NAND2_X1 U837 ( .A1(n743), .A2(n516), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n744), .A2(G8), .ZN(n745) );
  XOR2_X1 U839 ( .A(KEYINPUT32), .B(n745), .Z(n756) );
  NAND2_X1 U840 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U841 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U842 ( .A1(G8), .A2(n750), .ZN(n751) );
  NAND2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n757), .A2(n767), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n939), .A2(n758), .ZN(n761) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n934) );
  NOR2_X1 U848 ( .A1(n770), .A2(n759), .ZN(n760) );
  XNOR2_X1 U849 ( .A(G1981), .B(G305), .ZN(n945) );
  NOR2_X1 U850 ( .A1(n939), .A2(n770), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n517), .A2(n764), .ZN(n773) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n765) );
  XOR2_X1 U853 ( .A(KEYINPUT99), .B(n765), .Z(n766) );
  NAND2_X1 U854 ( .A1(G8), .A2(n766), .ZN(n769) );
  INV_X1 U855 ( .A(n767), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G160), .A2(G40), .ZN(n776) );
  NOR2_X1 U860 ( .A1(n777), .A2(n776), .ZN(n820) );
  NAND2_X1 U861 ( .A1(G140), .A2(n881), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G104), .A2(n882), .ZN(n778) );
  NAND2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U864 ( .A(KEYINPUT34), .B(n780), .ZN(n786) );
  NAND2_X1 U865 ( .A1(n877), .A2(G128), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G116), .A2(n878), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U868 ( .A(KEYINPUT91), .B(n783), .ZN(n784) );
  XNOR2_X1 U869 ( .A(KEYINPUT35), .B(n784), .ZN(n785) );
  NOR2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U871 ( .A(KEYINPUT36), .B(n787), .ZN(n891) );
  XNOR2_X1 U872 ( .A(G2067), .B(KEYINPUT37), .ZN(n809) );
  NOR2_X1 U873 ( .A1(n891), .A2(n809), .ZN(n991) );
  NAND2_X1 U874 ( .A1(n820), .A2(n991), .ZN(n817) );
  NAND2_X1 U875 ( .A1(G131), .A2(n881), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G107), .A2(n878), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U878 ( .A1(G95), .A2(n882), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G119), .A2(n877), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n868) );
  INV_X1 U882 ( .A(G1991), .ZN(n811) );
  NOR2_X1 U883 ( .A1(n868), .A2(n811), .ZN(n804) );
  NAND2_X1 U884 ( .A1(G105), .A2(n882), .ZN(n794) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n794), .Z(n800) );
  NAND2_X1 U886 ( .A1(G117), .A2(n878), .ZN(n795) );
  XNOR2_X1 U887 ( .A(n795), .B(KEYINPUT92), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G129), .A2(n877), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U890 ( .A(KEYINPUT93), .B(n798), .Z(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n881), .A2(G141), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n888) );
  AND2_X1 U894 ( .A1(n888), .A2(G1996), .ZN(n803) );
  NOR2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n993) );
  INV_X1 U896 ( .A(n820), .ZN(n805) );
  NOR2_X1 U897 ( .A1(n993), .A2(n805), .ZN(n814) );
  INV_X1 U898 ( .A(n814), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n817), .A2(n806), .ZN(n807) );
  XNOR2_X1 U900 ( .A(G1986), .B(G290), .ZN(n931) );
  NAND2_X1 U901 ( .A1(n518), .A2(n808), .ZN(n823) );
  NAND2_X1 U902 ( .A1(n809), .A2(n891), .ZN(n810) );
  XNOR2_X1 U903 ( .A(n810), .B(KEYINPUT100), .ZN(n1001) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n888), .ZN(n996) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n812) );
  AND2_X1 U906 ( .A1(n811), .A2(n868), .ZN(n988) );
  NOR2_X1 U907 ( .A1(n812), .A2(n988), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U909 ( .A1(n996), .A2(n815), .ZN(n816) );
  XNOR2_X1 U910 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n1001), .A2(n819), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U915 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U918 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U921 ( .A(n829), .B(KEYINPUT102), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XOR2_X1 U928 ( .A(KEYINPUT42), .B(G2078), .Z(n833) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2072), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U931 ( .A(n834), .B(G2096), .Z(n836) );
  XNOR2_X1 U932 ( .A(G2084), .B(G2090), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U934 ( .A(G2100), .B(KEYINPUT43), .Z(n838) );
  XNOR2_X1 U935 ( .A(KEYINPUT103), .B(G2678), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U937 ( .A(n840), .B(n839), .Z(G227) );
  XNOR2_X1 U938 ( .A(G1991), .B(KEYINPUT41), .ZN(n850) );
  XOR2_X1 U939 ( .A(G1981), .B(G1966), .Z(n842) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1986), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U942 ( .A(G1976), .B(G1971), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1956), .B(G1961), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U945 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U946 ( .A(KEYINPUT104), .B(G2474), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(G229) );
  NAND2_X1 U949 ( .A1(G124), .A2(n877), .ZN(n851) );
  XOR2_X1 U950 ( .A(KEYINPUT105), .B(n851), .Z(n852) );
  XNOR2_X1 U951 ( .A(n852), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U952 ( .A1(G112), .A2(n878), .ZN(n853) );
  NAND2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U954 ( .A1(G136), .A2(n881), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G100), .A2(n882), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U957 ( .A1(n858), .A2(n857), .ZN(G162) );
  XNOR2_X1 U958 ( .A(G160), .B(G162), .ZN(n867) );
  NAND2_X1 U959 ( .A1(G139), .A2(n881), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G103), .A2(n882), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U962 ( .A(KEYINPUT106), .B(n861), .ZN(n866) );
  NAND2_X1 U963 ( .A1(n877), .A2(G127), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G115), .A2(n878), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U966 ( .A(KEYINPUT47), .B(n864), .Z(n865) );
  NOR2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n1002) );
  XNOR2_X1 U968 ( .A(n867), .B(n1002), .ZN(n871) );
  XOR2_X1 U969 ( .A(G164), .B(n868), .Z(n869) );
  XNOR2_X1 U970 ( .A(n869), .B(n985), .ZN(n870) );
  XOR2_X1 U971 ( .A(n871), .B(n870), .Z(n876) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT107), .B(n874), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n893) );
  NAND2_X1 U977 ( .A1(n877), .A2(G130), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U980 ( .A1(G142), .A2(n881), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G106), .A2(n882), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U986 ( .A(n891), .B(n890), .Z(n892) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U988 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U989 ( .A(n895), .B(G286), .Z(n897) );
  XNOR2_X1 U990 ( .A(n928), .B(G301), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G397) );
  NOR2_X1 U993 ( .A1(G227), .A2(G229), .ZN(n899) );
  XOR2_X1 U994 ( .A(KEYINPUT49), .B(n899), .Z(n900) );
  NAND2_X1 U995 ( .A1(G319), .A2(n900), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G401), .A2(n901), .ZN(n902) );
  XNOR2_X1 U997 ( .A(KEYINPUT110), .B(n902), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U999 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1002 ( .A(G1991), .B(G25), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(G2072), .B(G33), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(G28), .A2(n907), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(KEYINPUT116), .B(G2067), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(G26), .B(n908), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n916) );
  XNOR2_X1 U1009 ( .A(n911), .B(G32), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n912), .B(G27), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(KEYINPUT53), .B(n917), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(G2090), .B(G35), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n918), .B(KEYINPUT115), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n921), .B(KEYINPUT117), .ZN(n924) );
  XOR2_X1 U1018 ( .A(G2084), .B(G34), .Z(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT54), .B(n922), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(KEYINPUT55), .B(KEYINPUT113), .ZN(n1009) );
  XOR2_X1 U1022 ( .A(n925), .B(n1009), .Z(n927) );
  XNOR2_X1 U1023 ( .A(KEYINPUT118), .B(G29), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n983) );
  XNOR2_X1 U1025 ( .A(n928), .B(G1348), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(G1341), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n942) );
  XNOR2_X1 U1029 ( .A(G166), .B(G1971), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(G1956), .B(G299), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1034 ( .A(KEYINPUT121), .B(n940), .Z(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n948) );
  XOR2_X1 U1036 ( .A(G1966), .B(G168), .Z(n943) );
  XNOR2_X1 U1037 ( .A(KEYINPUT120), .B(n943), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1039 ( .A(KEYINPUT57), .B(n946), .Z(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(G1961), .B(G301), .ZN(n949) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G16), .B(KEYINPUT119), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT56), .B(n951), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(n954), .B(KEYINPUT122), .ZN(n980) );
  XNOR2_X1 U1047 ( .A(G5), .B(G1961), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n955), .B(KEYINPUT123), .ZN(n976) );
  XOR2_X1 U1049 ( .A(G1966), .B(G21), .Z(n967) );
  XOR2_X1 U1050 ( .A(G1348), .B(KEYINPUT59), .Z(n956) );
  XNOR2_X1 U1051 ( .A(G4), .B(n956), .ZN(n964) );
  XNOR2_X1 U1052 ( .A(G1341), .B(G19), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G1981), .B(G6), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(KEYINPUT124), .B(n959), .Z(n961) );
  XNOR2_X1 U1056 ( .A(G1956), .B(G20), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(n962), .B(KEYINPUT125), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n965), .B(KEYINPUT60), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G22), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(G23), .B(G1976), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n971) );
  XOR2_X1 U1065 ( .A(G1986), .B(G24), .Z(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(KEYINPUT58), .B(n972), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT61), .B(n977), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n978), .A2(G16), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT126), .B(n984), .ZN(n1014) );
  XNOR2_X1 U1076 ( .A(G160), .B(G2084), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(KEYINPUT111), .B(n989), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n999) );
  XOR2_X1 U1082 ( .A(G2090), .B(G162), .Z(n994) );
  XNOR2_X1 U1083 ( .A(KEYINPUT112), .B(n994), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(KEYINPUT51), .B(n997), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1007) );
  XOR2_X1 U1088 ( .A(G2072), .B(n1002), .Z(n1004) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(KEYINPUT50), .B(n1005), .Z(n1006) );
  NOR2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(KEYINPUT52), .B(n1008), .ZN(n1010) );
  NAND2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1095 ( .A1(n1011), .A2(G29), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(KEYINPUT114), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1097 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(n1015), .B(KEYINPUT62), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(KEYINPUT127), .B(n1016), .ZN(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

