

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734;

  XNOR2_X1 U366 ( .A(n411), .B(n565), .ZN(n711) );
  NOR2_X1 U367 ( .A1(n703), .A2(n707), .ZN(n415) );
  XNOR2_X2 U368 ( .A(n432), .B(KEYINPUT75), .ZN(n642) );
  OR2_X2 U369 ( .A1(n610), .A2(n521), .ZN(n425) );
  NOR2_X2 U370 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X2 U371 ( .A(n526), .B(KEYINPUT0), .ZN(n546) );
  INV_X1 U372 ( .A(n572), .ZN(n669) );
  AND2_X2 U373 ( .A1(n407), .A2(n445), .ZN(n705) );
  AND2_X1 U374 ( .A1(n396), .A2(n393), .ZN(n411) );
  XNOR2_X1 U375 ( .A(n384), .B(KEYINPUT39), .ZN(n612) );
  XNOR2_X1 U376 ( .A(n453), .B(KEYINPUT22), .ZN(n392) );
  NOR2_X1 U377 ( .A1(n546), .A2(n352), .ZN(n453) );
  NOR2_X1 U378 ( .A1(n594), .A2(n669), .ZN(n578) );
  AND2_X1 U379 ( .A1(n425), .A2(n348), .ZN(n424) );
  XNOR2_X1 U380 ( .A(n402), .B(n714), .ZN(n693) );
  XNOR2_X1 U381 ( .A(n404), .B(n403), .ZN(n402) );
  XNOR2_X1 U382 ( .A(G116), .B(KEYINPUT3), .ZN(n431) );
  XNOR2_X1 U383 ( .A(n430), .B(n429), .ZN(n387) );
  XNOR2_X1 U384 ( .A(G113), .B(KEYINPUT70), .ZN(n429) );
  XNOR2_X1 U385 ( .A(n502), .B(n431), .ZN(n430) );
  XNOR2_X1 U386 ( .A(G119), .B(KEYINPUT84), .ZN(n502) );
  XNOR2_X1 U387 ( .A(n488), .B(n487), .ZN(n516) );
  INV_X1 U388 ( .A(KEYINPUT4), .ZN(n487) );
  AND2_X1 U389 ( .A1(n616), .A2(n446), .ZN(n407) );
  INV_X1 U390 ( .A(n617), .ZN(n446) );
  XNOR2_X1 U391 ( .A(n540), .B(n493), .ZN(n722) );
  XNOR2_X1 U392 ( .A(n490), .B(n489), .ZN(n512) );
  XNOR2_X1 U393 ( .A(n498), .B(n497), .ZN(n386) );
  NOR2_X1 U394 ( .A1(G902), .A2(n698), .ZN(n498) );
  OR2_X1 U395 ( .A1(n359), .A2(n356), .ZN(n549) );
  NAND2_X1 U396 ( .A1(n361), .A2(n360), .ZN(n359) );
  NAND2_X1 U397 ( .A1(n362), .A2(G902), .ZN(n360) );
  XNOR2_X1 U398 ( .A(n721), .B(n419), .ZN(n621) );
  XNOR2_X1 U399 ( .A(n506), .B(n501), .ZN(n419) );
  XNOR2_X1 U400 ( .A(n387), .B(n505), .ZN(n506) );
  XNOR2_X1 U401 ( .A(n516), .B(n444), .ZN(n721) );
  XNOR2_X1 U402 ( .A(G131), .B(G134), .ZN(n444) );
  NAND2_X1 U403 ( .A1(n615), .A2(n711), .ZN(n616) );
  AND2_X1 U404 ( .A1(n385), .A2(n343), .ZN(n615) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n541) );
  XOR2_X1 U406 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n535) );
  XNOR2_X1 U407 ( .A(G104), .B(G143), .ZN(n534) );
  XNOR2_X1 U408 ( .A(n364), .B(G113), .ZN(n462) );
  INV_X1 U409 ( .A(G140), .ZN(n364) );
  NAND2_X1 U410 ( .A1(n366), .A2(KEYINPUT48), .ZN(n365) );
  INV_X1 U411 ( .A(n654), .ZN(n374) );
  INV_X1 U412 ( .A(G122), .ZN(n401) );
  INV_X1 U413 ( .A(KEYINPUT72), .ZN(n383) );
  NAND2_X1 U414 ( .A1(n571), .A2(n383), .ZN(n382) );
  XNOR2_X1 U415 ( .A(n437), .B(n722), .ZN(n706) );
  XNOR2_X1 U416 ( .A(n484), .B(n438), .ZN(n437) );
  XNOR2_X1 U417 ( .A(n483), .B(n439), .ZN(n438) );
  XNOR2_X1 U418 ( .A(n459), .B(n539), .ZN(n700) );
  XNOR2_X1 U419 ( .A(n460), .B(n540), .ZN(n459) );
  INV_X1 U420 ( .A(n516), .ZN(n403) );
  NAND2_X1 U421 ( .A1(n600), .A2(n574), .ZN(n384) );
  NAND2_X1 U422 ( .A1(n363), .A2(n641), .ZN(n607) );
  AND2_X1 U423 ( .A1(n418), .A2(n655), .ZN(n363) );
  BUF_X1 U424 ( .A(n670), .Z(n413) );
  AND2_X1 U425 ( .A1(n545), .A2(n550), .ZN(n592) );
  XNOR2_X1 U426 ( .A(n443), .B(n441), .ZN(n601) );
  XNOR2_X1 U427 ( .A(n573), .B(n442), .ZN(n441) );
  NAND2_X1 U428 ( .A1(n572), .A2(n655), .ZN(n443) );
  INV_X1 U429 ( .A(KEYINPUT107), .ZN(n442) );
  XNOR2_X1 U430 ( .A(n549), .B(n457), .ZN(n545) );
  INV_X1 U431 ( .A(KEYINPUT98), .ZN(n457) );
  XNOR2_X1 U432 ( .A(n621), .B(KEYINPUT62), .ZN(n623) );
  NAND2_X1 U433 ( .A1(n705), .A2(G217), .ZN(n452) );
  XNOR2_X1 U434 ( .A(n492), .B(n496), .ZN(n391) );
  XNOR2_X1 U435 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U436 ( .A(n491), .B(n501), .ZN(n492) );
  NOR2_X1 U437 ( .A1(n355), .A2(n354), .ZN(n422) );
  NOR2_X1 U438 ( .A1(n689), .A2(n345), .ZN(n408) );
  INV_X2 U439 ( .A(G953), .ZN(n416) );
  NOR2_X1 U440 ( .A1(n642), .A2(n587), .ZN(n390) );
  NAND2_X1 U441 ( .A1(n458), .A2(n358), .ZN(n357) );
  INV_X1 U442 ( .A(G902), .ZN(n358) );
  NAND2_X1 U443 ( .A1(n700), .A2(n362), .ZN(n361) );
  XOR2_X1 U444 ( .A(G137), .B(KEYINPUT5), .Z(n504) );
  INV_X1 U445 ( .A(KEYINPUT44), .ZN(n564) );
  AND2_X1 U446 ( .A1(n394), .A2(n628), .ZN(n393) );
  XNOR2_X1 U447 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n439) );
  XNOR2_X1 U448 ( .A(n511), .B(n480), .ZN(n540) );
  XNOR2_X1 U449 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n480) );
  XNOR2_X1 U450 ( .A(n543), .B(n461), .ZN(n460) );
  XNOR2_X1 U451 ( .A(n462), .B(n542), .ZN(n461) );
  XOR2_X1 U452 ( .A(KEYINPUT66), .B(G101), .Z(n510) );
  XNOR2_X1 U453 ( .A(G137), .B(G140), .ZN(n493) );
  NAND2_X1 U454 ( .A1(n373), .A2(KEYINPUT48), .ZN(n372) );
  AND2_X1 U455 ( .A1(n711), .A2(n455), .ZN(n454) );
  INV_X1 U456 ( .A(KEYINPUT77), .ZN(n455) );
  XNOR2_X1 U457 ( .A(n596), .B(KEYINPUT38), .ZN(n656) );
  OR2_X1 U458 ( .A1(G902), .A2(G237), .ZN(n518) );
  XNOR2_X1 U459 ( .A(G902), .B(KEYINPUT15), .ZN(n617) );
  NOR2_X1 U460 ( .A1(G902), .A2(n706), .ZN(n485) );
  XNOR2_X1 U461 ( .A(n512), .B(n400), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n513), .B(n401), .ZN(n400) );
  INV_X1 U463 ( .A(KEYINPUT16), .ZN(n513) );
  XNOR2_X1 U464 ( .A(n347), .B(n464), .ZN(n488) );
  XNOR2_X1 U465 ( .A(G128), .B(KEYINPUT64), .ZN(n464) );
  XNOR2_X1 U466 ( .A(G107), .B(KEYINPUT7), .ZN(n466) );
  XOR2_X1 U467 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n467) );
  XNOR2_X1 U468 ( .A(G116), .B(G122), .ZN(n465) );
  NAND2_X1 U469 ( .A1(n380), .A2(n378), .ZN(n600) );
  NAND2_X1 U470 ( .A1(n379), .A2(n350), .ZN(n378) );
  AND2_X1 U471 ( .A1(n382), .A2(n381), .ZN(n380) );
  OR2_X1 U472 ( .A1(n655), .A2(n521), .ZN(n428) );
  AND2_X1 U473 ( .A1(n655), .A2(n521), .ZN(n427) );
  NOR2_X1 U474 ( .A1(G902), .A2(n621), .ZN(n508) );
  XNOR2_X1 U475 ( .A(n700), .B(n463), .ZN(n701) );
  XNOR2_X1 U476 ( .A(n580), .B(n414), .ZN(n734) );
  INV_X1 U477 ( .A(KEYINPUT42), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n412), .B(KEYINPUT40), .ZN(n377) );
  NOR2_X1 U479 ( .A1(n607), .A2(n596), .ZN(n598) );
  XNOR2_X1 U480 ( .A(n410), .B(n409), .ZN(n731) );
  INV_X1 U481 ( .A(KEYINPUT35), .ZN(n409) );
  NOR2_X1 U482 ( .A1(n624), .A2(n707), .ZN(n627) );
  INV_X1 U483 ( .A(KEYINPUT122), .ZN(n448) );
  NAND2_X1 U484 ( .A1(n450), .A2(n420), .ZN(n449) );
  XNOR2_X1 U485 ( .A(n452), .B(n451), .ZN(n450) );
  XNOR2_X1 U486 ( .A(n696), .B(n406), .ZN(n699) );
  XNOR2_X1 U487 ( .A(n698), .B(n697), .ZN(n406) );
  AND2_X1 U488 ( .A1(n421), .A2(n420), .ZN(n695) );
  XNOR2_X1 U489 ( .A(n422), .B(n440), .ZN(n421) );
  XNOR2_X1 U490 ( .A(n694), .B(n692), .ZN(n440) );
  AND2_X1 U491 ( .A1(n417), .A2(n416), .ZN(n691) );
  AND2_X1 U492 ( .A1(n688), .A2(n408), .ZN(n690) );
  XNOR2_X1 U493 ( .A(n500), .B(n499), .ZN(n571) );
  XOR2_X1 U494 ( .A(n486), .B(n485), .Z(n576) );
  AND2_X1 U495 ( .A1(n614), .A2(KEYINPUT2), .ZN(n343) );
  AND2_X1 U496 ( .A1(n426), .A2(n428), .ZN(n344) );
  XOR2_X1 U497 ( .A(n687), .B(KEYINPUT117), .Z(n345) );
  XOR2_X1 U498 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n346) );
  XOR2_X1 U499 ( .A(G143), .B(KEYINPUT76), .Z(n347) );
  OR2_X1 U500 ( .A1(n570), .A2(n525), .ZN(n348) );
  NOR2_X1 U501 ( .A1(n577), .A2(n435), .ZN(n349) );
  INV_X1 U502 ( .A(n458), .ZN(n362) );
  XNOR2_X1 U503 ( .A(n544), .B(G475), .ZN(n458) );
  NOR2_X1 U504 ( .A1(n577), .A2(n383), .ZN(n350) );
  AND2_X1 U505 ( .A1(n344), .A2(n425), .ZN(n351) );
  OR2_X1 U506 ( .A1(n659), .A2(n435), .ZN(n352) );
  XNOR2_X1 U507 ( .A(n391), .B(n721), .ZN(n698) );
  XOR2_X1 U508 ( .A(n531), .B(KEYINPUT120), .Z(n353) );
  INV_X1 U509 ( .A(KEYINPUT48), .ZN(n375) );
  INV_X1 U510 ( .A(KEYINPUT2), .ZN(n613) );
  NOR2_X1 U511 ( .A1(G952), .A2(n416), .ZN(n707) );
  INV_X1 U512 ( .A(n707), .ZN(n420) );
  INV_X1 U513 ( .A(n445), .ZN(n354) );
  NAND2_X1 U514 ( .A1(n407), .A2(G210), .ZN(n355) );
  NOR2_X1 U515 ( .A1(n700), .A2(n357), .ZN(n356) );
  NAND2_X1 U516 ( .A1(n365), .A2(n374), .ZN(n370) );
  NAND2_X1 U517 ( .A1(n367), .A2(n591), .ZN(n366) );
  INV_X1 U518 ( .A(n366), .ZN(n376) );
  AND2_X1 U519 ( .A1(n590), .A2(n640), .ZN(n367) );
  NAND2_X1 U520 ( .A1(n372), .A2(n368), .ZN(n371) );
  NAND2_X1 U521 ( .A1(n376), .A2(n369), .ZN(n368) );
  AND2_X1 U522 ( .A1(n606), .A2(n375), .ZN(n369) );
  NOR2_X2 U523 ( .A1(n371), .A2(n370), .ZN(n385) );
  INV_X1 U524 ( .A(n606), .ZN(n373) );
  NAND2_X1 U525 ( .A1(n377), .A2(n734), .ZN(n582) );
  XNOR2_X1 U526 ( .A(n377), .B(G131), .ZN(G33) );
  INV_X1 U527 ( .A(n571), .ZN(n379) );
  NAND2_X1 U528 ( .A1(n577), .A2(n383), .ZN(n381) );
  NAND2_X1 U529 ( .A1(n385), .A2(n652), .ZN(n723) );
  NAND2_X1 U530 ( .A1(n386), .A2(n671), .ZN(n500) );
  XNOR2_X1 U531 ( .A(n386), .B(KEYINPUT1), .ZN(n670) );
  NAND2_X1 U532 ( .A1(n579), .A2(n386), .ZN(n583) );
  XNOR2_X1 U533 ( .A(n399), .B(n387), .ZN(n714) );
  NAND2_X1 U534 ( .A1(n388), .A2(n585), .ZN(n589) );
  XNOR2_X1 U535 ( .A(n390), .B(n389), .ZN(n388) );
  INV_X1 U536 ( .A(KEYINPUT78), .ZN(n389) );
  NAND2_X1 U537 ( .A1(n392), .A2(n593), .ZN(n562) );
  NAND2_X1 U538 ( .A1(n392), .A2(n436), .ZN(n557) );
  NAND2_X1 U539 ( .A1(n395), .A2(n586), .ZN(n394) );
  NAND2_X1 U540 ( .A1(n648), .A2(n632), .ZN(n395) );
  XNOR2_X1 U541 ( .A(n397), .B(n564), .ZN(n396) );
  NAND2_X1 U542 ( .A1(n398), .A2(n731), .ZN(n397) );
  NOR2_X1 U543 ( .A1(n733), .A2(n423), .ZN(n398) );
  XNOR2_X1 U544 ( .A(n517), .B(n405), .ZN(n404) );
  XNOR2_X1 U545 ( .A(n515), .B(KEYINPUT81), .ZN(n405) );
  XNOR2_X1 U546 ( .A(n618), .B(n353), .ZN(n619) );
  XNOR2_X1 U547 ( .A(n622), .B(n623), .ZN(n624) );
  NAND2_X2 U548 ( .A1(n447), .A2(n613), .ZN(n445) );
  NAND2_X1 U549 ( .A1(n424), .A2(n344), .ZN(n526) );
  NAND2_X1 U550 ( .A1(n556), .A2(n604), .ZN(n410) );
  NAND2_X1 U551 ( .A1(n656), .A2(n655), .ZN(n660) );
  INV_X1 U552 ( .A(n666), .ZN(n435) );
  NAND2_X1 U553 ( .A1(n612), .A2(n592), .ZN(n412) );
  XNOR2_X1 U554 ( .A(n415), .B(n704), .ZN(G60) );
  XNOR2_X1 U555 ( .A(n690), .B(KEYINPUT118), .ZN(n417) );
  XNOR2_X1 U556 ( .A(n651), .B(KEYINPUT80), .ZN(n606) );
  NAND2_X1 U557 ( .A1(n599), .A2(n413), .ZN(n651) );
  XNOR2_X1 U558 ( .A(n595), .B(KEYINPUT106), .ZN(n418) );
  INV_X1 U559 ( .A(n636), .ZN(n423) );
  NAND2_X1 U560 ( .A1(n610), .A2(n427), .ZN(n426) );
  XNOR2_X2 U561 ( .A(n520), .B(n519), .ZN(n610) );
  NAND2_X1 U562 ( .A1(n433), .A2(n351), .ZN(n432) );
  INV_X1 U563 ( .A(n583), .ZN(n433) );
  XNOR2_X1 U564 ( .A(n434), .B(KEYINPUT68), .ZN(n594) );
  NAND2_X1 U565 ( .A1(n436), .A2(n349), .ZN(n434) );
  INV_X1 U566 ( .A(n576), .ZN(n436) );
  XNOR2_X2 U567 ( .A(n508), .B(n507), .ZN(n572) );
  NAND2_X1 U568 ( .A1(n445), .A2(n616), .ZN(n688) );
  NAND2_X1 U569 ( .A1(n454), .A2(n456), .ZN(n447) );
  XNOR2_X1 U570 ( .A(n449), .B(n448), .ZN(G66) );
  INV_X1 U571 ( .A(n706), .ZN(n451) );
  INV_X1 U572 ( .A(n723), .ZN(n456) );
  XNOR2_X1 U573 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U574 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n463) );
  XNOR2_X1 U575 ( .A(KEYINPUT46), .B(KEYINPUT79), .ZN(n581) );
  INV_X1 U576 ( .A(n512), .ZN(n491) );
  INV_X1 U577 ( .A(KEYINPUT45), .ZN(n565) );
  NAND2_X1 U578 ( .A1(n705), .A2(G472), .ZN(n622) );
  INV_X1 U579 ( .A(KEYINPUT63), .ZN(n625) );
  XNOR2_X1 U580 ( .A(n625), .B(KEYINPUT82), .ZN(n626) );
  NAND2_X1 U581 ( .A1(n619), .A2(n420), .ZN(n620) );
  XNOR2_X1 U582 ( .A(n620), .B(KEYINPUT121), .ZN(G63) );
  XNOR2_X1 U583 ( .A(n465), .B(G134), .ZN(n469) );
  XNOR2_X1 U584 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U585 ( .A(n469), .B(n468), .Z(n472) );
  NAND2_X1 U586 ( .A1(G234), .A2(n416), .ZN(n470) );
  XOR2_X1 U587 ( .A(KEYINPUT8), .B(n470), .Z(n479) );
  NAND2_X1 U588 ( .A1(G217), .A2(n479), .ZN(n471) );
  XNOR2_X1 U589 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U590 ( .A(n488), .B(n473), .ZN(n531) );
  NAND2_X1 U591 ( .A1(G234), .A2(n617), .ZN(n474) );
  XNOR2_X1 U592 ( .A(KEYINPUT20), .B(n474), .ZN(n476) );
  NAND2_X1 U593 ( .A1(n476), .A2(G221), .ZN(n475) );
  XOR2_X1 U594 ( .A(KEYINPUT21), .B(n475), .Z(n666) );
  XOR2_X1 U595 ( .A(KEYINPUT25), .B(KEYINPUT90), .Z(n478) );
  NAND2_X1 U596 ( .A1(n476), .A2(G217), .ZN(n477) );
  XNOR2_X1 U597 ( .A(n478), .B(n477), .ZN(n486) );
  NAND2_X1 U598 ( .A1(n479), .A2(G221), .ZN(n484) );
  XOR2_X1 U599 ( .A(G125), .B(G146), .Z(n511) );
  XOR2_X1 U600 ( .A(KEYINPUT89), .B(G128), .Z(n482) );
  XNOR2_X1 U601 ( .A(G119), .B(G110), .ZN(n481) );
  XNOR2_X1 U602 ( .A(n482), .B(n481), .ZN(n483) );
  AND2_X1 U603 ( .A1(n666), .A2(n576), .ZN(n671) );
  XOR2_X1 U604 ( .A(G104), .B(G107), .Z(n490) );
  XNOR2_X1 U605 ( .A(G110), .B(KEYINPUT83), .ZN(n489) );
  XNOR2_X1 U606 ( .A(G146), .B(n510), .ZN(n501) );
  INV_X1 U607 ( .A(n493), .ZN(n495) );
  NAND2_X1 U608 ( .A1(G227), .A2(n416), .ZN(n494) );
  XNOR2_X1 U609 ( .A(KEYINPUT69), .B(G469), .ZN(n497) );
  INV_X1 U610 ( .A(KEYINPUT91), .ZN(n499) );
  NAND2_X1 U611 ( .A1(n541), .A2(G210), .ZN(n503) );
  XNOR2_X1 U612 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U613 ( .A(KEYINPUT71), .B(G472), .ZN(n507) );
  NAND2_X1 U614 ( .A1(n518), .A2(G214), .ZN(n509) );
  XOR2_X1 U615 ( .A(KEYINPUT85), .B(n509), .Z(n655) );
  XNOR2_X1 U616 ( .A(n511), .B(n510), .ZN(n517) );
  NAND2_X1 U617 ( .A1(G224), .A2(n416), .ZN(n514) );
  XNOR2_X1 U618 ( .A(n346), .B(n514), .ZN(n515) );
  NAND2_X1 U619 ( .A1(n693), .A2(n617), .ZN(n520) );
  AND2_X1 U620 ( .A1(G210), .A2(n518), .ZN(n519) );
  XOR2_X1 U621 ( .A(KEYINPUT73), .B(KEYINPUT19), .Z(n521) );
  NAND2_X1 U622 ( .A1(G237), .A2(G234), .ZN(n522) );
  XNOR2_X1 U623 ( .A(n522), .B(KEYINPUT86), .ZN(n523) );
  XNOR2_X1 U624 ( .A(KEYINPUT14), .B(n523), .ZN(n524) );
  NAND2_X1 U625 ( .A1(G952), .A2(n524), .ZN(n684) );
  NOR2_X1 U626 ( .A1(G953), .A2(n684), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G902), .A2(n524), .ZN(n566) );
  XNOR2_X1 U628 ( .A(G898), .B(KEYINPUT87), .ZN(n710) );
  NAND2_X1 U629 ( .A1(G953), .A2(n710), .ZN(n715) );
  NOR2_X1 U630 ( .A1(n566), .A2(n715), .ZN(n525) );
  XNOR2_X1 U631 ( .A(n546), .B(KEYINPUT88), .ZN(n553) );
  NOR2_X1 U632 ( .A1(n572), .A2(n553), .ZN(n527) );
  NAND2_X1 U633 ( .A1(n379), .A2(n527), .ZN(n632) );
  NAND2_X1 U634 ( .A1(n670), .A2(n671), .ZN(n551) );
  OR2_X1 U635 ( .A1(n669), .A2(n551), .ZN(n676) );
  NOR2_X1 U636 ( .A1(n546), .A2(n676), .ZN(n529) );
  XNOR2_X1 U637 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n528) );
  XNOR2_X1 U638 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U639 ( .A(KEYINPUT92), .B(n530), .Z(n648) );
  NOR2_X1 U640 ( .A1(G902), .A2(n531), .ZN(n533) );
  XNOR2_X1 U641 ( .A(KEYINPUT100), .B(G478), .ZN(n532) );
  XNOR2_X1 U642 ( .A(n533), .B(n532), .ZN(n550) );
  XNOR2_X1 U643 ( .A(n535), .B(n534), .ZN(n543) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n537) );
  XNOR2_X1 U645 ( .A(G131), .B(KEYINPUT94), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U647 ( .A(n538), .B(G122), .Z(n539) );
  NAND2_X1 U648 ( .A1(n541), .A2(G214), .ZN(n542) );
  XNOR2_X1 U649 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n544) );
  NOR2_X1 U650 ( .A1(n550), .A2(n545), .ZN(n637) );
  XOR2_X1 U651 ( .A(KEYINPUT101), .B(n637), .Z(n611) );
  NOR2_X1 U652 ( .A1(n592), .A2(n611), .ZN(n661) );
  INV_X1 U653 ( .A(n661), .ZN(n586) );
  INV_X1 U654 ( .A(n413), .ZN(n559) );
  XOR2_X1 U655 ( .A(KEYINPUT102), .B(n436), .Z(n665) );
  INV_X1 U656 ( .A(n665), .ZN(n547) );
  XNOR2_X1 U657 ( .A(n572), .B(KEYINPUT6), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n550), .A2(n549), .ZN(n659) );
  NOR2_X1 U659 ( .A1(n547), .A2(n562), .ZN(n548) );
  NAND2_X1 U660 ( .A1(n559), .A2(n548), .ZN(n628) );
  NOR2_X1 U661 ( .A1(n550), .A2(n549), .ZN(n604) );
  NOR2_X1 U662 ( .A1(n551), .A2(n593), .ZN(n552) );
  XNOR2_X1 U663 ( .A(n552), .B(KEYINPUT33), .ZN(n685) );
  NOR2_X1 U664 ( .A1(n553), .A2(n685), .ZN(n555) );
  XNOR2_X1 U665 ( .A(KEYINPUT34), .B(KEYINPUT74), .ZN(n554) );
  XNOR2_X1 U666 ( .A(n555), .B(n554), .ZN(n556) );
  NOR2_X1 U667 ( .A1(n572), .A2(n557), .ZN(n558) );
  NAND2_X1 U668 ( .A1(n559), .A2(n558), .ZN(n636) );
  NOR2_X1 U669 ( .A1(n559), .A2(n665), .ZN(n560) );
  XNOR2_X1 U670 ( .A(n560), .B(KEYINPUT103), .ZN(n561) );
  XNOR2_X1 U671 ( .A(KEYINPUT32), .B(n563), .ZN(n733) );
  NOR2_X1 U672 ( .A1(G900), .A2(n566), .ZN(n567) );
  NAND2_X1 U673 ( .A1(G953), .A2(n567), .ZN(n568) );
  XNOR2_X1 U674 ( .A(KEYINPUT105), .B(n568), .ZN(n569) );
  NOR2_X1 U675 ( .A1(n570), .A2(n569), .ZN(n577) );
  XOR2_X1 U676 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n573) );
  INV_X1 U677 ( .A(n610), .ZN(n596) );
  AND2_X1 U678 ( .A1(n601), .A2(n656), .ZN(n574) );
  NOR2_X1 U679 ( .A1(n659), .A2(n660), .ZN(n575) );
  XNOR2_X1 U680 ( .A(n575), .B(KEYINPUT41), .ZN(n686) );
  XNOR2_X1 U681 ( .A(n578), .B(KEYINPUT28), .ZN(n579) );
  NOR2_X1 U682 ( .A1(n686), .A2(n583), .ZN(n580) );
  XNOR2_X1 U683 ( .A(n582), .B(n581), .ZN(n591) );
  INV_X1 U684 ( .A(KEYINPUT47), .ZN(n587) );
  NOR2_X1 U685 ( .A1(KEYINPUT47), .A2(n661), .ZN(n584) );
  NAND2_X1 U686 ( .A1(n642), .A2(n584), .ZN(n585) );
  NOR2_X1 U687 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U688 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U689 ( .A(KEYINPUT104), .B(n592), .ZN(n641) );
  INV_X1 U690 ( .A(n641), .ZN(n645) );
  NOR2_X1 U691 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U692 ( .A(KEYINPUT36), .B(KEYINPUT110), .ZN(n597) );
  XNOR2_X1 U693 ( .A(n598), .B(n597), .ZN(n599) );
  AND2_X1 U694 ( .A1(n600), .A2(n601), .ZN(n602) );
  NAND2_X1 U695 ( .A1(n610), .A2(n602), .ZN(n603) );
  XNOR2_X1 U696 ( .A(KEYINPUT109), .B(n603), .ZN(n605) );
  NAND2_X1 U697 ( .A1(n605), .A2(n604), .ZN(n640) );
  NOR2_X1 U698 ( .A1(n413), .A2(n607), .ZN(n608) );
  XNOR2_X1 U699 ( .A(n608), .B(KEYINPUT43), .ZN(n609) );
  NOR2_X1 U700 ( .A1(n610), .A2(n609), .ZN(n654) );
  NAND2_X1 U701 ( .A1(n612), .A2(n611), .ZN(n652) );
  XOR2_X1 U702 ( .A(n652), .B(KEYINPUT77), .Z(n614) );
  NAND2_X1 U703 ( .A1(G478), .A2(n705), .ZN(n618) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(G57) );
  XNOR2_X1 U705 ( .A(G101), .B(n628), .ZN(G3) );
  NOR2_X1 U706 ( .A1(n645), .A2(n632), .ZN(n630) );
  XNOR2_X1 U707 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U709 ( .A(G104), .B(n631), .ZN(G6) );
  INV_X1 U710 ( .A(n637), .ZN(n647) );
  NOR2_X1 U711 ( .A1(n647), .A2(n632), .ZN(n634) );
  XNOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U714 ( .A(G107), .B(n635), .ZN(G9) );
  XNOR2_X1 U715 ( .A(G110), .B(n636), .ZN(G12) );
  XOR2_X1 U716 ( .A(G128), .B(KEYINPUT29), .Z(n639) );
  NAND2_X1 U717 ( .A1(n637), .A2(n642), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n639), .B(n638), .ZN(G30) );
  XNOR2_X1 U719 ( .A(G143), .B(n640), .ZN(G45) );
  XOR2_X1 U720 ( .A(G146), .B(KEYINPUT113), .Z(n644) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n644), .B(n643), .ZN(G48) );
  NOR2_X1 U723 ( .A1(n645), .A2(n648), .ZN(n646) );
  XOR2_X1 U724 ( .A(G113), .B(n646), .Z(G15) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U726 ( .A(G116), .B(n649), .Z(G18) );
  XOR2_X1 U727 ( .A(G125), .B(KEYINPUT37), .Z(n650) );
  XNOR2_X1 U728 ( .A(n651), .B(n650), .ZN(G27) );
  XNOR2_X1 U729 ( .A(G134), .B(KEYINPUT114), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(G36) );
  XOR2_X1 U731 ( .A(G140), .B(n654), .Z(G42) );
  NOR2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n657), .B(KEYINPUT116), .ZN(n658) );
  NOR2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n663) );
  NOR2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U737 ( .A1(n664), .A2(n685), .ZN(n681) );
  NOR2_X1 U738 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n667), .B(KEYINPUT49), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n674) );
  NOR2_X1 U741 ( .A1(n671), .A2(n413), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(KEYINPUT50), .ZN(n673) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n675), .B(KEYINPUT115), .ZN(n677) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U746 ( .A(KEYINPUT51), .B(n678), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n679), .A2(n686), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U752 ( .A(KEYINPUT53), .B(n691), .ZN(G75) );
  XOR2_X1 U753 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n692) );
  INV_X1 U754 ( .A(n693), .ZN(n694) );
  XNOR2_X1 U755 ( .A(KEYINPUT56), .B(n695), .ZN(G51) );
  XOR2_X1 U756 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n697) );
  NAND2_X1 U757 ( .A1(n705), .A2(G469), .ZN(n696) );
  NOR2_X1 U758 ( .A1(n707), .A2(n699), .ZN(G54) );
  NAND2_X1 U759 ( .A1(n705), .A2(G475), .ZN(n702) );
  XOR2_X1 U760 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n704) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n708) );
  XOR2_X1 U762 ( .A(KEYINPUT61), .B(n708), .Z(n709) );
  NOR2_X1 U763 ( .A1(n710), .A2(n709), .ZN(n713) );
  AND2_X1 U764 ( .A1(n711), .A2(n416), .ZN(n712) );
  NOR2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n720) );
  XOR2_X1 U766 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n718) );
  XOR2_X1 U767 ( .A(n714), .B(G101), .Z(n716) );
  NAND2_X1 U768 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(G69) );
  XNOR2_X1 U771 ( .A(n721), .B(n722), .ZN(n725) );
  XOR2_X1 U772 ( .A(n723), .B(n725), .Z(n724) );
  NAND2_X1 U773 ( .A1(n724), .A2(n416), .ZN(n730) );
  XNOR2_X1 U774 ( .A(n725), .B(G227), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n726), .B(KEYINPUT125), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U777 ( .A1(G953), .A2(n728), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n730), .A2(n729), .ZN(G72) );
  XNOR2_X1 U779 ( .A(n731), .B(G122), .ZN(G24) );
  XOR2_X1 U780 ( .A(G119), .B(KEYINPUT126), .Z(n732) );
  XNOR2_X1 U781 ( .A(n733), .B(n732), .ZN(G21) );
  XNOR2_X1 U782 ( .A(n734), .B(G137), .ZN(G39) );
endmodule

