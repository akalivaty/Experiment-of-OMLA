//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n203), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(G58), .A2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n206), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  INV_X1    g0039(.A(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G77), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(G1698), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT66), .ZN(new_n263));
  INV_X1    g0063(.A(G223), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n254), .B(new_n261), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(G1), .A2(G13), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(G274), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n275), .A2(new_n274), .B1(new_n266), .B2(new_n267), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n218), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n270), .A2(new_n271), .A3(new_n276), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n217), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n226), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G50), .A3(new_n282), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n227), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G150), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI22_X1  g0094(.A1(new_n290), .A2(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n296));
  OAI21_X1  g0096(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n286), .A2(new_n226), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n285), .B(new_n289), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI211_X1 g0104(.A(new_n304), .B(new_n279), .C1(new_n265), .C2(new_n269), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n281), .B(new_n301), .C1(new_n305), .C2(G169), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n270), .A2(new_n276), .A3(new_n280), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G200), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT9), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n270), .A2(G190), .A3(new_n276), .A4(new_n280), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n301), .A2(new_n310), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n309), .A2(new_n311), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n308), .A2(G200), .B1(new_n310), .B2(new_n301), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n311), .A4(new_n312), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n307), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n259), .A2(G226), .A3(new_n260), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n304), .B1(new_n323), .B2(new_n269), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n277), .A2(G238), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  OAI211_X1 g0130(.A(KEYINPUT70), .B(KEYINPUT14), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(G179), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT70), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  OAI221_X1 g0134(.A(G169), .B1(new_n333), .B2(new_n334), .C1(new_n327), .C2(new_n328), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n294), .A2(new_n217), .B1(new_n227), .B2(G68), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n291), .A2(new_n219), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n287), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT69), .B(KEYINPUT11), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n227), .A2(G1), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G13), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n300), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT68), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n300), .A2(new_n343), .A3(KEYINPUT68), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G68), .ZN(new_n349));
  INV_X1    g0149(.A(G68), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n284), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT12), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n341), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n336), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n353), .B1(new_n329), .B2(G190), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n355), .B1(new_n356), .B2(new_n329), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(G77), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT15), .B(G87), .Z(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n291), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n290), .A2(new_n294), .B1(new_n227), .B2(new_n219), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n287), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n358), .B(new_n363), .C1(G77), .C2(new_n343), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n278), .A2(new_n220), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n366));
  INV_X1    g0166(.A(G238), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n213), .B2(new_n259), .C1(new_n263), .C2(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n304), .B(new_n365), .C1(new_n368), .C2(new_n269), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n364), .B1(new_n369), .B2(G190), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n269), .ZN(new_n371));
  INV_X1    g0171(.A(new_n365), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n276), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n319), .A2(new_n354), .A3(new_n357), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n257), .A2(new_n227), .A3(new_n258), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n258), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n350), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G58), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n350), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n229), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n293), .A2(G159), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n377), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT7), .B1(new_n253), .B2(new_n227), .ZN(new_n389));
  INV_X1    g0189(.A(new_n381), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n387), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n393), .A3(new_n287), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n290), .A2(new_n342), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT71), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n288), .B1(new_n284), .B2(new_n290), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n264), .A2(new_n260), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n218), .A2(G1698), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n251), .C2(new_n252), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n269), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n304), .B1(new_n277), .B2(G232), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n271), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n268), .B1(new_n401), .B2(new_n402), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n268), .A2(G232), .A3(new_n302), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n276), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n330), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT18), .B1(new_n398), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  AOI211_X1 g0214(.A(new_n414), .B(new_n411), .C1(new_n394), .C2(new_n397), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT72), .ZN(new_n417));
  OAI21_X1  g0217(.A(G200), .B1(new_n407), .B2(new_n409), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n404), .A2(G190), .A3(new_n405), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n394), .A2(new_n397), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n420), .A2(new_n421), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n417), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n394), .A2(new_n397), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n425), .A2(KEYINPUT17), .A3(new_n418), .A4(new_n419), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n420), .A2(new_n421), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(KEYINPUT72), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n416), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n371), .A2(new_n271), .A3(new_n276), .A4(new_n372), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n364), .C1(new_n369), .C2(G169), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n376), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G283), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n220), .B1(new_n257), .B2(new_n258), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(KEYINPUT4), .ZN(new_n436));
  OAI211_X1 g0236(.A(G244), .B(new_n260), .C1(new_n251), .C2(new_n252), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT4), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n259), .A2(G250), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT4), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G1698), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n268), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT74), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n275), .A2(G45), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G41), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT74), .A3(new_n275), .A4(G45), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(G257), .A3(new_n268), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n448), .A2(new_n452), .A3(G274), .A4(new_n449), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n269), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(G200), .B1(new_n444), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT75), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n456), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n438), .B1(new_n253), .B2(new_n220), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n434), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n260), .B1(new_n441), .B2(KEYINPUT4), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n269), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(G190), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n343), .A2(G97), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n256), .A2(G1), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n344), .A2(new_n209), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT73), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT6), .A2(G97), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(G107), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n213), .A2(KEYINPUT73), .A3(KEYINPUT6), .A4(G97), .ZN(new_n473));
  XOR2_X1   g0273(.A(G97), .B(G107), .Z(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(KEYINPUT6), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G20), .ZN(new_n476));
  OAI21_X1  g0276(.A(G107), .B1(new_n389), .B2(new_n390), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n293), .A2(G77), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n467), .B(new_n469), .C1(new_n479), .C2(new_n287), .ZN(new_n480));
  OAI211_X1 g0280(.A(KEYINPUT75), .B(G200), .C1(new_n444), .C2(new_n456), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n459), .A2(new_n466), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n469), .B1(new_n479), .B2(new_n287), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(G97), .B2(new_n343), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n455), .A2(new_n269), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n465), .A2(new_n486), .A3(new_n454), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n330), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n460), .A2(new_n271), .A3(new_n465), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n259), .A2(new_n227), .A3(G68), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n207), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n322), .A2(new_n227), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(KEYINPUT19), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT19), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n322), .B2(G20), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n491), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n287), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n344), .A2(new_n468), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n360), .A2(new_n284), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G238), .B(new_n260), .C1(new_n251), .C2(new_n252), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT76), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT76), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n259), .A2(new_n506), .A3(G238), .A4(new_n260), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n259), .A2(G244), .A3(G1698), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n505), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n269), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n447), .A2(new_n208), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n275), .A2(new_n303), .A3(G45), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n268), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n503), .B1(new_n515), .B2(G200), .ZN(new_n516));
  INV_X1    g0316(.A(new_n514), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n510), .B2(new_n269), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n498), .A2(new_n287), .B1(new_n284), .B2(new_n360), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n500), .A2(new_n359), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n518), .A2(new_n271), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n515), .A2(new_n330), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n516), .A2(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n482), .A2(new_n490), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT25), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n343), .B2(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n500), .A2(G107), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT23), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(G20), .B2(new_n213), .ZN(new_n532));
  INV_X1    g0332(.A(G116), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n291), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n213), .A3(G20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT81), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n227), .A2(G107), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT81), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(new_n531), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n532), .B(new_n534), .C1(new_n536), .C2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT82), .ZN(new_n542));
  AND2_X1   g0342(.A1(KEYINPUT80), .A2(G87), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n227), .B(new_n543), .C1(new_n251), .C2(new_n252), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n259), .A2(KEYINPUT22), .A3(new_n227), .A4(new_n543), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n540), .A2(new_n542), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n542), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n539), .A2(new_n536), .ZN(new_n550));
  INV_X1    g0350(.A(new_n534), .ZN(new_n551));
  INV_X1    g0351(.A(new_n532), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n546), .A2(new_n547), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n541), .A2(KEYINPUT82), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n530), .B1(new_n559), .B2(new_n287), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n453), .A2(G264), .A3(new_n268), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n251), .A2(new_n252), .B1(G250), .B2(G1698), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n260), .A2(G257), .ZN(new_n563));
  INV_X1    g0363(.A(G294), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n562), .A2(new_n563), .B1(new_n256), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n269), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n486), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n330), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n561), .A2(new_n566), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n485), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n271), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n567), .A2(G190), .A3(new_n486), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n557), .B1(new_n548), .B2(new_n555), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n529), .B(new_n574), .C1(new_n575), .C2(new_n300), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n571), .A2(new_n356), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n560), .A2(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n525), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n453), .A2(new_n268), .ZN(new_n580));
  OAI22_X1  g0380(.A1(new_n580), .A2(new_n240), .B1(new_n269), .B2(new_n455), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n260), .A2(G264), .ZN(new_n583));
  NOR2_X1   g0383(.A1(G257), .A2(G1698), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n583), .A2(new_n584), .B1(new_n251), .B2(new_n252), .ZN(new_n585));
  INV_X1    g0385(.A(G303), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n257), .A2(new_n586), .A3(new_n258), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n585), .A2(KEYINPUT77), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT77), .B1(new_n585), .B2(new_n587), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT78), .B1(new_n590), .B2(new_n269), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n214), .A2(G1698), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n210), .A2(new_n260), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n593), .A2(new_n594), .B1(new_n257), .B2(new_n258), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n251), .A2(new_n252), .A3(G303), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n585), .A2(KEYINPUT77), .A3(new_n587), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n597), .A2(KEYINPUT78), .A3(new_n269), .A4(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n582), .B1(new_n591), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n286), .A2(new_n226), .B1(G20), .B2(new_n533), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n434), .B(new_n227), .C1(G33), .C2(new_n209), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT20), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n284), .A2(new_n533), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n468), .B1(new_n346), .B2(new_n347), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G116), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n330), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n601), .A2(KEYINPUT21), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n597), .A2(new_n269), .A3(new_n598), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT78), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n581), .B1(new_n619), .B2(new_n599), .ZN(new_n620));
  AOI211_X1 g0420(.A(new_n533), .B(new_n468), .C1(new_n346), .C2(new_n347), .ZN(new_n621));
  OAI21_X1  g0421(.A(G169), .B1(new_n621), .B2(new_n610), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n616), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n611), .A2(new_n613), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(G179), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n615), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT79), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n619), .A2(new_n599), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(G190), .A3(new_n582), .ZN(new_n629));
  INV_X1    g0429(.A(new_n624), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n620), .A2(new_n356), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n627), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n601), .A2(G200), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(KEYINPUT79), .A3(new_n630), .A4(new_n629), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n626), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n433), .A2(new_n579), .A3(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n416), .ZN(new_n638));
  INV_X1    g0438(.A(new_n431), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n357), .B1(new_n336), .B2(new_n353), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n424), .A2(new_n428), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n638), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n315), .A2(new_n318), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n307), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n433), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n522), .A2(new_n523), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT83), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n516), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n516), .A2(new_n648), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n519), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n490), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n576), .A2(new_n577), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n656), .A3(new_n482), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n560), .A2(new_n573), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n626), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n654), .B(new_n655), .C1(new_n657), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n516), .A2(new_n519), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n653), .A2(KEYINPUT26), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n647), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n645), .B1(new_n646), .B2(new_n663), .ZN(G369));
  NOR3_X1   g0464(.A1(new_n283), .A2(G1), .A3(G20), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT84), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT27), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G213), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n665), .B2(new_n667), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n630), .A2(new_n675), .ZN(new_n676));
  MUX2_X1   g0476(.A(new_n636), .B(new_n626), .S(new_n676), .Z(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G330), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT85), .Z(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n560), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n578), .B1(new_n681), .B2(new_n674), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT86), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n658), .A2(new_n674), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(KEYINPUT86), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT87), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n680), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n658), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n674), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n626), .A2(new_n675), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n691), .A2(new_n696), .ZN(G399));
  NAND2_X1  g0497(.A1(new_n204), .A2(new_n272), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G1), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n492), .A2(new_n207), .A3(new_n533), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(new_n231), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g0501(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n702));
  XNOR2_X1  g0502(.A(new_n701), .B(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(G179), .B1(new_n628), .B2(new_n582), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(new_n568), .A3(new_n487), .A4(new_n515), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n567), .A2(new_n518), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n487), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(KEYINPUT30), .A3(G179), .A4(new_n620), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n628), .A2(G179), .A3(new_n582), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n460), .A2(new_n567), .A3(new_n465), .A4(new_n518), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n705), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n713), .A2(new_n714), .A3(new_n674), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n713), .B2(new_n674), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n579), .A2(new_n636), .A3(new_n675), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT89), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n720), .A2(new_n721), .A3(G330), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n720), .B2(G330), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n653), .A2(new_n655), .A3(new_n661), .ZN(new_n725));
  INV_X1    g0525(.A(new_n647), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n725), .B(new_n726), .C1(new_n655), .C2(new_n652), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n655), .B1(new_n657), .B2(new_n659), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(new_n490), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT29), .B1(new_n729), .B2(new_n674), .ZN(new_n730));
  OR3_X1    g0530(.A1(new_n663), .A2(KEYINPUT29), .A3(new_n674), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n724), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n703), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n677), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n226), .B1(G20), .B2(new_n330), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  NAND3_X1  g0541(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT94), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n350), .ZN(new_n746));
  INV_X1    g0546(.A(G190), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n227), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n356), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G87), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n227), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n749), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n752), .B(new_n259), .C1(new_n213), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT97), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n743), .A2(new_n747), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n755), .A2(new_n756), .B1(G50), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n271), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n748), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n753), .A2(new_n759), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G58), .A2(new_n761), .B1(new_n763), .B2(G77), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n758), .B1(KEYINPUT93), .B2(new_n764), .C1(new_n756), .C2(new_n755), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n746), .B(new_n765), .C1(KEYINPUT93), .C2(new_n764), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n753), .B1(new_n768), .B2(G20), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(KEYINPUT98), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(KEYINPUT98), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G97), .ZN(new_n774));
  INV_X1    g0574(.A(new_n753), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n778));
  XNOR2_X1  g0578(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n766), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT99), .ZN(new_n781));
  INV_X1    g0581(.A(new_n754), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n776), .A2(G329), .B1(G283), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G322), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT33), .B(G317), .Z(new_n785));
  OAI221_X1 g0585(.A(new_n783), .B1(new_n784), .B2(new_n760), .C1(new_n745), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G311), .B2(new_n763), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n259), .B1(new_n757), .B2(G326), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n586), .C2(new_n750), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G294), .B2(new_n773), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n741), .B1(new_n781), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n283), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n699), .B1(G45), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n259), .A2(new_n204), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT90), .Z(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G355), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n253), .A2(new_n204), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT91), .Z(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n231), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n249), .A2(new_n273), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n797), .B1(G116), .B2(new_n204), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n741), .A2(new_n737), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n794), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n739), .B1(new_n805), .B2(KEYINPUT100), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(KEYINPUT100), .B2(new_n805), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT101), .Z(new_n808));
  OAI211_X1 g0608(.A(new_n679), .B(new_n794), .C1(G330), .C2(new_n677), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(G396));
  NOR2_X1   g0610(.A1(new_n754), .A2(new_n350), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n253), .B(new_n811), .C1(G50), .C2(new_n751), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  INV_X1    g0613(.A(new_n776), .ZN(new_n814));
  INV_X1    g0614(.A(new_n773), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n812), .B1(new_n813), .B2(new_n814), .C1(new_n815), .C2(new_n383), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT102), .Z(new_n817));
  AOI22_X1  g0617(.A1(new_n744), .A2(G150), .B1(G143), .B2(new_n761), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n762), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G137), .B2(new_n757), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT34), .Z(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n757), .A2(G303), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n761), .A2(G294), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n782), .A2(G87), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G283), .B2(new_n744), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n774), .A2(new_n825), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n762), .A2(new_n533), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n750), .A2(new_n213), .ZN(new_n833));
  NOR4_X1   g0633(.A1(new_n831), .A2(new_n259), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n741), .B1(new_n824), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n741), .A2(new_n735), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n219), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n373), .A2(new_n330), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n840), .A2(new_n364), .A3(new_n430), .A4(new_n675), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n364), .A2(new_n674), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n370), .B2(new_n374), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(new_n843), .B2(new_n639), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n736), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n836), .A2(new_n794), .A3(new_n839), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n724), .A2(new_n844), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n722), .B2(new_n723), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n663), .A2(new_n674), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n850), .B(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n847), .B1(new_n852), .B2(new_n794), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n579), .A2(new_n636), .A3(new_n675), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT106), .B1(new_n717), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT106), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n719), .B(new_n858), .C1(new_n716), .C2(new_n715), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n353), .A2(new_n674), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n354), .A2(new_n357), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n336), .A2(new_n353), .A3(new_n674), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n844), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n857), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n422), .A2(new_n423), .A3(new_n417), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT72), .B1(new_n426), .B2(new_n427), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n638), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n672), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n398), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n398), .A2(new_n412), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT104), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n872), .A2(new_n869), .A3(new_n420), .A4(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n877), .B(KEYINPUT38), .C1(new_n429), .C2(new_n869), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n855), .B1(new_n864), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n420), .B(KEYINPUT17), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT105), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n416), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT105), .B1(new_n422), .B2(new_n423), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n869), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n875), .B(new_n876), .Z(new_n889));
  OAI21_X1  g0689(.A(new_n883), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n855), .B1(new_n890), .B2(new_n879), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n891), .A2(new_n857), .A3(new_n859), .A4(new_n863), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT107), .Z(new_n894));
  AND2_X1   g0694(.A1(new_n857), .A2(new_n859), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n433), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n894), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(G330), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n881), .A2(KEYINPUT39), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n890), .A2(new_n879), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n354), .A2(new_n674), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n861), .A2(new_n862), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n663), .A2(new_n674), .A3(new_n844), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n841), .B(KEYINPUT103), .Z(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n909), .A2(new_n881), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n416), .A2(new_n672), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n731), .A2(new_n730), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n433), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n645), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n912), .B(new_n915), .Z(new_n916));
  XNOR2_X1  g0716(.A(new_n898), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n275), .B2(new_n792), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n533), .B1(new_n475), .B2(KEYINPUT35), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n228), .C1(KEYINPUT35), .C2(new_n475), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT36), .ZN(new_n921));
  OAI21_X1  g0721(.A(G77), .B1(new_n383), .B2(new_n350), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n231), .A2(new_n922), .B1(G50), .B2(new_n350), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(G1), .A3(new_n283), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n918), .A2(new_n921), .A3(new_n924), .ZN(G367));
  NAND2_X1  g0725(.A1(new_n690), .A2(new_n695), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n482), .B(new_n490), .C1(new_n480), .C2(new_n675), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n653), .A2(new_n674), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT42), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n490), .B1(new_n927), .B2(new_n692), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n675), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n694), .B1(new_n688), .B2(new_n689), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT42), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n934), .A2(new_n935), .A3(new_n929), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n931), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n652), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n503), .A2(new_n674), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n726), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n726), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT43), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n942), .A3(new_n941), .ZN(new_n945));
  INV_X1    g0745(.A(new_n691), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n929), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n941), .A2(new_n942), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n937), .A2(new_n949), .A3(new_n943), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n945), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n948), .B1(new_n945), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n698), .B(KEYINPUT41), .Z(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n696), .A2(new_n929), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR4_X1   g0758(.A1(new_n934), .A2(new_n957), .A3(new_n693), .A4(new_n930), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT44), .B1(new_n696), .B2(new_n929), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT44), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(new_n930), .C1(new_n934), .C2(new_n693), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n961), .A2(new_n691), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n688), .A2(new_n689), .A3(new_n694), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n926), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(new_n679), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n732), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT45), .B1(new_n696), .B2(new_n929), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n959), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n962), .A2(new_n964), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n946), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n965), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n955), .B1(new_n974), .B2(new_n733), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n792), .A2(G45), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(G1), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT108), .Z(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n953), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n253), .B1(new_n757), .B2(G143), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n383), .B2(new_n750), .C1(new_n219), .C2(new_n754), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n773), .A2(G68), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n292), .B2(new_n760), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT110), .Z(new_n985));
  AOI211_X1 g0785(.A(new_n982), .B(new_n985), .C1(G50), .C2(new_n763), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n819), .B2(new_n745), .ZN(new_n987));
  XNOR2_X1  g0787(.A(KEYINPUT111), .B(G137), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n987), .B1(new_n776), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT112), .Z(new_n990));
  AOI21_X1  g0790(.A(new_n259), .B1(new_n757), .B2(G311), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n776), .A2(G317), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT46), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n750), .B2(new_n533), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n751), .A2(KEYINPUT46), .A3(G116), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n745), .C2(new_n564), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n991), .B(new_n992), .C1(new_n996), .C2(KEYINPUT109), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n815), .B2(new_n213), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(G303), .C2(new_n761), .ZN(new_n1000));
  INV_X1    g0800(.A(G283), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n209), .B2(new_n754), .C1(new_n1001), .C2(new_n762), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n990), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n741), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n941), .A2(new_n737), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n799), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n803), .B1(new_n204), .B2(new_n360), .C1(new_n241), .C2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1005), .A2(new_n793), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n980), .A2(new_n1009), .ZN(G387));
  AOI21_X1  g0810(.A(new_n698), .B1(new_n968), .B2(new_n732), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n969), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1007), .B1(new_n237), .B2(G45), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n700), .B2(new_n796), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n290), .A2(G50), .ZN(new_n1016));
  XOR2_X1   g0816(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n350), .A2(new_n219), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n1018), .A2(G45), .A3(new_n1019), .A4(new_n700), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1015), .A2(new_n1020), .B1(G107), .B2(new_n204), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n794), .B1(new_n1021), .B2(new_n803), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n690), .B2(new_n738), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n773), .A2(new_n359), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n350), .B2(new_n762), .C1(new_n292), .C2(new_n814), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n745), .A2(new_n290), .B1(new_n209), .B2(new_n754), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n253), .B1(new_n761), .B2(G50), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n757), .A2(G159), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n751), .A2(G77), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n744), .A2(G311), .B1(G317), .B2(new_n761), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n757), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n586), .B2(new_n762), .C1(new_n784), .C2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT48), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n1001), .B2(new_n815), .C1(new_n564), .C2(new_n750), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT49), .Z(new_n1037));
  AOI21_X1  g0837(.A(new_n259), .B1(new_n776), .B2(G326), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n533), .B2(new_n754), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1031), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1023), .B1(new_n741), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n968), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n979), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1013), .A2(new_n1043), .ZN(G393));
  NAND3_X1  g0844(.A1(new_n965), .A2(new_n973), .A3(new_n979), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n757), .A2(G150), .B1(G159), .B2(new_n761), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n773), .A2(G77), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n217), .B2(new_n745), .C1(new_n290), .C2(new_n762), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT114), .Z(new_n1050));
  AOI211_X1 g0850(.A(new_n253), .B(new_n1050), .C1(G68), .C2(new_n751), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n827), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1047), .B(new_n1052), .C1(G143), .C2(new_n776), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n757), .A2(G317), .B1(G311), .B2(new_n761), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G283), .B2(new_n751), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n213), .A2(new_n754), .B1(new_n762), .B2(new_n564), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n259), .B(new_n1057), .C1(new_n744), .C2(G303), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(new_n533), .C2(new_n815), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G322), .B2(new_n776), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n741), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n930), .A2(new_n737), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n803), .B1(new_n209), .B2(new_n204), .C1(new_n246), .C2(new_n1007), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1061), .A2(new_n793), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1045), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n965), .A2(new_n973), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n698), .B1(new_n1066), .B2(new_n1012), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1065), .B1(new_n1067), .B2(new_n974), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(G390));
  AND3_X1   g0869(.A1(new_n857), .A2(G330), .A3(new_n859), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n845), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n906), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n845), .B(new_n906), .C1(new_n722), .C2(new_n723), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n843), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n431), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n728), .A2(new_n490), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n675), .B(new_n1076), .C1(new_n1077), .C2(new_n727), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(new_n841), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1073), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1070), .A2(new_n863), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n849), .B2(new_n1072), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n907), .A2(new_n908), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n895), .A2(G330), .A3(new_n433), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n914), .A2(new_n645), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n904), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n900), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1078), .A2(new_n841), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n906), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n909), .A2(new_n1090), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1074), .C1(new_n1095), .C2(new_n903), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n909), .A2(new_n1090), .B1(new_n902), .B2(new_n899), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1082), .B1(new_n1097), .B2(new_n1093), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1089), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n698), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1089), .A2(new_n1099), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1096), .A2(new_n1098), .A3(new_n979), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n751), .A2(G150), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT53), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n259), .B1(new_n815), .B2(new_n819), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n744), .C2(new_n988), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n757), .A2(G128), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n776), .A2(G125), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n760), .A2(new_n813), .B1(new_n754), .B2(new_n217), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n763), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n253), .B1(new_n745), .B2(new_n213), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1048), .B1(new_n533), .B2(new_n760), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT116), .Z(new_n1117));
  AOI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(G294), .C2(new_n776), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n757), .A2(G283), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n763), .A2(G97), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1118), .A2(new_n752), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1114), .B1(new_n1121), .B2(new_n811), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n741), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n794), .B1(new_n837), .B2(new_n290), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT115), .Z(new_n1125));
  OAI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(new_n736), .C2(new_n903), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1104), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(KEYINPUT117), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1103), .B1(new_n1128), .B2(new_n1129), .ZN(G378));
  NAND2_X1  g0930(.A1(new_n849), .A2(new_n1072), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1084), .B1(new_n1131), .B2(new_n1081), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1080), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1088), .B1(new_n1134), .B2(new_n1099), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n644), .A2(new_n306), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1137), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n319), .A2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1138), .A2(new_n1140), .B1(new_n301), .B2(new_n868), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n319), .A2(new_n1139), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n307), .B(new_n1137), .C1(new_n315), .C2(new_n318), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n301), .A2(new_n868), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n882), .A2(G330), .A3(new_n892), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(KEYINPUT120), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT121), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT120), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n882), .A2(new_n1150), .A3(new_n892), .A4(G330), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n882), .A2(G330), .A3(new_n892), .A4(new_n1146), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT121), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n912), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1152), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1147), .A2(KEYINPUT120), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1146), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1151), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1154), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n912), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(KEYINPUT57), .B(new_n1135), .C1(new_n1157), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT122), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1135), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1156), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1162), .A2(new_n912), .A3(new_n1163), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1173), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n1135), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1167), .A2(new_n1170), .A3(new_n1101), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n978), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n773), .A2(G150), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n744), .A2(G132), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n757), .A2(G125), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G128), .A2(new_n761), .B1(new_n763), .B2(G137), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n751), .B2(new_n1112), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT59), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G41), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT118), .B(G124), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1184), .B1(new_n814), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1186), .A2(G33), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n1183), .B2(new_n1182), .C1(new_n819), .C2(new_n754), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n744), .A2(G97), .B1(G77), .B2(new_n751), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n983), .B(new_n1189), .C1(new_n1001), .C2(new_n814), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n253), .B1(new_n1033), .B2(new_n533), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n754), .A2(new_n383), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1190), .A2(G41), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n213), .B2(new_n760), .C1(new_n360), .C2(new_n762), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT58), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n217), .B1(new_n251), .B2(G41), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT119), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n741), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1159), .A2(new_n735), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n837), .A2(new_n217), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1199), .A2(new_n793), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1176), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1175), .A2(new_n1204), .ZN(G375));
  OAI211_X1 g1005(.A(new_n1080), .B(new_n1087), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1089), .A2(new_n954), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1072), .A2(new_n735), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n744), .A2(new_n1112), .B1(new_n761), .B2(new_n988), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n813), .B2(new_n1033), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT123), .Z(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G150), .B2(new_n763), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n253), .B(new_n1192), .C1(G159), .C2(new_n751), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n217), .C2(new_n815), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G128), .B2(new_n776), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n750), .A2(new_n209), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n763), .A2(G107), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n776), .A2(G303), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n760), .A2(new_n1001), .B1(new_n754), .B2(new_n219), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n259), .B(new_n1219), .C1(new_n757), .C2(G294), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1024), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1216), .B(new_n1221), .C1(G116), .C2(new_n744), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n741), .B1(new_n1215), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n837), .A2(new_n350), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1208), .A2(new_n1223), .A3(new_n793), .A4(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1134), .B2(new_n978), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1207), .A2(new_n1227), .ZN(G381));
  AND3_X1   g1028(.A1(new_n1103), .A2(new_n1104), .A3(new_n1126), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1175), .A2(new_n1204), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n853), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(G381), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n980), .A2(new_n1009), .A3(new_n1068), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(G407));
  AOI21_X1  g1035(.A(new_n669), .B1(new_n1230), .B2(new_n673), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G407), .A2(new_n1236), .ZN(G409));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(G2897), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n669), .A2(G343), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(G2897), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1175), .A2(G378), .A3(new_n1204), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1173), .A2(new_n979), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(KEYINPUT124), .A3(new_n1202), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1173), .A2(new_n954), .A3(new_n1135), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT124), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1176), .B2(new_n1203), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1229), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1240), .B1(new_n1243), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  OR3_X1    g1052(.A1(new_n1206), .A2(KEYINPUT125), .A3(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT125), .B1(new_n1206), .B2(new_n1252), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n698), .B1(new_n1206), .B2(new_n1252), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1256), .A2(new_n1089), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1258), .B2(new_n1227), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1226), .B(new_n853), .C1(new_n1255), .C2(new_n1257), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1242), .B1(new_n1251), .B2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G2897), .B(new_n1240), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT127), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1263), .B(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1251), .A2(new_n1261), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1251), .A2(new_n1270), .A3(new_n1261), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .A4(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(G393), .A2(G396), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(new_n1234), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1068), .B1(new_n980), .B2(new_n1009), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1233), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(G390), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n980), .A2(new_n1009), .A3(new_n1068), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1273), .A2(new_n1234), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1272), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1268), .B2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1251), .A2(KEYINPUT63), .A3(new_n1261), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1284), .A2(new_n1267), .A3(new_n1266), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1229), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1288), .A2(new_n1243), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1281), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1281), .A2(new_n1289), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1261), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1290), .A2(new_n1261), .A3(new_n1291), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G402));
endmodule


