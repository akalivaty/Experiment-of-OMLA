

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(n713), .B(n712), .ZN(n715) );
  AND2_X1 U556 ( .A1(n998), .A2(n837), .ZN(n523) );
  NOR2_X1 U557 ( .A1(n826), .A2(n523), .ZN(n524) );
  AND2_X1 U558 ( .A1(n772), .A2(n976), .ZN(n525) );
  INV_X1 U559 ( .A(KEYINPUT26), .ZN(n718) );
  INV_X1 U560 ( .A(KEYINPUT27), .ZN(n711) );
  XNOR2_X1 U561 ( .A(n711), .B(KEYINPUT99), .ZN(n712) );
  OR2_X1 U562 ( .A1(n728), .A2(n729), .ZN(n727) );
  INV_X1 U563 ( .A(n745), .ZN(n740) );
  NAND2_X1 U564 ( .A1(n744), .A2(n743), .ZN(n759) );
  NAND2_X1 U565 ( .A1(n794), .A2(n704), .ZN(n745) );
  INV_X1 U566 ( .A(n787), .ZN(n773) );
  XOR2_X1 U567 ( .A(KEYINPUT65), .B(n541), .Z(n652) );
  NOR2_X2 U568 ( .A1(G2104), .A2(n555), .ZN(n882) );
  NOR2_X1 U569 ( .A1(G651), .A2(n666), .ZN(n661) );
  XOR2_X1 U570 ( .A(G2430), .B(G2443), .Z(n527) );
  XNOR2_X1 U571 ( .A(KEYINPUT105), .B(G2451), .ZN(n526) );
  XNOR2_X1 U572 ( .A(n527), .B(n526), .ZN(n534) );
  XOR2_X1 U573 ( .A(G2435), .B(G2427), .Z(n529) );
  XNOR2_X1 U574 ( .A(G2446), .B(G2454), .ZN(n528) );
  XNOR2_X1 U575 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U576 ( .A(n530), .B(G2438), .Z(n532) );
  XNOR2_X1 U577 ( .A(G1348), .B(G1341), .ZN(n531) );
  XNOR2_X1 U578 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U579 ( .A(n534), .B(n533), .ZN(n535) );
  AND2_X1 U580 ( .A1(n535), .A2(G14), .ZN(G401) );
  INV_X1 U581 ( .A(G651), .ZN(n540) );
  NOR2_X1 U582 ( .A1(G543), .A2(n540), .ZN(n537) );
  XNOR2_X1 U583 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n536) );
  XNOR2_X1 U584 ( .A(n537), .B(n536), .ZN(n665) );
  NAND2_X1 U585 ( .A1(G64), .A2(n665), .ZN(n539) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n666) );
  NAND2_X1 U587 ( .A1(G52), .A2(n661), .ZN(n538) );
  NAND2_X1 U588 ( .A1(n539), .A2(n538), .ZN(n547) );
  NOR2_X1 U589 ( .A1(n666), .A2(n540), .ZN(n650) );
  NAND2_X1 U590 ( .A1(G77), .A2(n650), .ZN(n543) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G90), .A2(n652), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U594 ( .A(KEYINPUT70), .B(n544), .Z(n545) );
  XNOR2_X1 U595 ( .A(KEYINPUT9), .B(n545), .ZN(n546) );
  NOR2_X1 U596 ( .A1(n547), .A2(n546), .ZN(G171) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  NOR2_X1 U598 ( .A1(G2104), .A2(G2105), .ZN(n548) );
  XOR2_X2 U599 ( .A(KEYINPUT17), .B(n548), .Z(n878) );
  NAND2_X1 U600 ( .A1(G135), .A2(n878), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G2105), .A2(G2104), .ZN(n549) );
  XOR2_X1 U602 ( .A(KEYINPUT66), .B(n549), .Z(n883) );
  NAND2_X1 U603 ( .A1(G111), .A2(n883), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n554) );
  INV_X1 U605 ( .A(G2105), .ZN(n555) );
  NAND2_X1 U606 ( .A1(n882), .A2(G123), .ZN(n552) );
  XOR2_X1 U607 ( .A(KEYINPUT18), .B(n552), .Z(n553) );
  NOR2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n557) );
  AND2_X1 U609 ( .A1(n555), .A2(G2104), .ZN(n879) );
  NAND2_X1 U610 ( .A1(n879), .A2(G99), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n946) );
  XNOR2_X1 U612 ( .A(G2096), .B(n946), .ZN(n558) );
  OR2_X1 U613 ( .A1(G2100), .A2(n558), .ZN(G156) );
  INV_X1 U614 ( .A(G108), .ZN(G238) );
  INV_X1 U615 ( .A(G120), .ZN(G236) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  NAND2_X1 U618 ( .A1(G75), .A2(n650), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G88), .A2(n652), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U621 ( .A1(G62), .A2(n665), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G50), .A2(n661), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(G166) );
  NAND2_X1 U625 ( .A1(n879), .A2(G102), .ZN(n571) );
  NAND2_X1 U626 ( .A1(G126), .A2(n882), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT90), .B(n565), .Z(n569) );
  NAND2_X1 U628 ( .A1(G138), .A2(n878), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G114), .A2(n883), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U633 ( .A(n572), .B(KEYINPUT91), .ZN(G164) );
  NAND2_X1 U634 ( .A1(G89), .A2(n652), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT79), .B(n573), .Z(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT4), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G76), .A2(n650), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U639 ( .A(n577), .B(KEYINPUT5), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G63), .A2(n665), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G51), .A2(n661), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT6), .B(n580), .Z(n581) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U645 ( .A(n583), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U646 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G567), .ZN(n692) );
  NOR2_X1 U650 ( .A1(G223), .A2(n692), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n585), .Z(n586) );
  XNOR2_X1 U652 ( .A(KEYINPUT73), .B(n586), .ZN(G234) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n588) );
  NAND2_X1 U654 ( .A1(G56), .A2(n665), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n588), .B(n587), .ZN(n602) );
  NAND2_X1 U656 ( .A1(G81), .A2(n652), .ZN(n590) );
  XOR2_X1 U657 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n589) );
  XNOR2_X1 U658 ( .A(n590), .B(n589), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G68), .A2(n650), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U661 ( .A(n593), .B(KEYINPUT13), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n594), .A2(KEYINPUT76), .ZN(n598) );
  INV_X1 U663 ( .A(n594), .ZN(n596) );
  INV_X1 U664 ( .A(KEYINPUT76), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G43), .A2(n661), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X2 U669 ( .A1(n602), .A2(n601), .ZN(n978) );
  NAND2_X1 U670 ( .A1(G860), .A2(n978), .ZN(n603) );
  XOR2_X1 U671 ( .A(KEYINPUT77), .B(n603), .Z(G153) );
  INV_X1 U672 ( .A(G171), .ZN(G301) );
  NAND2_X1 U673 ( .A1(G868), .A2(G301), .ZN(n613) );
  NAND2_X1 U674 ( .A1(n661), .A2(G54), .ZN(n610) );
  NAND2_X1 U675 ( .A1(G66), .A2(n665), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G79), .A2(n650), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U678 ( .A1(n652), .A2(G92), .ZN(n606) );
  XOR2_X1 U679 ( .A(KEYINPUT78), .B(n606), .Z(n607) );
  NOR2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U682 ( .A(KEYINPUT15), .B(n611), .Z(n728) );
  INV_X1 U683 ( .A(G868), .ZN(n679) );
  NAND2_X1 U684 ( .A1(n728), .A2(n679), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(G284) );
  NAND2_X1 U686 ( .A1(G65), .A2(n665), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G91), .A2(n652), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G78), .A2(n650), .ZN(n616) );
  XNOR2_X1 U690 ( .A(KEYINPUT71), .B(n616), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n661), .A2(G53), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(G299) );
  NOR2_X1 U694 ( .A1(G286), .A2(n679), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT80), .ZN(n623) );
  NOR2_X1 U696 ( .A1(G299), .A2(G868), .ZN(n622) );
  NOR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(G297) );
  INV_X1 U698 ( .A(G860), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n624), .A2(G559), .ZN(n625) );
  INV_X1 U700 ( .A(n728), .ZN(n989) );
  NAND2_X1 U701 ( .A1(n625), .A2(n989), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n626), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U703 ( .A1(n728), .A2(n679), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n627), .B(KEYINPUT81), .ZN(n628) );
  NOR2_X1 U705 ( .A1(G559), .A2(n628), .ZN(n630) );
  AND2_X1 U706 ( .A1(n679), .A2(n978), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n630), .A2(n629), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G559), .A2(n989), .ZN(n631) );
  XOR2_X1 U709 ( .A(n978), .B(n631), .Z(n675) );
  NOR2_X1 U710 ( .A1(n675), .A2(G860), .ZN(n641) );
  NAND2_X1 U711 ( .A1(G93), .A2(n652), .ZN(n632) );
  XNOR2_X1 U712 ( .A(n632), .B(KEYINPUT82), .ZN(n637) );
  NAND2_X1 U713 ( .A1(G67), .A2(n665), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G55), .A2(n661), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U716 ( .A(KEYINPUT84), .B(n635), .Z(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U718 ( .A1(G80), .A2(n650), .ZN(n638) );
  XNOR2_X1 U719 ( .A(KEYINPUT83), .B(n638), .ZN(n639) );
  OR2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n678) );
  XOR2_X1 U721 ( .A(n641), .B(n678), .Z(G145) );
  NAND2_X1 U722 ( .A1(G72), .A2(n650), .ZN(n643) );
  NAND2_X1 U723 ( .A1(G85), .A2(n652), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n661), .A2(G47), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n665), .A2(G60), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U728 ( .A(KEYINPUT68), .B(n646), .ZN(n647) );
  NOR2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(KEYINPUT69), .ZN(G290) );
  NAND2_X1 U731 ( .A1(G73), .A2(n650), .ZN(n651) );
  XNOR2_X1 U732 ( .A(n651), .B(KEYINPUT2), .ZN(n659) );
  NAND2_X1 U733 ( .A1(G61), .A2(n665), .ZN(n654) );
  NAND2_X1 U734 ( .A1(G86), .A2(n652), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U736 ( .A1(G48), .A2(n661), .ZN(n655) );
  XNOR2_X1 U737 ( .A(KEYINPUT85), .B(n655), .ZN(n656) );
  NOR2_X1 U738 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(KEYINPUT86), .B(n660), .ZN(G305) );
  NAND2_X1 U741 ( .A1(G49), .A2(n661), .ZN(n663) );
  NAND2_X1 U742 ( .A1(G74), .A2(G651), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U745 ( .A1(n666), .A2(G87), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n668), .A2(n667), .ZN(G288) );
  XOR2_X1 U747 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n669) );
  XNOR2_X1 U748 ( .A(G288), .B(n669), .ZN(n670) );
  XNOR2_X1 U749 ( .A(n670), .B(n678), .ZN(n672) );
  INV_X1 U750 ( .A(G299), .ZN(n992) );
  XNOR2_X1 U751 ( .A(n992), .B(G166), .ZN(n671) );
  XNOR2_X1 U752 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U753 ( .A(G305), .B(n673), .Z(n674) );
  XNOR2_X1 U754 ( .A(G290), .B(n674), .ZN(n893) );
  XNOR2_X1 U755 ( .A(KEYINPUT88), .B(n675), .ZN(n676) );
  XNOR2_X1 U756 ( .A(n893), .B(n676), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n677), .A2(G868), .ZN(n681) );
  NAND2_X1 U758 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U759 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U760 ( .A1(G2084), .A2(G2078), .ZN(n682) );
  XOR2_X1 U761 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U766 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U767 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U768 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U769 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U770 ( .A1(G96), .A2(n688), .ZN(n846) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n846), .ZN(n689) );
  XNOR2_X1 U772 ( .A(n689), .B(KEYINPUT89), .ZN(n694) );
  NOR2_X1 U773 ( .A1(G236), .A2(G238), .ZN(n690) );
  NAND2_X1 U774 ( .A1(G69), .A2(n690), .ZN(n691) );
  NOR2_X1 U775 ( .A1(G237), .A2(n691), .ZN(n848) );
  NOR2_X1 U776 ( .A1(n692), .A2(n848), .ZN(n693) );
  NOR2_X1 U777 ( .A1(n694), .A2(n693), .ZN(G319) );
  INV_X1 U778 ( .A(G319), .ZN(n696) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n695) );
  NOR2_X1 U780 ( .A1(n696), .A2(n695), .ZN(n845) );
  NAND2_X1 U781 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U782 ( .A1(n878), .A2(G137), .ZN(n699) );
  NAND2_X1 U783 ( .A1(G101), .A2(n879), .ZN(n697) );
  XOR2_X1 U784 ( .A(KEYINPUT23), .B(n697), .Z(n698) );
  NAND2_X1 U785 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U786 ( .A1(G125), .A2(n882), .ZN(n701) );
  NAND2_X1 U787 ( .A1(G113), .A2(n883), .ZN(n700) );
  NAND2_X1 U788 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U789 ( .A1(n703), .A2(n702), .ZN(G160) );
  INV_X1 U790 ( .A(G166), .ZN(G303) );
  NOR2_X1 U791 ( .A1(G164), .A2(G1384), .ZN(n794) );
  NAND2_X1 U792 ( .A1(G160), .A2(G40), .ZN(n793) );
  INV_X1 U793 ( .A(n793), .ZN(n704) );
  NOR2_X1 U794 ( .A1(G2090), .A2(n745), .ZN(n705) );
  XNOR2_X1 U795 ( .A(KEYINPUT103), .B(n705), .ZN(n708) );
  NAND2_X1 U796 ( .A1(G8), .A2(n745), .ZN(n787) );
  NOR2_X1 U797 ( .A1(G1971), .A2(n787), .ZN(n706) );
  NOR2_X1 U798 ( .A1(G166), .A2(n706), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n753) );
  INV_X1 U800 ( .A(n753), .ZN(n709) );
  OR2_X1 U801 ( .A1(n709), .A2(G286), .ZN(n710) );
  AND2_X1 U802 ( .A1(G8), .A2(n710), .ZN(n756) );
  NAND2_X1 U803 ( .A1(G2072), .A2(n740), .ZN(n713) );
  AND2_X1 U804 ( .A1(n745), .A2(G1956), .ZN(n714) );
  NOR2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n992), .A2(n734), .ZN(n733) );
  NAND2_X1 U807 ( .A1(n745), .A2(G1341), .ZN(n716) );
  XNOR2_X1 U808 ( .A(n716), .B(KEYINPUT100), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n717), .A2(n978), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n740), .A2(G1996), .ZN(n719) );
  XNOR2_X1 U811 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n723) );
  INV_X1 U813 ( .A(KEYINPUT64), .ZN(n722) );
  XNOR2_X1 U814 ( .A(n723), .B(n722), .ZN(n729) );
  NOR2_X1 U815 ( .A1(n740), .A2(G1348), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G2067), .A2(n745), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n737) );
  NOR2_X1 U822 ( .A1(n992), .A2(n734), .ZN(n735) );
  XOR2_X1 U823 ( .A(n735), .B(KEYINPUT28), .Z(n736) );
  NAND2_X1 U824 ( .A1(n737), .A2(n736), .ZN(n739) );
  XNOR2_X1 U825 ( .A(KEYINPUT101), .B(KEYINPUT29), .ZN(n738) );
  XNOR2_X1 U826 ( .A(n739), .B(n738), .ZN(n744) );
  XOR2_X1 U827 ( .A(G1961), .B(KEYINPUT98), .Z(n1005) );
  NAND2_X1 U828 ( .A1(n1005), .A2(n745), .ZN(n742) );
  XNOR2_X1 U829 ( .A(KEYINPUT25), .B(G2078), .ZN(n927) );
  NAND2_X1 U830 ( .A1(n740), .A2(n927), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n749) );
  NAND2_X1 U832 ( .A1(n749), .A2(G171), .ZN(n743) );
  NOR2_X1 U833 ( .A1(G1966), .A2(n787), .ZN(n764) );
  NOR2_X1 U834 ( .A1(G2084), .A2(n745), .ZN(n761) );
  NOR2_X1 U835 ( .A1(n764), .A2(n761), .ZN(n746) );
  NAND2_X1 U836 ( .A1(G8), .A2(n746), .ZN(n747) );
  XNOR2_X1 U837 ( .A(KEYINPUT30), .B(n747), .ZN(n748) );
  NOR2_X1 U838 ( .A1(G168), .A2(n748), .ZN(n751) );
  NOR2_X1 U839 ( .A1(G171), .A2(n749), .ZN(n750) );
  NOR2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U841 ( .A(KEYINPUT31), .B(n752), .Z(n758) );
  AND2_X1 U842 ( .A1(n758), .A2(n753), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n759), .A2(n754), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U845 ( .A(n757), .B(KEYINPUT32), .ZN(n768) );
  NAND2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U847 ( .A(n760), .B(KEYINPUT102), .ZN(n766) );
  NAND2_X1 U848 ( .A1(n761), .A2(G8), .ZN(n762) );
  XNOR2_X1 U849 ( .A(KEYINPUT97), .B(n762), .ZN(n763) );
  NOR2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n768), .A2(n767), .ZN(n783) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n991) );
  NOR2_X1 U854 ( .A1(G1971), .A2(G303), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n991), .A2(n769), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n783), .A2(n770), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT104), .ZN(n772) );
  NAND2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NAND2_X1 U859 ( .A1(n525), .A2(n773), .ZN(n775) );
  INV_X1 U860 ( .A(KEYINPUT33), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n780) );
  NAND2_X1 U862 ( .A1(n991), .A2(KEYINPUT33), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n776), .A2(n787), .ZN(n778) );
  XOR2_X1 U864 ( .A(G305), .B(G1981), .Z(n984) );
  INV_X1 U865 ( .A(n984), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  AND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n791) );
  NOR2_X1 U868 ( .A1(G2090), .A2(G303), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G8), .A2(n781), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n784), .A2(n787), .ZN(n789) );
  NOR2_X1 U872 ( .A1(G305), .A2(G1981), .ZN(n785) );
  XOR2_X1 U873 ( .A(n785), .B(KEYINPUT24), .Z(n786) );
  OR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U876 ( .A1(n791), .A2(n790), .ZN(n792) );
  INV_X1 U877 ( .A(n792), .ZN(n827) );
  NOR2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n837) );
  NAND2_X1 U879 ( .A1(G140), .A2(n878), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G104), .A2(n879), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U882 ( .A(n797), .B(KEYINPUT93), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n798), .B(KEYINPUT34), .ZN(n804) );
  XNOR2_X1 U884 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n802) );
  NAND2_X1 U885 ( .A1(G128), .A2(n882), .ZN(n800) );
  NAND2_X1 U886 ( .A1(G116), .A2(n883), .ZN(n799) );
  NAND2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n802), .B(n801), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U890 ( .A(KEYINPUT36), .B(n805), .Z(n860) );
  XNOR2_X1 U891 ( .A(G2067), .B(KEYINPUT37), .ZN(n835) );
  NOR2_X1 U892 ( .A1(n860), .A2(n835), .ZN(n966) );
  NAND2_X1 U893 ( .A1(n837), .A2(n966), .ZN(n833) );
  NAND2_X1 U894 ( .A1(G131), .A2(n878), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G95), .A2(n879), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U897 ( .A(KEYINPUT95), .B(n808), .ZN(n812) );
  NAND2_X1 U898 ( .A1(n883), .A2(G107), .ZN(n810) );
  NAND2_X1 U899 ( .A1(G119), .A2(n882), .ZN(n809) );
  AND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n858) );
  AND2_X1 U902 ( .A1(n858), .A2(G1991), .ZN(n822) );
  NAND2_X1 U903 ( .A1(G129), .A2(n882), .ZN(n814) );
  NAND2_X1 U904 ( .A1(G117), .A2(n883), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n817) );
  NAND2_X1 U906 ( .A1(n879), .A2(G105), .ZN(n815) );
  XOR2_X1 U907 ( .A(KEYINPUT38), .B(n815), .Z(n816) );
  NOR2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U909 ( .A(n818), .B(KEYINPUT96), .ZN(n820) );
  NAND2_X1 U910 ( .A1(G141), .A2(n878), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n820), .A2(n819), .ZN(n859) );
  AND2_X1 U912 ( .A1(n859), .A2(G1996), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n963) );
  INV_X1 U914 ( .A(n837), .ZN(n823) );
  NOR2_X1 U915 ( .A1(n963), .A2(n823), .ZN(n830) );
  INV_X1 U916 ( .A(n830), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n833), .A2(n824), .ZN(n826) );
  XNOR2_X1 U918 ( .A(G1986), .B(KEYINPUT92), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(G290), .ZN(n998) );
  NAND2_X1 U920 ( .A1(n827), .A2(n524), .ZN(n840) );
  NOR2_X1 U921 ( .A1(G1996), .A2(n859), .ZN(n957) );
  NOR2_X1 U922 ( .A1(G1986), .A2(G290), .ZN(n828) );
  NOR2_X1 U923 ( .A1(G1991), .A2(n858), .ZN(n949) );
  NOR2_X1 U924 ( .A1(n828), .A2(n949), .ZN(n829) );
  NOR2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U926 ( .A1(n957), .A2(n831), .ZN(n832) );
  XNOR2_X1 U927 ( .A(n832), .B(KEYINPUT39), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n860), .A2(n835), .ZN(n950) );
  NAND2_X1 U930 ( .A1(n836), .A2(n950), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U933 ( .A(n841), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U934 ( .A(G223), .ZN(n842) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U939 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(n846), .ZN(n847) );
  NAND2_X1 U943 ( .A1(n848), .A2(n847), .ZN(G261) );
  INV_X1 U944 ( .A(G261), .ZN(G325) );
  NAND2_X1 U945 ( .A1(G124), .A2(n882), .ZN(n849) );
  XNOR2_X1 U946 ( .A(n849), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U947 ( .A1(n879), .A2(G100), .ZN(n851) );
  NAND2_X1 U948 ( .A1(G112), .A2(n883), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(KEYINPUT110), .B(n852), .Z(n853) );
  NAND2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G136), .A2(n878), .ZN(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(n855), .ZN(n856) );
  NOR2_X1 U954 ( .A1(n857), .A2(n856), .ZN(G162) );
  XOR2_X1 U955 ( .A(n858), .B(G162), .Z(n862) );
  XOR2_X1 U956 ( .A(n860), .B(n859), .Z(n861) );
  XNOR2_X1 U957 ( .A(n862), .B(n861), .ZN(n877) );
  NAND2_X1 U958 ( .A1(G130), .A2(n882), .ZN(n864) );
  NAND2_X1 U959 ( .A1(G118), .A2(n883), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n870) );
  NAND2_X1 U961 ( .A1(G142), .A2(n878), .ZN(n866) );
  NAND2_X1 U962 ( .A1(G106), .A2(n879), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U964 ( .A(KEYINPUT111), .B(n867), .ZN(n868) );
  XNOR2_X1 U965 ( .A(KEYINPUT45), .B(n868), .ZN(n869) );
  NOR2_X1 U966 ( .A1(n870), .A2(n869), .ZN(n874) );
  XOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n872) );
  XNOR2_X1 U968 ( .A(G160), .B(KEYINPUT113), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U970 ( .A(n874), .B(n873), .Z(n875) );
  XNOR2_X1 U971 ( .A(n946), .B(n875), .ZN(n876) );
  XOR2_X1 U972 ( .A(n877), .B(n876), .Z(n891) );
  NAND2_X1 U973 ( .A1(G139), .A2(n878), .ZN(n881) );
  NAND2_X1 U974 ( .A1(G103), .A2(n879), .ZN(n880) );
  NAND2_X1 U975 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U976 ( .A1(G127), .A2(n882), .ZN(n885) );
  NAND2_X1 U977 ( .A1(G115), .A2(n883), .ZN(n884) );
  NAND2_X1 U978 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n886), .Z(n887) );
  NOR2_X1 U980 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U981 ( .A(KEYINPUT112), .B(n889), .Z(n952) );
  XNOR2_X1 U982 ( .A(G164), .B(n952), .ZN(n890) );
  XNOR2_X1 U983 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U984 ( .A1(G37), .A2(n892), .ZN(G395) );
  XOR2_X1 U985 ( .A(n893), .B(G286), .Z(n895) );
  XNOR2_X1 U986 ( .A(n989), .B(G171), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U988 ( .A(n978), .B(n896), .Z(n897) );
  NOR2_X1 U989 ( .A1(G37), .A2(n897), .ZN(G397) );
  XNOR2_X1 U990 ( .A(G1991), .B(G2474), .ZN(n907) );
  XOR2_X1 U991 ( .A(G1976), .B(G1971), .Z(n899) );
  XNOR2_X1 U992 ( .A(G1996), .B(G1986), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U994 ( .A(G1981), .B(G1961), .Z(n901) );
  XNOR2_X1 U995 ( .A(G1966), .B(G1956), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U997 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U998 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(G229) );
  XOR2_X1 U1001 ( .A(KEYINPUT43), .B(G2678), .Z(n909) );
  XNOR2_X1 U1002 ( .A(KEYINPUT107), .B(KEYINPUT106), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1004 ( .A(KEYINPUT42), .B(G2090), .Z(n911) );
  XNOR2_X1 U1005 ( .A(G2067), .B(G2072), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1007 ( .A(n913), .B(n912), .Z(n915) );
  XNOR2_X1 U1008 ( .A(G2096), .B(G2100), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1010 ( .A(G2084), .B(G2078), .Z(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(G227) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n918) );
  XOR2_X1 U1013 ( .A(KEYINPUT115), .B(n918), .Z(n924) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n919) );
  XOR2_X1 U1015 ( .A(KEYINPUT49), .B(n919), .Z(n920) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n920), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT114), .B(n922), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1022 ( .A(G2090), .B(G35), .ZN(n938) );
  XOR2_X1 U1023 ( .A(G2067), .B(G26), .Z(n926) );
  XOR2_X1 U1024 ( .A(G1991), .B(G25), .Z(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n935) );
  XNOR2_X1 U1026 ( .A(G27), .B(n927), .ZN(n933) );
  XOR2_X1 U1027 ( .A(G32), .B(G1996), .Z(n928) );
  NAND2_X1 U1028 ( .A1(n928), .A2(G28), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G33), .B(G2072), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT118), .B(n929), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(KEYINPUT53), .B(n936), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n941) );
  XOR2_X1 U1036 ( .A(G2084), .B(G34), .Z(n939) );
  XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(n939), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1039 ( .A(KEYINPUT55), .B(n942), .Z(n943) );
  INV_X1 U1040 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n971), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(G11), .A2(n944), .ZN(n973) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(KEYINPUT117), .ZN(n968) );
  XNOR2_X1 U1044 ( .A(G160), .B(G2084), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(n945), .B(KEYINPUT116), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n962) );
  XOR2_X1 U1049 ( .A(G164), .B(G2078), .Z(n954) );
  XNOR2_X1 U1050 ( .A(G2072), .B(n952), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(KEYINPUT50), .B(n955), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G2090), .B(G162), .Z(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1055 ( .A(KEYINPUT51), .B(n958), .Z(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n968), .B(n967), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n969), .A2(KEYINPUT55), .ZN(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n1004) );
  XOR2_X1 U1064 ( .A(G16), .B(KEYINPUT119), .Z(n974) );
  XNOR2_X1 U1065 ( .A(KEYINPUT56), .B(n974), .ZN(n1002) );
  XNOR2_X1 U1066 ( .A(G1971), .B(G166), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n975), .B(KEYINPUT122), .ZN(n983) );
  XNOR2_X1 U1068 ( .A(G171), .B(G1961), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n978), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(KEYINPUT123), .B(n979), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n988) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n986), .Z(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n1000) );
  XNOR2_X1 U1078 ( .A(G1348), .B(n989), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(n990), .B(KEYINPUT120), .ZN(n996) );
  XOR2_X1 U1080 ( .A(n991), .B(KEYINPUT121), .Z(n994) );
  XOR2_X1 U1081 ( .A(n992), .B(G1956), .Z(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1086 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1087 ( .A1(n1004), .A2(n1003), .ZN(n1032) );
  XNOR2_X1 U1088 ( .A(n1005), .B(G5), .ZN(n1021) );
  XNOR2_X1 U1089 ( .A(G1956), .B(G20), .ZN(n1011) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(n1006), .B(KEYINPUT124), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1007) );
  NOR2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(KEYINPUT125), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1095 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(KEYINPUT126), .B(n1012), .ZN(n1015) );
  XNOR2_X1 U1097 ( .A(G1348), .B(KEYINPUT59), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1013), .B(G4), .ZN(n1014) );
  NAND2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(n1016), .B(KEYINPUT60), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(KEYINPUT127), .B(n1017), .Z(n1019) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1018) );
  NOR2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1104 ( .A1(n1021), .A2(n1020), .ZN(n1028) );
  XNOR2_X1 U1105 ( .A(G1971), .B(G22), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(G23), .B(G1976), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  XOR2_X1 U1108 ( .A(G1986), .B(G24), .Z(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(KEYINPUT58), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1029), .Z(n1030) );
  NOR2_X1 U1113 ( .A1(G16), .A2(n1030), .ZN(n1031) );
  NOR2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1115 ( .A(n1033), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

