//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT0), .A3(G128), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G134), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n201));
  AOI22_X1  g015(.A1(KEYINPUT65), .A2(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(new_n201), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n198), .B2(G134), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n202), .A2(new_n203), .A3(new_n208), .A4(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n201), .B1(new_n204), .B2(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(KEYINPUT65), .A3(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n200), .B1(new_n215), .B2(new_n201), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(KEYINPUT66), .B(G131), .C1(new_n214), .C2(new_n216), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT69), .B1(new_n219), .B2(new_n220), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n197), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G116), .B(G119), .ZN(new_n224));
  INV_X1    g038(.A(G113), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(KEYINPUT2), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n224), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G116), .ZN(new_n230));
  INV_X1    g044(.A(G116), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n239), .A2(new_n188), .A3(new_n190), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT68), .A2(G128), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT68), .A2(G128), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n240), .B1(new_n244), .B2(new_n191), .ZN(new_n245));
  INV_X1    g059(.A(new_n199), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n205), .B1(new_n246), .B2(KEYINPUT67), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(KEYINPUT67), .B2(new_n246), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(G131), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n211), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n223), .A2(new_n237), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n223), .A2(KEYINPUT30), .A3(new_n250), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n219), .A2(new_n220), .ZN(new_n260));
  INV_X1    g074(.A(new_n197), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n250), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT30), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n236), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n259), .A2(new_n267), .A3(new_n236), .A4(new_n264), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n258), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  INV_X1    g084(.A(new_n257), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n251), .A2(KEYINPUT28), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n223), .A2(new_n273), .A3(new_n237), .A4(new_n250), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n262), .A2(new_n236), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n269), .A2(new_n270), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n268), .ZN(new_n279));
  INV_X1    g093(.A(new_n258), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT71), .B1(new_n281), .B2(KEYINPUT31), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n269), .A2(new_n283), .A3(new_n270), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n278), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n251), .A2(new_n271), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n291), .B1(new_n266), .B2(new_n268), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n237), .B1(new_n223), .B2(new_n250), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n297));
  AOI211_X1 g111(.A(new_n296), .B(new_n297), .C1(new_n272), .C2(new_n274), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n295), .B1(new_n298), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n296), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n275), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT72), .B(new_n300), .C1(new_n302), .C2(new_n297), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n294), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n285), .A2(new_n289), .B1(G472), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n279), .A2(new_n270), .A3(new_n280), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n277), .A2(new_n271), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n283), .B1(new_n269), .B2(new_n270), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n281), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n288), .B1(new_n311), .B2(new_n287), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G217), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(G234), .B2(new_n300), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n317));
  OR2_X1    g131(.A1(KEYINPUT68), .A2(G128), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT68), .A2(G128), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n318), .A2(new_n319), .A3(G119), .A4(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n243), .A2(new_n242), .A3(new_n229), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT73), .B1(new_n238), .B2(G119), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT24), .B(G110), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G110), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT23), .B1(new_n238), .B2(G119), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n238), .A2(G119), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n318), .A2(KEYINPUT23), .A3(G119), .A4(new_n320), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(KEYINPUT74), .A2(G125), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(KEYINPUT74), .A2(G125), .A3(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(KEYINPUT16), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(G125), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n338), .A2(new_n187), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n187), .B1(new_n338), .B2(new_n341), .ZN(new_n343));
  OAI221_X1 g157(.A(new_n327), .B1(new_n328), .B2(new_n333), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n325), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n332), .A3(new_n328), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G140), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n339), .A2(new_n349), .A3(new_n187), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n347), .A2(new_n351), .A3(KEYINPUT75), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT75), .B1(new_n347), .B2(new_n351), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n344), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n355), .B(new_n356), .Z(new_n357));
  AND2_X1   g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(KEYINPUT76), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n344), .B(new_n360), .C1(new_n352), .C2(new_n353), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n357), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n317), .B1(new_n364), .B2(G902), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT25), .B(new_n300), .C1(new_n366), .C2(new_n358), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n316), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n315), .A2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  OR3_X1    g185(.A1(new_n368), .A2(KEYINPUT77), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT77), .B1(new_n368), .B2(new_n371), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n252), .A2(new_n253), .A3(G214), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(G143), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT18), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n377), .B1(new_n378), .B2(new_n203), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n339), .A2(new_n349), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n336), .A2(new_n337), .ZN(new_n381));
  MUX2_X1   g195(.A(new_n380), .B(new_n381), .S(G146), .Z(new_n382));
  XNOR2_X1  g196(.A(new_n376), .B(new_n189), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT18), .A3(G131), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT93), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT93), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(new_n379), .A3(new_n384), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n342), .A2(new_n343), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n383), .A2(KEYINPUT17), .A3(G131), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n377), .B(new_n203), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n390), .B(new_n391), .C1(new_n392), .C2(KEYINPUT17), .ZN(new_n393));
  XNOR2_X1  g207(.A(G113), .B(G122), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT94), .B(G104), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n389), .B2(new_n393), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n300), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G475), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT19), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n380), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(KEYINPUT19), .B2(new_n381), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n343), .B1(new_n404), .B2(new_n187), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n386), .A2(new_n388), .B1(new_n405), .B2(new_n392), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n397), .B1(new_n406), .B2(new_n396), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT20), .ZN(new_n408));
  NOR2_X1   g222(.A1(G475), .A2(G902), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n407), .B2(new_n409), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n401), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G107), .ZN(new_n416));
  INV_X1    g230(.A(G122), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G116), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n416), .B1(new_n418), .B2(KEYINPUT14), .ZN(new_n419));
  XNOR2_X1  g233(.A(G116), .B(G122), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n318), .A2(G143), .A3(new_n320), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n189), .A2(G128), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n204), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n204), .B1(new_n422), .B2(new_n423), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n420), .B(new_n416), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT13), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT95), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n423), .A2(new_n429), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT95), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(new_n189), .A3(KEYINPUT13), .A4(G128), .ZN(new_n433));
  AND4_X1   g247(.A1(new_n430), .A2(new_n422), .A3(new_n431), .A4(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n424), .B(new_n428), .C1(new_n434), .C2(new_n204), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT9), .B(G234), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n436), .A2(new_n314), .A3(G953), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n427), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n427), .B2(new_n435), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n300), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n441), .A2(new_n446), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n415), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G952), .ZN(new_n451));
  AOI211_X1 g265(.A(G953), .B(new_n451), .C1(G234), .C2(G237), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n300), .B(new_n253), .C1(G234), .C2(G237), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n253), .A2(G227), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT78), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G140), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n460), .B(KEYINPUT79), .Z(new_n461));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n462));
  XNOR2_X1  g276(.A(G104), .B(G107), .ZN(new_n463));
  INV_X1    g277(.A(G101), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n416), .A2(G104), .ZN(new_n466));
  INV_X1    g280(.A(G104), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G107), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT82), .A3(G101), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT3), .B1(new_n467), .B2(G107), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT3), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n416), .A3(G104), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n471), .A2(new_n473), .A3(new_n464), .A4(new_n468), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n245), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT83), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n241), .A2(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n240), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT82), .B1(new_n469), .B2(G101), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n462), .B(new_n464), .C1(new_n466), .C2(new_n468), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n195), .A2(new_n239), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n238), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n486), .B2(new_n195), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(KEYINPUT83), .A3(new_n474), .A4(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n477), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n489), .A2(new_n490), .A3(new_n260), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n260), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n220), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n488), .A2(new_n481), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n494), .A2(new_n495), .B1(new_n496), .B2(new_n476), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n492), .B1(new_n497), .B2(KEYINPUT12), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n221), .A2(new_n222), .ZN(new_n499));
  OAI211_X1 g313(.A(KEYINPUT84), .B(new_n490), .C1(new_n499), .C2(new_n489), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n491), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n471), .A2(new_n473), .A3(new_n468), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G101), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT4), .A3(new_n474), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(G101), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n197), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT81), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT81), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n504), .A2(new_n197), .A3(new_n509), .A4(new_n506), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n245), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n465), .A2(new_n470), .A3(new_n474), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT10), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n488), .A2(new_n481), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n511), .B(new_n514), .C1(new_n515), .C2(KEYINPUT10), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n494), .A2(new_n495), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n461), .B1(new_n501), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  INV_X1    g334(.A(new_n460), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n516), .B2(new_n517), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(G469), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G469), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(new_n300), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n491), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n497), .A2(new_n492), .A3(KEYINPUT12), .ZN(new_n530));
  OAI22_X1  g344(.A1(new_n515), .A2(new_n477), .B1(new_n221), .B2(new_n222), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT84), .B1(new_n531), .B2(new_n490), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT85), .ZN(new_n534));
  INV_X1    g348(.A(new_n522), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT85), .B1(new_n501), .B2(new_n522), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n460), .B1(new_n520), .B2(new_n518), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n525), .A3(new_n300), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n528), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G221), .B1(new_n436), .B2(G902), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n233), .A2(new_n234), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT5), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n229), .A3(G116), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT86), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n544), .A2(new_n229), .A3(KEYINPUT86), .A4(G116), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n225), .B1(new_n224), .B2(KEYINPUT5), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n513), .ZN(new_n552));
  XNOR2_X1  g366(.A(G110), .B(G122), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n502), .A2(G101), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n474), .A2(KEYINPUT4), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n236), .B(new_n506), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n236), .A2(new_n506), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n558), .A2(new_n504), .B1(new_n551), .B2(new_n513), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n553), .B(KEYINPUT87), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n557), .B(KEYINPUT6), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n244), .A2(new_n191), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT89), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n348), .A4(new_n485), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n318), .A2(new_n320), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n348), .B(new_n485), .C1(new_n568), .C2(new_n195), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT89), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n348), .B1(new_n194), .B2(new_n196), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G224), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(G953), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n574), .B(new_n567), .C1(new_n570), .C2(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OR3_X1    g392(.A1(new_n559), .A2(KEYINPUT6), .A3(new_n561), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n552), .A2(new_n556), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n560), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n581), .A2(KEYINPUT88), .A3(KEYINPUT6), .A4(new_n557), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n564), .A2(new_n578), .A3(new_n579), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n572), .A2(KEYINPUT7), .A3(new_n575), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n567), .C1(new_n570), .C2(new_n571), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n553), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT5), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n589), .A2(new_n547), .A3(G113), .A4(new_n548), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n228), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n591), .A2(new_n475), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n475), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n584), .A2(new_n586), .A3(new_n577), .A4(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n557), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n583), .B(new_n300), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(G210), .B1(G237), .B2(G902), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n594), .A2(new_n577), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(KEYINPUT91), .A3(new_n584), .A4(new_n586), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n597), .A3(new_n557), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n606), .A2(new_n300), .A3(new_n601), .A4(new_n583), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G214), .B1(G237), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND4_X1   g426(.A1(new_n456), .A2(new_n541), .A3(new_n542), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n313), .A2(new_n375), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  NAND2_X1  g429(.A1(new_n541), .A2(new_n542), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n374), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n285), .A2(new_n286), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n285), .A2(new_n300), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n603), .A2(new_n622), .A3(new_n607), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n600), .A2(KEYINPUT97), .A3(new_n602), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n610), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n439), .A2(KEYINPUT33), .A3(new_n440), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n437), .A2(KEYINPUT99), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n427), .B2(new_n435), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n629), .A2(new_n631), .B1(new_n438), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n629), .B2(new_n631), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n442), .B(new_n628), .C1(new_n634), .C2(KEYINPUT33), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n442), .A2(new_n300), .ZN(new_n636));
  INV_X1    g450(.A(new_n441), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n636), .B1(new_n637), .B2(new_n442), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT100), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n634), .A2(KEYINPUT33), .ZN(new_n641));
  INV_X1    g455(.A(new_n628), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(G478), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n644), .A3(new_n638), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n415), .ZN(new_n647));
  INV_X1    g461(.A(new_n455), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n621), .A2(new_n627), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT101), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NAND3_X1  g467(.A1(new_n407), .A2(new_n412), .A3(new_n409), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n401), .B1(new_n655), .B2(new_n413), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n656), .A2(new_n455), .A3(new_n449), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n603), .A2(new_n607), .A3(new_n622), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n658), .A3(new_n610), .A4(new_n624), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n621), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  INV_X1    g476(.A(new_n542), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n528), .B2(new_n540), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n664), .A2(new_n612), .ZN(new_n665));
  OR3_X1    g479(.A1(new_n362), .A2(KEYINPUT36), .A3(new_n363), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n362), .B1(KEYINPUT36), .B2(new_n363), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n370), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n365), .A2(new_n367), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n668), .B1(new_n669), .B2(new_n315), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n456), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n665), .A2(new_n620), .A3(new_n673), .A4(new_n618), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n304), .A2(G472), .ZN(new_n678));
  INV_X1    g492(.A(new_n289), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n678), .B1(new_n311), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT32), .B1(new_n285), .B2(new_n286), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n623), .A2(new_n670), .A3(new_n625), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT102), .B(G900), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n453), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n452), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n401), .B(new_n687), .C1(new_n655), .C2(new_n413), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n449), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n664), .A2(new_n683), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n677), .B1(new_n682), .B2(new_n690), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n664), .A2(new_n683), .A3(new_n689), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n313), .A2(new_n692), .A3(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  NAND2_X1  g509(.A1(new_n285), .A2(new_n289), .ZN(new_n696));
  INV_X1    g510(.A(new_n251), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n266), .B2(new_n268), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(new_n271), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n301), .A2(new_n251), .A3(new_n271), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT105), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n700), .B(KEYINPUT105), .C1(new_n698), .C2(new_n271), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n300), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n312), .A2(new_n696), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n671), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n608), .B(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n415), .A2(new_n449), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n610), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n687), .B(KEYINPUT39), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n664), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n711), .B1(new_n713), .B2(KEYINPUT40), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n707), .B(new_n714), .C1(KEYINPUT40), .C2(new_n713), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT106), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  NAND4_X1  g531(.A1(new_n640), .A2(new_n414), .A3(new_n645), .A4(new_n687), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT107), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n664), .A3(new_n683), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n682), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n187), .ZN(G48));
  NAND2_X1  g536(.A1(new_n539), .A2(new_n300), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n626), .A2(new_n724), .A3(new_n542), .A4(new_n540), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n649), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n313), .A2(new_n726), .A3(new_n375), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND2_X1  g543(.A1(new_n724), .A2(new_n540), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n730), .A2(new_n659), .A3(new_n663), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n313), .A2(new_n375), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NOR2_X1   g547(.A1(new_n725), .A2(new_n672), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n313), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  INV_X1    g550(.A(new_n710), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n725), .A2(new_n455), .A3(new_n737), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n269), .A2(new_n270), .B1(new_n271), .B2(new_n302), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n281), .A2(KEYINPUT31), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n287), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n619), .B2(G472), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n368), .A2(new_n371), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT108), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(G472), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n285), .B2(new_n300), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  INV_X1    g561(.A(new_n743), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n741), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n738), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  INV_X1    g565(.A(new_n725), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n742), .A2(new_n671), .A3(new_n752), .A4(new_n719), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  NOR2_X1   g568(.A1(new_n608), .A2(new_n611), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT109), .B1(new_n616), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n664), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n719), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n313), .A2(new_n743), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT42), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n719), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(KEYINPUT42), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n374), .B1(new_n305), .B2(new_n312), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n757), .A4(new_n759), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n203), .ZN(G33));
  XOR2_X1   g582(.A(new_n689), .B(KEYINPUT110), .Z(new_n769));
  NAND4_X1  g583(.A1(new_n765), .A2(new_n757), .A3(new_n759), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  NAND2_X1  g585(.A1(new_n620), .A2(new_n618), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n415), .A2(new_n640), .A3(new_n645), .ZN(new_n773));
  NAND2_X1  g587(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n772), .A2(new_n671), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n756), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n772), .A2(KEYINPUT44), .A3(new_n671), .A4(new_n777), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(KEYINPUT112), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n519), .B2(new_n523), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n525), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n519), .A2(KEYINPUT45), .A3(new_n523), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT46), .B1(new_n786), .B2(new_n527), .ZN(new_n787));
  INV_X1    g601(.A(new_n540), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n527), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n663), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n712), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT112), .B1(new_n780), .B2(new_n781), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n198), .ZN(G39));
  NAND4_X1  g610(.A1(new_n682), .A2(new_n374), .A3(new_n719), .A4(new_n755), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n791), .A2(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n791), .A2(KEYINPUT47), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n335), .ZN(G42));
  OR4_X1    g615(.A1(new_n748), .A2(new_n773), .A3(new_n663), .A4(new_n611), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n709), .B(new_n802), .C1(KEYINPUT49), .C2(new_n730), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n803), .B(new_n706), .C1(KEYINPUT49), .C2(new_n730), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n646), .A2(new_n414), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n648), .A2(new_n612), .A3(new_n450), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n617), .A2(new_n620), .A3(new_n806), .A4(new_n618), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n727), .A2(new_n732), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n614), .A2(new_n674), .A3(new_n735), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n750), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n746), .A2(new_n670), .A3(new_n741), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n719), .A3(new_n757), .A4(new_n759), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n670), .A2(new_n447), .A3(new_n448), .A4(new_n688), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n313), .A2(new_n664), .A3(new_n755), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n770), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n810), .A2(new_n767), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n682), .A2(new_n720), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n313), .A2(new_n692), .A3(KEYINPUT103), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT103), .B1(new_n313), .B2(new_n692), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n687), .B(KEYINPUT113), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n664), .A2(new_n626), .A3(new_n710), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n705), .A2(new_n823), .A3(new_n670), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n753), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n817), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n721), .B1(new_n691), .B2(new_n693), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n824), .A2(new_n753), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(KEYINPUT52), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n808), .A2(new_n809), .A3(new_n750), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n767), .A2(new_n815), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n821), .A2(new_n817), .A3(new_n825), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n826), .B1(new_n835), .B2(KEYINPUT114), .ZN(new_n836));
  AOI211_X1 g650(.A(KEYINPUT114), .B(KEYINPUT52), .C1(new_n827), .C2(new_n828), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n834), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n831), .B1(new_n839), .B2(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT54), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT52), .B1(new_n827), .B2(new_n828), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n843), .B1(new_n844), .B2(new_n829), .ZN(new_n845));
  OAI211_X1 g659(.A(KEYINPUT53), .B(new_n816), .C1(new_n845), .C2(new_n837), .ZN(new_n846));
  AOI211_X1 g660(.A(KEYINPUT115), .B(KEYINPUT53), .C1(new_n816), .C2(new_n830), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n832), .B(new_n833), .C1(new_n835), .C2(new_n843), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n842), .B(new_n846), .C1(new_n847), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n798), .B(new_n799), .C1(new_n542), .C2(new_n730), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n777), .A2(new_n452), .ZN(new_n855));
  INV_X1    g669(.A(new_n744), .ZN(new_n856));
  INV_X1    g670(.A(new_n749), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n755), .A3(new_n858), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n730), .A2(new_n686), .A3(new_n756), .A4(new_n663), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n706), .A2(new_n375), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n415), .A3(new_n646), .ZN(new_n862));
  INV_X1    g676(.A(new_n811), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n777), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n730), .A2(new_n663), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n709), .A2(new_n610), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(KEYINPUT50), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n858), .A2(new_n866), .A3(new_n868), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT50), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n865), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n874));
  OAI211_X1 g688(.A(KEYINPUT51), .B(new_n859), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n874), .B2(new_n873), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n861), .A2(new_n647), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(G952), .A3(new_n253), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n864), .A2(new_n761), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT48), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n878), .B(new_n880), .C1(new_n626), .C2(new_n867), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n873), .A2(new_n859), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n853), .A2(new_n876), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(G952), .A2(G953), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT118), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n804), .B1(new_n885), .B2(new_n887), .ZN(G75));
  NAND2_X1  g702(.A1(new_n451), .A2(G953), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT119), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n846), .B1(new_n847), .B2(new_n851), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(G902), .ZN(new_n893));
  INV_X1    g707(.A(G210), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n564), .A2(new_n579), .A3(new_n582), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(new_n578), .Z(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n890), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n895), .B2(new_n898), .ZN(G51));
  INV_X1    g714(.A(new_n890), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n852), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n892), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n526), .B(KEYINPUT57), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n539), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n893), .A2(new_n786), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND4_X1  g724(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n911));
  INV_X1    g725(.A(new_n407), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n911), .A2(KEYINPUT121), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT121), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n901), .B1(new_n911), .B2(new_n912), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G60));
  NAND2_X1  g730(.A1(new_n641), .A2(new_n642), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n636), .B(KEYINPUT59), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n917), .A2(new_n904), .A3(new_n905), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n841), .B2(new_n852), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n890), .B1(new_n921), .B2(new_n917), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n922), .ZN(G63));
  XNOR2_X1  g737(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n314), .A2(new_n300), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n892), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n364), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n666), .A2(new_n667), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n892), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n890), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G66));
  OAI21_X1  g748(.A(G953), .B1(new_n454), .B2(new_n573), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n832), .B2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n896), .B1(G898), .B2(new_n253), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G69));
  AOI21_X1  g752(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n259), .A2(new_n264), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n404), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n694), .A2(new_n818), .A3(new_n753), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT124), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n761), .A2(new_n627), .A3(new_n737), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n792), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n800), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n793), .B2(new_n794), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n762), .A2(new_n766), .A3(new_n770), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT125), .Z(new_n952));
  AOI21_X1  g766(.A(G953), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n253), .A2(G900), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n942), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n949), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n956), .A2(new_n944), .A3(new_n952), .A4(new_n946), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n253), .ZN(new_n958));
  INV_X1    g772(.A(new_n954), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n958), .A2(KEYINPUT126), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n941), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n941), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n944), .A2(new_n716), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n944), .A2(new_n965), .A3(new_n716), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n805), .A2(new_n755), .A3(new_n450), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n713), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n765), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n964), .A2(new_n966), .A3(new_n969), .A4(new_n956), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n962), .B1(new_n970), .B2(new_n253), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n939), .B1(new_n961), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT126), .B1(new_n958), .B2(new_n959), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n942), .B(new_n954), .C1(new_n957), .C2(new_n253), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n962), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n939), .ZN(new_n976));
  INV_X1    g790(.A(new_n971), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n972), .A2(new_n978), .ZN(G72));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n970), .B2(new_n810), .ZN(new_n982));
  INV_X1    g796(.A(new_n699), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n981), .B1(new_n957), .B2(new_n810), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n292), .ZN(new_n986));
  INV_X1    g800(.A(new_n292), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n699), .A2(new_n987), .A3(new_n981), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n901), .B1(new_n840), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n984), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n984), .A2(new_n989), .A3(new_n992), .A4(new_n986), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(G57));
endmodule


