

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781;

  NOR2_X1 U374 ( .A1(n418), .A2(n417), .ZN(n416) );
  NOR2_X1 U375 ( .A1(n694), .A2(n695), .ZN(n699) );
  XNOR2_X1 U376 ( .A(n528), .B(n474), .ZN(n766) );
  XNOR2_X1 U377 ( .A(n611), .B(n580), .ZN(n711) );
  XNOR2_X1 U378 ( .A(n634), .B(n482), .ZN(n637) );
  NAND2_X1 U379 ( .A1(n450), .A2(n448), .ZN(n769) );
  NAND2_X1 U380 ( .A1(n637), .A2(n642), .ZN(n644) );
  INV_X1 U381 ( .A(n638), .ZN(n694) );
  XNOR2_X2 U382 ( .A(n451), .B(KEYINPUT108), .ZN(n714) );
  NOR2_X1 U383 ( .A1(n700), .A2(n636), .ZN(n675) );
  NAND2_X1 U384 ( .A1(n700), .A2(n699), .ZN(n650) );
  NAND2_X1 U385 ( .A1(n426), .A2(n777), .ZN(n655) );
  NAND2_X1 U386 ( .A1(n391), .A2(n387), .ZN(n647) );
  XOR2_X1 U387 ( .A(G146), .B(G125), .Z(n527) );
  XNOR2_X1 U388 ( .A(KEYINPUT97), .B(n649), .ZN(n672) );
  AND2_X1 U389 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U390 ( .A1(n651), .A2(n633), .ZN(n634) );
  NAND2_X1 U391 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U392 ( .A1(n488), .A2(n486), .ZN(n709) );
  NOR2_X1 U393 ( .A1(n443), .A2(n368), .ZN(n587) );
  XNOR2_X1 U394 ( .A(n739), .B(n738), .ZN(n741) );
  OR2_X1 U395 ( .A1(n639), .A2(n638), .ZN(n494) );
  XNOR2_X1 U396 ( .A(n564), .B(n563), .ZN(n638) );
  XNOR2_X1 U397 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U398 ( .A(n360), .B(n446), .ZN(n746) );
  XNOR2_X1 U399 ( .A(n520), .B(n457), .ZN(n743) );
  INV_X1 U400 ( .A(n754), .ZN(n479) );
  XNOR2_X1 U401 ( .A(n538), .B(n766), .ZN(n446) );
  XNOR2_X1 U402 ( .A(n768), .B(G146), .ZN(n520) );
  XNOR2_X1 U403 ( .A(n544), .B(n543), .ZN(n556) );
  XNOR2_X1 U404 ( .A(n548), .B(n483), .ZN(n768) );
  NAND2_X1 U405 ( .A1(n507), .A2(n506), .ZN(n547) );
  BUF_X1 U406 ( .A(n542), .Z(n497) );
  XNOR2_X1 U407 ( .A(n498), .B(n484), .ZN(n483) );
  XNOR2_X1 U408 ( .A(n485), .B(G137), .ZN(n484) );
  XNOR2_X1 U409 ( .A(n514), .B(G134), .ZN(n548) );
  XNOR2_X1 U410 ( .A(n496), .B(KEYINPUT64), .ZN(n542) );
  INV_X1 U411 ( .A(G953), .ZN(n496) );
  XNOR2_X1 U412 ( .A(G143), .B(G128), .ZN(n514) );
  XNOR2_X1 U413 ( .A(n640), .B(KEYINPUT32), .ZN(n353) );
  NAND2_X1 U414 ( .A1(n428), .A2(n427), .ZN(n356) );
  NAND2_X1 U415 ( .A1(n354), .A2(n355), .ZN(n357) );
  NAND2_X1 U416 ( .A1(n356), .A2(n357), .ZN(n760) );
  INV_X1 U417 ( .A(n428), .ZN(n354) );
  INV_X1 U418 ( .A(n427), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n640), .B(KEYINPUT32), .ZN(n779) );
  XNOR2_X2 U420 ( .A(G101), .B(G113), .ZN(n429) );
  XNOR2_X2 U421 ( .A(n453), .B(G119), .ZN(n430) );
  INV_X2 U422 ( .A(KEYINPUT3), .ZN(n453) );
  NAND2_X1 U423 ( .A1(n416), .A2(n413), .ZN(n412) );
  XNOR2_X2 U424 ( .A(n630), .B(n629), .ZN(n651) );
  XNOR2_X2 U425 ( .A(n430), .B(n429), .ZN(n447) );
  NAND2_X1 U426 ( .A1(n421), .A2(n375), .ZN(n419) );
  NAND2_X1 U427 ( .A1(n406), .A2(n405), .ZN(n404) );
  OR2_X1 U428 ( .A1(n585), .A2(KEYINPUT107), .ZN(n468) );
  AND2_X1 U429 ( .A1(n490), .A2(n489), .ZN(n488) );
  NAND2_X1 U430 ( .A1(n487), .A2(n358), .ZN(n486) );
  NAND2_X1 U431 ( .A1(n642), .A2(n371), .ZN(n489) );
  XNOR2_X1 U432 ( .A(n571), .B(KEYINPUT21), .ZN(n695) );
  INV_X1 U433 ( .A(KEYINPUT10), .ZN(n474) );
  INV_X1 U434 ( .A(KEYINPUT77), .ZN(n432) );
  NAND2_X1 U435 ( .A1(n400), .A2(n399), .ZN(n398) );
  XNOR2_X1 U436 ( .A(n473), .B(n590), .ZN(n621) );
  NAND2_X1 U437 ( .A1(n655), .A2(n374), .ZN(n415) );
  AND2_X1 U438 ( .A1(n695), .A2(n471), .ZN(n466) );
  NOR2_X1 U439 ( .A1(n411), .A2(n408), .ZN(n407) );
  XNOR2_X1 U440 ( .A(n404), .B(n593), .ZN(n403) );
  OR2_X1 U441 ( .A1(n599), .A2(n617), .ZN(n411) );
  XOR2_X1 U442 ( .A(G122), .B(G104), .Z(n529) );
  XNOR2_X1 U443 ( .A(n522), .B(n460), .ZN(n459) );
  INV_X1 U444 ( .A(G101), .ZN(n460) );
  XOR2_X1 U445 ( .A(G107), .B(G104), .Z(n522) );
  XOR2_X1 U446 ( .A(G140), .B(G110), .Z(n523) );
  INV_X1 U447 ( .A(n555), .ZN(n390) );
  INV_X1 U448 ( .A(G902), .ZN(n389) );
  NAND2_X1 U449 ( .A1(n555), .A2(G902), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n561), .B(n444), .ZN(n570) );
  XNOR2_X1 U451 ( .A(KEYINPUT20), .B(KEYINPUT94), .ZN(n444) );
  XNOR2_X1 U452 ( .A(n647), .B(n370), .ZN(n642) );
  INV_X1 U453 ( .A(n401), .ZN(n397) );
  NAND2_X1 U454 ( .A1(n641), .A2(n384), .ZN(n382) );
  NAND2_X1 U455 ( .A1(n709), .A2(n384), .ZN(n383) );
  NAND2_X1 U456 ( .A1(n380), .A2(n379), .ZN(n378) );
  NOR2_X1 U457 ( .A1(n641), .A2(n384), .ZN(n379) );
  AND2_X1 U458 ( .A1(n589), .A2(n362), .ZN(n609) );
  INV_X1 U459 ( .A(n647), .ZN(n698) );
  NOR2_X1 U460 ( .A1(n743), .A2(G902), .ZN(n526) );
  XNOR2_X1 U461 ( .A(n475), .B(n766), .ZN(n753) );
  INV_X1 U462 ( .A(KEYINPUT123), .ZN(n463) );
  NOR2_X1 U463 ( .A1(n497), .A2(G952), .ZN(n754) );
  NAND2_X1 U464 ( .A1(n731), .A2(n369), .ZN(n456) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n408) );
  INV_X1 U466 ( .A(KEYINPUT85), .ZN(n409) );
  INV_X1 U467 ( .A(KEYINPUT4), .ZN(n485) );
  OR2_X1 U468 ( .A1(G237), .A2(G902), .ZN(n574) );
  XNOR2_X1 U469 ( .A(n547), .B(KEYINPUT16), .ZN(n431) );
  XNOR2_X1 U470 ( .A(G902), .B(KEYINPUT15), .ZN(n658) );
  XOR2_X1 U471 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n512) );
  XNOR2_X1 U472 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n509) );
  NAND2_X1 U473 ( .A1(G234), .A2(G237), .ZN(n565) );
  INV_X1 U474 ( .A(KEYINPUT34), .ZN(n384) );
  NAND2_X1 U475 ( .A1(n469), .A2(n468), .ZN(n443) );
  NOR2_X1 U476 ( .A1(n449), .A2(n778), .ZN(n448) );
  INV_X1 U477 ( .A(n693), .ZN(n449) );
  XNOR2_X1 U478 ( .A(n529), .B(n508), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n447), .B(n431), .ZN(n428) );
  XOR2_X1 U480 ( .A(G110), .B(KEYINPUT74), .Z(n508) );
  XOR2_X1 U481 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n559) );
  XNOR2_X1 U482 ( .A(KEYINPUT98), .B(KEYINPUT12), .ZN(n531) );
  XOR2_X1 U483 ( .A(G131), .B(KEYINPUT100), .Z(n537) );
  XNOR2_X1 U484 ( .A(G113), .B(G143), .ZN(n530) );
  XNOR2_X1 U485 ( .A(n521), .B(n458), .ZN(n457) );
  XNOR2_X1 U486 ( .A(n459), .B(n523), .ZN(n458) );
  NAND2_X1 U487 ( .A1(n367), .A2(n398), .ZN(n733) );
  INV_X1 U488 ( .A(KEYINPUT105), .ZN(n436) );
  BUF_X1 U489 ( .A(n594), .Z(n611) );
  XNOR2_X1 U490 ( .A(KEYINPUT22), .B(KEYINPUT73), .ZN(n482) );
  OR2_X1 U491 ( .A1(n554), .A2(n388), .ZN(n387) );
  NAND2_X1 U492 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U493 ( .A(n562), .B(KEYINPUT25), .ZN(n563) );
  NOR2_X1 U494 ( .A1(n753), .A2(G902), .ZN(n564) );
  XNOR2_X1 U495 ( .A(n554), .B(KEYINPUT62), .ZN(n662) );
  AND2_X1 U496 ( .A1(n398), .A2(n394), .ZN(n584) );
  AND2_X1 U497 ( .A1(n396), .A2(n395), .ZN(n394) );
  NOR2_X1 U498 ( .A1(n600), .A2(n397), .ZN(n396) );
  XNOR2_X1 U499 ( .A(n592), .B(n591), .ZN(n780) );
  INV_X1 U500 ( .A(KEYINPUT35), .ZN(n492) );
  NAND2_X1 U501 ( .A1(n381), .A2(n378), .ZN(n386) );
  XNOR2_X1 U502 ( .A(n464), .B(n462), .ZN(n461) );
  XNOR2_X1 U503 ( .A(n753), .B(n463), .ZN(n462) );
  XNOR2_X1 U504 ( .A(n750), .B(n433), .ZN(n752) );
  XNOR2_X1 U505 ( .A(n751), .B(KEYINPUT122), .ZN(n433) );
  AND2_X1 U506 ( .A1(n454), .A2(n622), .ZN(n735) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n454) );
  INV_X1 U508 ( .A(KEYINPUT120), .ZN(n455) );
  NOR2_X1 U509 ( .A1(n642), .A2(n371), .ZN(n358) );
  OR2_X1 U510 ( .A1(n734), .A2(n733), .ZN(n359) );
  XOR2_X1 U511 ( .A(n534), .B(n533), .Z(n360) );
  XOR2_X1 U512 ( .A(n500), .B(n499), .Z(n361) );
  XOR2_X1 U513 ( .A(KEYINPUT30), .B(n588), .Z(n362) );
  OR2_X1 U514 ( .A1(n695), .A2(n471), .ZN(n363) );
  OR2_X1 U515 ( .A1(n715), .A2(n653), .ZN(n364) );
  AND2_X1 U516 ( .A1(n699), .A2(n585), .ZN(n365) );
  AND2_X1 U517 ( .A1(n491), .A2(n666), .ZN(n366) );
  AND2_X1 U518 ( .A1(n395), .A2(n401), .ZN(n367) );
  NAND2_X1 U519 ( .A1(n467), .A2(n465), .ZN(n368) );
  AND2_X1 U520 ( .A1(n732), .A2(n359), .ZN(n369) );
  XOR2_X1 U521 ( .A(KEYINPUT6), .B(KEYINPUT103), .Z(n370) );
  XOR2_X1 U522 ( .A(KEYINPUT104), .B(KEYINPUT33), .Z(n371) );
  XOR2_X1 U523 ( .A(KEYINPUT45), .B(KEYINPUT66), .Z(n372) );
  XOR2_X1 U524 ( .A(n743), .B(n744), .Z(n373) );
  AND2_X1 U525 ( .A1(n423), .A2(n654), .ZN(n374) );
  AND2_X1 U526 ( .A1(KEYINPUT44), .A2(n654), .ZN(n375) );
  AND2_X1 U527 ( .A1(KEYINPUT44), .A2(n423), .ZN(n376) );
  INV_X1 U528 ( .A(KEYINPUT2), .ZN(n438) );
  OR2_X1 U529 ( .A1(n658), .A2(n438), .ZN(n377) );
  INV_X1 U530 ( .A(n709), .ZN(n380) );
  XNOR2_X2 U531 ( .A(n385), .B(n492), .ZN(n777) );
  NAND2_X1 U532 ( .A1(n386), .A2(n643), .ZN(n385) );
  AND2_X1 U533 ( .A1(n393), .A2(n392), .ZN(n391) );
  NAND2_X1 U534 ( .A1(n554), .A2(n555), .ZN(n393) );
  NAND2_X1 U535 ( .A1(n714), .A2(n402), .ZN(n395) );
  NOR2_X1 U536 ( .A1(n713), .A2(n402), .ZN(n399) );
  INV_X1 U537 ( .A(n714), .ZN(n400) );
  NAND2_X1 U538 ( .A1(n713), .A2(n402), .ZN(n401) );
  INV_X1 U539 ( .A(KEYINPUT41), .ZN(n402) );
  NAND2_X1 U540 ( .A1(n407), .A2(n403), .ZN(n472) );
  INV_X1 U541 ( .A(n780), .ZN(n405) );
  INV_X1 U542 ( .A(n781), .ZN(n406) );
  NAND2_X1 U543 ( .A1(n616), .A2(n615), .ZN(n410) );
  XNOR2_X2 U544 ( .A(n412), .B(n372), .ZN(n726) );
  NAND2_X1 U545 ( .A1(n415), .A2(n414), .ZN(n413) );
  NAND2_X1 U546 ( .A1(n442), .A2(KEYINPUT44), .ZN(n414) );
  NAND2_X1 U547 ( .A1(n364), .A2(n419), .ZN(n417) );
  NAND2_X1 U548 ( .A1(n366), .A2(n420), .ZN(n418) );
  NAND2_X1 U549 ( .A1(n422), .A2(n376), .ZN(n420) );
  INV_X1 U550 ( .A(n777), .ZN(n421) );
  INV_X1 U551 ( .A(n656), .ZN(n422) );
  INV_X1 U552 ( .A(KEYINPUT67), .ZN(n423) );
  NAND2_X1 U553 ( .A1(n439), .A2(n377), .ZN(n441) );
  AND2_X1 U554 ( .A1(n441), .A2(n730), .ZN(n424) );
  AND2_X2 U555 ( .A1(n441), .A2(n730), .ZN(n452) );
  XNOR2_X1 U556 ( .A(n520), .B(n503), .ZN(n554) );
  XNOR2_X1 U557 ( .A(n472), .B(n620), .ZN(n450) );
  NAND2_X1 U558 ( .A1(n495), .A2(n659), .ZN(n660) );
  XNOR2_X1 U559 ( .A(n477), .B(n476), .ZN(n475) );
  INV_X1 U560 ( .A(n641), .ZN(n425) );
  NOR2_X1 U561 ( .A1(n779), .A2(n675), .ZN(n426) );
  XNOR2_X2 U562 ( .A(n660), .B(n432), .ZN(n730) );
  XNOR2_X1 U563 ( .A(n740), .B(n741), .ZN(n742) );
  XNOR2_X1 U564 ( .A(n661), .B(n662), .ZN(n663) );
  NAND2_X1 U565 ( .A1(n452), .A2(G475), .ZN(n748) );
  XNOR2_X1 U566 ( .A(n434), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U567 ( .A1(n749), .A2(n754), .ZN(n434) );
  NOR2_X2 U568 ( .A1(n726), .A2(n658), .ZN(n657) );
  INV_X1 U569 ( .A(n769), .ZN(n659) );
  NAND2_X1 U570 ( .A1(n435), .A2(n683), .ZN(n595) );
  XNOR2_X1 U571 ( .A(n573), .B(n436), .ZN(n435) );
  NAND2_X1 U572 ( .A1(n647), .A2(n710), .ZN(n588) );
  XNOR2_X1 U573 ( .A(n437), .B(n665), .ZN(G57) );
  NOR2_X2 U574 ( .A1(n663), .A2(n754), .ZN(n437) );
  XNOR2_X1 U575 ( .A(n657), .B(KEYINPUT88), .ZN(n440) );
  NOR2_X1 U576 ( .A1(n726), .A2(n438), .ZN(n495) );
  NAND2_X1 U577 ( .A1(n440), .A2(n659), .ZN(n439) );
  NAND2_X1 U578 ( .A1(n426), .A2(KEYINPUT67), .ZN(n442) );
  NOR2_X1 U579 ( .A1(n466), .A2(n586), .ZN(n465) );
  NAND2_X1 U580 ( .A1(n452), .A2(G210), .ZN(n740) );
  NOR2_X2 U581 ( .A1(n644), .A2(n494), .ZN(n640) );
  XNOR2_X1 U582 ( .A(n445), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U583 ( .A1(n742), .A2(n754), .ZN(n445) );
  AND2_X1 U584 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U585 ( .A(n447), .B(n361), .ZN(n502) );
  NAND2_X1 U586 ( .A1(n711), .A2(n710), .ZN(n451) );
  NAND2_X1 U587 ( .A1(n452), .A2(G472), .ZN(n661) );
  NAND2_X1 U588 ( .A1(n424), .A2(G478), .ZN(n750) );
  NAND2_X1 U589 ( .A1(n424), .A2(G469), .ZN(n481) );
  NAND2_X1 U590 ( .A1(n424), .A2(G217), .ZN(n464) );
  NOR2_X1 U591 ( .A1(n461), .A2(n754), .ZN(G66) );
  XNOR2_X2 U592 ( .A(n602), .B(n601), .ZN(n628) );
  NAND2_X2 U593 ( .A1(n594), .A2(n710), .ZN(n602) );
  XNOR2_X2 U594 ( .A(n519), .B(n518), .ZN(n594) );
  NAND2_X1 U595 ( .A1(n694), .A2(n471), .ZN(n467) );
  NAND2_X1 U596 ( .A1(n585), .A2(n470), .ZN(n469) );
  NOR2_X1 U597 ( .A1(n694), .A2(n363), .ZN(n470) );
  INV_X1 U598 ( .A(KEYINPUT107), .ZN(n471) );
  NAND2_X1 U599 ( .A1(n621), .A2(n683), .ZN(n592) );
  NAND2_X1 U600 ( .A1(n609), .A2(n711), .ZN(n473) );
  XNOR2_X1 U601 ( .A(n560), .B(n559), .ZN(n476) );
  NAND2_X1 U602 ( .A1(n556), .A2(G221), .ZN(n477) );
  XNOR2_X1 U603 ( .A(n478), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U604 ( .A1(n480), .A2(n479), .ZN(n478) );
  XNOR2_X1 U605 ( .A(n481), .B(n373), .ZN(n480) );
  NAND2_X1 U606 ( .A1(n650), .A2(n371), .ZN(n490) );
  INV_X1 U607 ( .A(n650), .ZN(n487) );
  NAND2_X1 U608 ( .A1(n777), .A2(KEYINPUT93), .ZN(n491) );
  BUF_X1 U609 ( .A(n709), .Z(n734) );
  AND2_X1 U610 ( .A1(n727), .A2(n438), .ZN(n493) );
  INV_X1 U611 ( .A(KEYINPUT93), .ZN(n654) );
  INV_X1 U612 ( .A(n695), .ZN(n631) );
  INV_X1 U613 ( .A(KEYINPUT89), .ZN(n618) );
  INV_X1 U614 ( .A(n723), .ZN(n626) );
  XNOR2_X1 U615 ( .A(n619), .B(n618), .ZN(n620) );
  AND2_X1 U616 ( .A1(n626), .A2(n625), .ZN(n627) );
  INV_X1 U617 ( .A(KEYINPUT0), .ZN(n629) );
  XNOR2_X1 U618 ( .A(n524), .B(G469), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U620 ( .A(n664), .B(KEYINPUT110), .ZN(n665) );
  XNOR2_X1 U621 ( .A(G131), .B(KEYINPUT69), .ZN(n498) );
  XOR2_X1 U622 ( .A(KEYINPUT95), .B(KEYINPUT76), .Z(n500) );
  XNOR2_X1 U623 ( .A(G116), .B(KEYINPUT5), .ZN(n499) );
  INV_X1 U624 ( .A(G953), .ZN(n622) );
  NOR2_X1 U625 ( .A1(G953), .A2(G237), .ZN(n535) );
  NAND2_X1 U626 ( .A1(n535), .A2(G210), .ZN(n501) );
  XNOR2_X1 U627 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U628 ( .A(G107), .ZN(n504) );
  NAND2_X1 U629 ( .A1(G116), .A2(n504), .ZN(n507) );
  INV_X1 U630 ( .A(G116), .ZN(n505) );
  NAND2_X1 U631 ( .A1(n505), .A2(G107), .ZN(n506) );
  XNOR2_X1 U632 ( .A(n509), .B(n527), .ZN(n510) );
  XNOR2_X1 U633 ( .A(n760), .B(n510), .ZN(n517) );
  NAND2_X1 U634 ( .A1(G224), .A2(n542), .ZN(n511) );
  XNOR2_X1 U635 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U636 ( .A(KEYINPUT17), .B(n513), .ZN(n515) );
  XNOR2_X1 U637 ( .A(n514), .B(n515), .ZN(n516) );
  XNOR2_X1 U638 ( .A(n517), .B(n516), .ZN(n736) );
  NAND2_X1 U639 ( .A1(n736), .A2(n658), .ZN(n519) );
  AND2_X1 U640 ( .A1(G210), .A2(n574), .ZN(n518) );
  NAND2_X1 U641 ( .A1(G227), .A2(n497), .ZN(n521) );
  XNOR2_X1 U642 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n524) );
  XNOR2_X2 U643 ( .A(n526), .B(n525), .ZN(n585) );
  XNOR2_X2 U644 ( .A(n585), .B(KEYINPUT1), .ZN(n700) );
  XNOR2_X1 U645 ( .A(n527), .B(G140), .ZN(n528) );
  XNOR2_X1 U646 ( .A(n530), .B(n529), .ZN(n534) );
  XOR2_X1 U647 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n532) );
  XNOR2_X1 U648 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U649 ( .A1(G214), .A2(n535), .ZN(n536) );
  XNOR2_X1 U650 ( .A(n537), .B(n536), .ZN(n538) );
  NOR2_X1 U651 ( .A1(G902), .A2(n746), .ZN(n540) );
  XNOR2_X1 U652 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n539) );
  XNOR2_X1 U653 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U654 ( .A(G475), .B(n541), .ZN(n608) );
  INV_X1 U655 ( .A(n608), .ZN(n605) );
  XOR2_X1 U656 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n546) );
  XOR2_X1 U657 ( .A(KEYINPUT86), .B(KEYINPUT8), .Z(n544) );
  NAND2_X1 U658 ( .A1(G234), .A2(n542), .ZN(n543) );
  NAND2_X1 U659 ( .A1(G217), .A2(n556), .ZN(n545) );
  XNOR2_X1 U660 ( .A(n546), .B(n545), .ZN(n552) );
  XOR2_X1 U661 ( .A(KEYINPUT7), .B(n547), .Z(n550) );
  XNOR2_X1 U662 ( .A(n548), .B(G122), .ZN(n549) );
  XNOR2_X1 U663 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U664 ( .A(n552), .B(n551), .Z(n751) );
  NOR2_X1 U665 ( .A1(n751), .A2(G902), .ZN(n553) );
  XNOR2_X1 U666 ( .A(n553), .B(G478), .ZN(n607) );
  AND2_X1 U667 ( .A1(n605), .A2(n607), .ZN(n683) );
  XNOR2_X1 U668 ( .A(G472), .B(KEYINPUT96), .ZN(n555) );
  XOR2_X1 U669 ( .A(G110), .B(G137), .Z(n558) );
  XNOR2_X1 U670 ( .A(G119), .B(G128), .ZN(n557) );
  XNOR2_X1 U671 ( .A(n558), .B(n557), .ZN(n560) );
  NAND2_X1 U672 ( .A1(n658), .A2(G234), .ZN(n561) );
  NAND2_X1 U673 ( .A1(G217), .A2(n570), .ZN(n562) );
  XOR2_X1 U674 ( .A(n565), .B(KEYINPUT14), .Z(n723) );
  NOR2_X1 U675 ( .A1(n497), .A2(G900), .ZN(n566) );
  NAND2_X1 U676 ( .A1(G902), .A2(n566), .ZN(n567) );
  NAND2_X1 U677 ( .A1(G952), .A2(n622), .ZN(n623) );
  NAND2_X1 U678 ( .A1(n567), .A2(n623), .ZN(n568) );
  NAND2_X1 U679 ( .A1(n626), .A2(n568), .ZN(n569) );
  XNOR2_X1 U680 ( .A(KEYINPUT82), .B(n569), .ZN(n586) );
  NAND2_X1 U681 ( .A1(n570), .A2(G221), .ZN(n571) );
  NOR2_X1 U682 ( .A1(n586), .A2(n695), .ZN(n572) );
  NAND2_X1 U683 ( .A1(n694), .A2(n572), .ZN(n581) );
  NOR2_X1 U684 ( .A1(n642), .A2(n581), .ZN(n573) );
  INV_X1 U685 ( .A(n595), .ZN(n575) );
  NAND2_X1 U686 ( .A1(G214), .A2(n574), .ZN(n710) );
  NAND2_X1 U687 ( .A1(n575), .A2(n710), .ZN(n576) );
  NOR2_X1 U688 ( .A1(n700), .A2(n576), .ZN(n577) );
  XNOR2_X1 U689 ( .A(n577), .B(KEYINPUT43), .ZN(n578) );
  NOR2_X1 U690 ( .A1(n611), .A2(n578), .ZN(n579) );
  XNOR2_X1 U691 ( .A(KEYINPUT106), .B(n579), .ZN(n778) );
  XNOR2_X1 U692 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n580) );
  NAND2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n713) );
  NOR2_X1 U694 ( .A1(n698), .A2(n581), .ZN(n582) );
  XNOR2_X1 U695 ( .A(n582), .B(KEYINPUT28), .ZN(n583) );
  NAND2_X1 U696 ( .A1(n583), .A2(n585), .ZN(n600) );
  XNOR2_X1 U697 ( .A(n584), .B(KEYINPUT42), .ZN(n781) );
  XNOR2_X1 U698 ( .A(n587), .B(KEYINPUT78), .ZN(n589) );
  XOR2_X1 U699 ( .A(KEYINPUT91), .B(KEYINPUT39), .Z(n590) );
  INV_X1 U700 ( .A(KEYINPUT40), .ZN(n591) );
  XNOR2_X1 U701 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n593) );
  NOR2_X1 U702 ( .A1(n595), .A2(n602), .ZN(n597) );
  XNOR2_X1 U703 ( .A(KEYINPUT109), .B(KEYINPUT36), .ZN(n596) );
  XNOR2_X1 U704 ( .A(n597), .B(n596), .ZN(n598) );
  INV_X1 U705 ( .A(n700), .ZN(n639) );
  NOR2_X1 U706 ( .A1(n598), .A2(n639), .ZN(n690) );
  XNOR2_X1 U707 ( .A(n690), .B(KEYINPUT90), .ZN(n599) );
  INV_X1 U708 ( .A(n600), .ZN(n603) );
  XNOR2_X1 U709 ( .A(KEYINPUT19), .B(KEYINPUT68), .ZN(n601) );
  NAND2_X1 U710 ( .A1(n603), .A2(n628), .ZN(n604) );
  XOR2_X1 U711 ( .A(n604), .B(KEYINPUT81), .Z(n614) );
  INV_X1 U712 ( .A(n614), .ZN(n681) );
  NOR2_X1 U713 ( .A1(n605), .A2(n607), .ZN(n686) );
  NOR2_X1 U714 ( .A1(n683), .A2(n686), .ZN(n715) );
  NOR2_X1 U715 ( .A1(KEYINPUT47), .A2(n715), .ZN(n606) );
  AND2_X1 U716 ( .A1(n681), .A2(n606), .ZN(n617) );
  NAND2_X1 U717 ( .A1(KEYINPUT47), .A2(n715), .ZN(n612) );
  NOR2_X1 U718 ( .A1(n608), .A2(n607), .ZN(n643) );
  AND2_X1 U719 ( .A1(n609), .A2(n643), .ZN(n610) );
  NAND2_X1 U720 ( .A1(n611), .A2(n610), .ZN(n680) );
  NAND2_X1 U721 ( .A1(n612), .A2(n680), .ZN(n613) );
  XNOR2_X1 U722 ( .A(n613), .B(KEYINPUT83), .ZN(n616) );
  NAND2_X1 U723 ( .A1(KEYINPUT47), .A2(n614), .ZN(n615) );
  XOR2_X1 U724 ( .A(KEYINPUT48), .B(KEYINPUT70), .Z(n619) );
  NAND2_X1 U725 ( .A1(n686), .A2(n621), .ZN(n693) );
  NOR2_X1 U726 ( .A1(G898), .A2(n622), .ZN(n763) );
  NAND2_X1 U727 ( .A1(G902), .A2(n763), .ZN(n624) );
  NAND2_X1 U728 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U729 ( .A(n651), .ZN(n641) );
  INV_X1 U730 ( .A(n713), .ZN(n632) );
  AND2_X1 U731 ( .A1(n637), .A2(n694), .ZN(n635) );
  NAND2_X1 U732 ( .A1(n698), .A2(n635), .ZN(n636) );
  NOR2_X1 U733 ( .A1(n675), .A2(n353), .ZN(n656) );
  NOR2_X1 U734 ( .A1(n700), .A2(n644), .ZN(n645) );
  XNOR2_X1 U735 ( .A(n645), .B(KEYINPUT92), .ZN(n646) );
  NAND2_X1 U736 ( .A1(n646), .A2(n638), .ZN(n666) );
  NOR2_X1 U737 ( .A1(n647), .A2(n641), .ZN(n648) );
  NAND2_X1 U738 ( .A1(n365), .A2(n648), .ZN(n649) );
  NOR2_X1 U739 ( .A1(n698), .A2(n650), .ZN(n705) );
  NAND2_X1 U740 ( .A1(n425), .A2(n705), .ZN(n652) );
  XNOR2_X1 U741 ( .A(n652), .B(KEYINPUT31), .ZN(n687) );
  NOR2_X1 U742 ( .A1(n672), .A2(n687), .ZN(n653) );
  INV_X1 U743 ( .A(KEYINPUT63), .ZN(n664) );
  XNOR2_X1 U744 ( .A(G101), .B(n666), .ZN(G3) );
  XOR2_X1 U745 ( .A(G104), .B(KEYINPUT111), .Z(n668) );
  NAND2_X1 U746 ( .A1(n672), .A2(n683), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n668), .B(n667), .ZN(G6) );
  XOR2_X1 U748 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n670) );
  XNOR2_X1 U749 ( .A(G107), .B(KEYINPUT112), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U751 ( .A(KEYINPUT26), .B(n671), .Z(n674) );
  NAND2_X1 U752 ( .A1(n672), .A2(n686), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n674), .B(n673), .ZN(G9) );
  XOR2_X1 U754 ( .A(n675), .B(G110), .Z(G12) );
  XOR2_X1 U755 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n677) );
  NAND2_X1 U756 ( .A1(n686), .A2(n681), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U758 ( .A(G128), .B(n678), .ZN(G30) );
  XOR2_X1 U759 ( .A(G143), .B(KEYINPUT115), .Z(n679) );
  XNOR2_X1 U760 ( .A(n680), .B(n679), .ZN(G45) );
  NAND2_X1 U761 ( .A1(n681), .A2(n683), .ZN(n682) );
  XNOR2_X1 U762 ( .A(n682), .B(G146), .ZN(G48) );
  NAND2_X1 U763 ( .A1(n687), .A2(n683), .ZN(n684) );
  XNOR2_X1 U764 ( .A(n684), .B(KEYINPUT116), .ZN(n685) );
  XNOR2_X1 U765 ( .A(G113), .B(n685), .ZN(G15) );
  XOR2_X1 U766 ( .A(G116), .B(KEYINPUT117), .Z(n689) );
  NAND2_X1 U767 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U768 ( .A(n689), .B(n688), .ZN(G18) );
  XNOR2_X1 U769 ( .A(n690), .B(KEYINPUT118), .ZN(n691) );
  XNOR2_X1 U770 ( .A(n691), .B(KEYINPUT37), .ZN(n692) );
  XNOR2_X1 U771 ( .A(G125), .B(n692), .ZN(G27) );
  XNOR2_X1 U772 ( .A(G134), .B(n693), .ZN(G36) );
  AND2_X1 U773 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U774 ( .A(n696), .B(KEYINPUT49), .ZN(n697) );
  NAND2_X1 U775 ( .A1(n698), .A2(n697), .ZN(n703) );
  NOR2_X1 U776 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U777 ( .A(n701), .B(KEYINPUT50), .ZN(n702) );
  NOR2_X1 U778 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U779 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U780 ( .A(KEYINPUT119), .B(n706), .Z(n707) );
  XOR2_X1 U781 ( .A(KEYINPUT51), .B(n707), .Z(n708) );
  NOR2_X1 U782 ( .A1(n733), .A2(n708), .ZN(n720) );
  NOR2_X1 U783 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U784 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U787 ( .A1(n734), .A2(n718), .ZN(n719) );
  NOR2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U789 ( .A(n721), .B(KEYINPUT52), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U791 ( .A1(G952), .A2(n724), .ZN(n732) );
  NAND2_X1 U792 ( .A1(n769), .A2(n438), .ZN(n725) );
  XNOR2_X1 U793 ( .A(KEYINPUT87), .B(n725), .ZN(n728) );
  BUF_X1 U794 ( .A(n726), .Z(n727) );
  NOR2_X1 U795 ( .A1(n728), .A2(n493), .ZN(n729) );
  NAND2_X1 U796 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U797 ( .A(KEYINPUT53), .B(n735), .ZN(G75) );
  XNOR2_X1 U798 ( .A(KEYINPUT55), .B(KEYINPUT84), .ZN(n739) );
  BUF_X1 U799 ( .A(n736), .Z(n737) );
  XNOR2_X1 U800 ( .A(n737), .B(KEYINPUT54), .ZN(n738) );
  XOR2_X1 U801 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n744) );
  INV_X1 U802 ( .A(KEYINPUT59), .ZN(n745) );
  NOR2_X1 U803 ( .A1(n754), .A2(n752), .ZN(G63) );
  OR2_X1 U804 ( .A1(n727), .A2(G953), .ZN(n759) );
  NAND2_X1 U805 ( .A1(G224), .A2(G953), .ZN(n755) );
  XNOR2_X1 U806 ( .A(n755), .B(KEYINPUT61), .ZN(n756) );
  XNOR2_X1 U807 ( .A(KEYINPUT124), .B(n756), .ZN(n757) );
  NAND2_X1 U808 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U809 ( .A1(n759), .A2(n758), .ZN(n765) );
  BUF_X1 U810 ( .A(n760), .Z(n761) );
  XOR2_X1 U811 ( .A(n761), .B(KEYINPUT125), .Z(n762) );
  NOR2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U813 ( .A(n765), .B(n764), .ZN(G69) );
  XOR2_X1 U814 ( .A(n766), .B(KEYINPUT126), .Z(n767) );
  XNOR2_X1 U815 ( .A(n768), .B(n767), .ZN(n771) );
  XNOR2_X1 U816 ( .A(n771), .B(n769), .ZN(n770) );
  NAND2_X1 U817 ( .A1(n770), .A2(n497), .ZN(n776) );
  XNOR2_X1 U818 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U819 ( .A1(n772), .A2(G900), .ZN(n773) );
  XOR2_X1 U820 ( .A(KEYINPUT127), .B(n773), .Z(n774) );
  NAND2_X1 U821 ( .A1(G953), .A2(n774), .ZN(n775) );
  NAND2_X1 U822 ( .A1(n776), .A2(n775), .ZN(G72) );
  XNOR2_X1 U823 ( .A(G122), .B(n777), .ZN(G24) );
  XOR2_X1 U824 ( .A(G140), .B(n778), .Z(G42) );
  XOR2_X1 U825 ( .A(n779), .B(G119), .Z(G21) );
  XOR2_X1 U826 ( .A(n780), .B(G131), .Z(G33) );
  XOR2_X1 U827 ( .A(n781), .B(G137), .Z(G39) );
endmodule

