//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1203,
    new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n465), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  OR2_X1    g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n470), .A2(new_n472), .B1(new_n478), .B2(G2105), .ZN(G160));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n475), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT69), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n474), .A2(new_n482), .A3(new_n475), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n462), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n462), .A3(new_n483), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(new_n467), .A2(G102), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n480), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(new_n462), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n497), .B(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT70), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n497), .B(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(G114), .A2(G2104), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n463), .A2(new_n464), .ZN(new_n503));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G2105), .B1(G102), .B2(new_n467), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n501), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n500), .A2(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n514), .A2(new_n516), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n511), .A2(new_n512), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n514), .A2(new_n516), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT71), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n514), .A2(new_n516), .A3(new_n528), .A4(G62), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n523), .B1(new_n530), .B2(G651), .ZN(G166));
  INV_X1    g106(.A(new_n521), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n514), .A2(new_n516), .A3(G63), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(G89), .B1(G651), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n510), .A2(G51), .A3(G543), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n514), .A2(new_n516), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n540), .A2(G89), .A3(new_n510), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n514), .A2(new_n516), .A3(G63), .A4(G651), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n541), .A2(new_n536), .A3(new_n542), .A4(new_n538), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT72), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n539), .A2(new_n544), .ZN(G168));
  NAND3_X1  g120(.A1(new_n514), .A2(new_n516), .A3(G64), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  NOR3_X1   g125(.A1(new_n549), .A2(new_n550), .A3(new_n517), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n511), .A2(new_n552), .B1(new_n521), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  INV_X1    g131(.A(G68), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n524), .A2(new_n556), .B1(new_n557), .B2(new_n513), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI221_X1 g135(.A(KEYINPUT74), .B1(new_n557), .B2(new_n513), .C1(new_n524), .C2(new_n556), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G651), .A3(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n510), .A2(G543), .ZN(new_n563));
  AOI22_X1  g138(.A1(G43), .A2(new_n563), .B1(new_n532), .B2(G81), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(G188));
  NAND4_X1  g146(.A1(new_n518), .A2(new_n520), .A3(G53), .A4(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n510), .A2(new_n574), .A3(G53), .A4(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n524), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n532), .A2(G91), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(new_n580), .A3(new_n581), .ZN(G299));
  NOR3_X1   g157(.A1(new_n551), .A2(KEYINPUT75), .A3(new_n554), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n546), .A2(new_n548), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT73), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(G651), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n554), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G301));
  INV_X1    g167(.A(G168), .ZN(G286));
  NAND2_X1  g168(.A1(new_n530), .A2(G651), .ZN(new_n594));
  INV_X1    g169(.A(new_n523), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G303));
  INV_X1    g171(.A(G87), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT76), .B1(new_n521), .B2(new_n597), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n598), .A2(new_n599), .B1(G49), .B2(new_n563), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n540), .B2(G74), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G288));
  NAND2_X1  g177(.A1(new_n540), .A2(G61), .ZN(new_n603));
  NAND2_X1  g178(.A1(G73), .A2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT77), .Z(new_n605));
  AOI21_X1  g180(.A(new_n517), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G48), .ZN(new_n607));
  INV_X1    g182(.A(G86), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n511), .A2(new_n607), .B1(new_n521), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G305));
  NAND3_X1  g186(.A1(new_n514), .A2(new_n516), .A3(G60), .ZN(new_n612));
  NAND2_X1  g187(.A1(G72), .A2(G543), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT78), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n612), .A2(new_n616), .A3(new_n613), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n615), .A2(G651), .A3(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(G47), .A2(new_n563), .B1(new_n532), .B2(G85), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G66), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n524), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G651), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G92), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n521), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n563), .A2(G54), .ZN(new_n629));
  NAND4_X1  g204(.A1(new_n540), .A2(new_n625), .A3(G92), .A4(new_n510), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n624), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n591), .B2(new_n632), .ZN(G284));
  OAI21_X1  g209(.A(new_n633), .B1(new_n591), .B2(new_n632), .ZN(G321));
  NAND2_X1  g210(.A1(G299), .A2(new_n632), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G168), .B2(new_n632), .ZN(G280));
  XNOR2_X1  g212(.A(G280), .B(KEYINPUT80), .ZN(G297));
  INV_X1    g213(.A(new_n631), .ZN(new_n639));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G860), .ZN(G148));
  NOR2_X1   g216(.A1(new_n565), .A2(G868), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(G868), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT82), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g222(.A1(new_n485), .A2(G123), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n488), .A2(G135), .ZN(new_n649));
  NOR2_X1   g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n480), .A2(new_n467), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT13), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2435), .ZN(new_n661));
  XOR2_X1   g236(.A(G2427), .B(G2438), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT14), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2451), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1341), .B(G1348), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(G14), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  INV_X1    g255(.A(new_n678), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(KEYINPUT17), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n675), .A2(new_n676), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(KEYINPUT17), .ZN(new_n684));
  NAND4_X1  g259(.A1(new_n682), .A2(new_n683), .A3(new_n677), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n678), .B(KEYINPUT85), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n680), .B(new_n685), .C1(new_n683), .C2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2096), .ZN(new_n690));
  INV_X1    g265(.A(G2100), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n697), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n695), .A2(new_n698), .A3(new_n700), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n703), .B(new_n704), .C1(new_n701), .C2(new_n702), .ZN(new_n705));
  XOR2_X1   g280(.A(G1991), .B(G1996), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(G229));
  INV_X1    g286(.A(G107), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n466), .B1(new_n712), .B2(G2105), .ZN(new_n713));
  OR2_X1    g288(.A1(G95), .A2(G2105), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT88), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n717), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n481), .A2(G119), .A3(G2105), .A4(new_n483), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n481), .A2(G131), .A3(new_n462), .A4(new_n483), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G25), .B(new_n722), .S(G29), .Z(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT35), .B(G1991), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n723), .B(new_n724), .Z(new_n725));
  INV_X1    g300(.A(G1986), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n618), .A2(new_n619), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(G24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n725), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(G23), .ZN(new_n732));
  INV_X1    g307(.A(G288), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n728), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT33), .ZN(new_n735));
  INV_X1    g310(.A(G1976), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n728), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n728), .ZN(new_n740));
  INV_X1    g315(.A(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n728), .A2(G6), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n610), .B2(new_n728), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT32), .B(G1981), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n737), .A2(new_n738), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n731), .B1(new_n747), .B2(KEYINPUT34), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n730), .A2(new_n726), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n748), .B(new_n749), .C1(KEYINPUT34), .C2(new_n747), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT36), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G26), .ZN(new_n753));
  INV_X1    g328(.A(G116), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n466), .B1(new_n754), .B2(G2105), .ZN(new_n755));
  OR2_X1    g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT89), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n755), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n481), .A2(G128), .A3(G2105), .A4(new_n483), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n481), .A2(G140), .A3(new_n462), .A4(new_n483), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(KEYINPUT90), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n753), .B1(new_n769), .B2(new_n752), .ZN(new_n770));
  MUX2_X1   g345(.A(new_n753), .B(new_n770), .S(KEYINPUT28), .Z(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(G2067), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n752), .A2(KEYINPUT94), .A3(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n752), .ZN(new_n774));
  AOI21_X1  g349(.A(KEYINPUT94), .B1(new_n752), .B2(G27), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT95), .B(G2078), .Z(new_n777));
  AND2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G1341), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n565), .A2(new_n728), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n728), .B2(G19), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n776), .A2(new_n777), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n778), .B(new_n782), .C1(new_n779), .C2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n728), .A2(G20), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT97), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT23), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G16), .B2(G299), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  NOR2_X1   g363(.A1(G29), .A2(G32), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n467), .A2(G105), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT91), .Z(new_n791));
  NAND4_X1  g366(.A1(new_n481), .A2(G141), .A3(new_n462), .A4(new_n483), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n481), .A2(G129), .A3(G2105), .A4(new_n483), .ZN(new_n793));
  NAND3_X1  g368(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT26), .Z(new_n795));
  NAND4_X1  g370(.A1(new_n791), .A2(new_n792), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n789), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT27), .B(G1996), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(KEYINPUT24), .A2(G34), .ZN(new_n801));
  NAND2_X1  g376(.A1(KEYINPUT24), .A2(G34), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n801), .A2(new_n752), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G160), .B2(new_n752), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G2084), .ZN(new_n805));
  NAND2_X1  g380(.A1(G171), .A2(G16), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G5), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1961), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n788), .A2(new_n800), .A3(new_n805), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n467), .A2(G103), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT25), .Z(new_n812));
  AOI22_X1  g387(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n813));
  INV_X1    g388(.A(G139), .ZN(new_n814));
  OAI221_X1 g389(.A(new_n812), .B1(new_n462), .B2(new_n813), .C1(new_n814), .C2(new_n487), .ZN(new_n815));
  MUX2_X1   g390(.A(G33), .B(new_n815), .S(G29), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2072), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n728), .A2(G4), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n639), .B2(new_n728), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1348), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n798), .A2(new_n799), .B1(new_n804), .B2(G2084), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n810), .A2(new_n817), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n752), .A2(G35), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G162), .B2(new_n752), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT96), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT29), .B(G2090), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n783), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G28), .ZN(new_n829));
  AOI21_X1  g404(.A(G29), .B1(new_n829), .B2(KEYINPUT30), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(KEYINPUT30), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n652), .B2(new_n752), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n807), .A2(new_n808), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n728), .A2(G21), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G168), .B2(new_n728), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n832), .B(new_n833), .C1(G1966), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(G1966), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT92), .Z(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT31), .B(G11), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT93), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(KEYINPUT93), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n771), .A2(G2067), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n828), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n751), .A2(new_n772), .A3(new_n844), .ZN(G150));
  INV_X1    g420(.A(G150), .ZN(G311));
  AOI22_X1  g421(.A1(new_n540), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n517), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  INV_X1    g424(.A(G93), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n511), .A2(new_n849), .B1(new_n521), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n565), .B(new_n852), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT39), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n639), .A2(G559), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT38), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n857), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n855), .B1(new_n860), .B2(G860), .ZN(G145));
  NAND2_X1  g436(.A1(new_n501), .A2(new_n506), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n766), .A2(new_n767), .A3(new_n796), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n796), .B1(new_n766), .B2(new_n767), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n768), .A2(new_n797), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n496), .A2(new_n499), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n868), .A3(new_n863), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n815), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n866), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n815), .A2(new_n870), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n866), .A2(new_n869), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n488), .A2(KEYINPUT101), .A3(G142), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n485), .A2(G130), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  INV_X1    g458(.A(G142), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n487), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n879), .A2(new_n880), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n887));
  INV_X1    g462(.A(new_n656), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n888), .B1(new_n887), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n886), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n887), .A2(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n656), .ZN(new_n896));
  INV_X1    g471(.A(new_n886), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n492), .B(KEYINPUT98), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n894), .A2(new_n898), .A3(KEYINPUT103), .A4(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n878), .A2(new_n901), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n866), .A2(new_n869), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n873), .A2(new_n876), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n901), .A2(new_n910), .A3(new_n874), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n652), .B(G160), .Z(new_n913));
  AND3_X1   g488(.A1(new_n906), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n906), .B2(new_n912), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g494(.A1(new_n853), .A2(new_n632), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n727), .A2(G303), .ZN(new_n921));
  NAND2_X1  g496(.A1(G290), .A2(G166), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n921), .A2(new_n922), .A3(G305), .ZN(new_n923));
  AOI21_X1  g498(.A(G305), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G288), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n610), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n921), .A2(new_n922), .A3(G305), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n733), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n856), .B(new_n643), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n631), .B(G299), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n639), .A2(G299), .ZN(new_n936));
  INV_X1    g511(.A(G299), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(new_n631), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT104), .B1(new_n639), .B2(G299), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n933), .B2(KEYINPUT104), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n942), .B2(new_n939), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n935), .B1(new_n932), .B2(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n931), .B(new_n944), .Z(new_n945));
  OAI21_X1  g520(.A(new_n920), .B1(new_n945), .B2(new_n632), .ZN(G295));
  OAI21_X1  g521(.A(new_n920), .B1(new_n945), .B2(new_n632), .ZN(G331));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n949));
  OAI21_X1  g524(.A(G168), .B1(new_n583), .B2(new_n590), .ZN(new_n950));
  NAND3_X1  g525(.A1(G171), .A2(new_n539), .A3(new_n544), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND4_X1   g527(.A1(new_n539), .A2(new_n544), .A3(new_n589), .A4(new_n588), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(KEYINPUT106), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n952), .A2(new_n856), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n565), .B(new_n853), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT75), .B1(new_n551), .B2(new_n554), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n588), .A2(new_n589), .A3(new_n584), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n957), .A2(new_n958), .B1(new_n539), .B2(new_n544), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT106), .B1(new_n959), .B2(new_n953), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n951), .A2(new_n949), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n933), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n856), .B1(new_n952), .B2(new_n954), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n956), .A3(new_n961), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n943), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n930), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n948), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(KEYINPUT107), .B(new_n930), .C1(new_n963), .C2(new_n966), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT41), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n933), .ZN(new_n973));
  INV_X1    g548(.A(new_n942), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n973), .B(new_n930), .C1(new_n974), .C2(new_n972), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n971), .A2(new_n917), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n964), .A2(new_n943), .A3(new_n965), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n934), .B1(new_n964), .B2(new_n965), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n968), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT107), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n967), .A2(new_n948), .A3(new_n968), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n963), .A2(new_n930), .A3(new_n966), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .A4(new_n917), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n976), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n978), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(KEYINPUT44), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n971), .A2(new_n917), .A3(new_n975), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n985), .B2(new_n976), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(KEYINPUT44), .B2(new_n991), .ZN(G397));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n500), .A2(new_n508), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(G160), .A2(KEYINPUT108), .A3(G40), .ZN(new_n996));
  OAI21_X1  g571(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n997));
  INV_X1    g572(.A(new_n472), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n471), .B1(new_n465), .B2(new_n468), .ZN(new_n999));
  OAI211_X1 g574(.A(G40), .B(new_n997), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n995), .A2(KEYINPUT50), .B1(new_n996), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G2090), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n862), .A2(new_n994), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1006));
  OR2_X1    g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n995), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1005), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n996), .A2(new_n1002), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1008), .A2(new_n1009), .B1(new_n741), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n993), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(G166), .A2(new_n993), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT55), .Z(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT112), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n993), .B1(new_n1015), .B2(new_n1013), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(G288), .B2(new_n736), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n733), .A2(KEYINPUT113), .A3(G1976), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT52), .ZN(new_n1028));
  INV_X1    g603(.A(G1981), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n610), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT49), .B1(new_n610), .B2(new_n1029), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n610), .A2(new_n1029), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1033), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n1036), .A3(new_n1031), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1023), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n736), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1028), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1022), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1015), .B(new_n1043), .C1(new_n1011), .C2(new_n995), .ZN(new_n1044));
  INV_X1    g619(.A(G1966), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G2084), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1003), .A2(new_n1047), .A3(new_n1007), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n993), .B(G286), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1020), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1018), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT63), .B1(new_n1051), .B2(new_n1041), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1041), .A2(KEYINPUT116), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1028), .A2(new_n1054), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n500), .A2(new_n508), .A3(new_n1057), .A4(new_n994), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1015), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1060), .A2(KEYINPUT115), .ZN(new_n1061));
  AOI21_X1  g636(.A(G2090), .B1(new_n1060), .B2(KEYINPUT115), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1061), .A2(new_n1062), .B1(new_n741), .B2(new_n1016), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1020), .B1(new_n1063), .B2(new_n993), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT63), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1049), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1056), .A2(new_n1022), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1038), .A2(new_n736), .A3(new_n733), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1034), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1023), .ZN(new_n1070));
  AND4_X1   g645(.A1(new_n1042), .A2(new_n1052), .A3(new_n1067), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT123), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1074));
  OAI211_X1 g649(.A(G8), .B(new_n1073), .C1(new_n1074), .C2(G286), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1072), .A2(KEYINPUT123), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(G8), .A3(G286), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT62), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1056), .A2(new_n1064), .A3(new_n1022), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n995), .A2(KEYINPUT50), .ZN(new_n1084));
  AND4_X1   g659(.A1(KEYINPUT118), .A2(new_n1084), .A3(new_n1007), .A4(new_n1015), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT118), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n808), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(G2078), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1087), .B(KEYINPUT124), .C1(new_n1089), .C2(new_n1044), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1088), .B1(new_n1016), .B2(G2078), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1084), .A2(new_n1007), .A3(new_n1015), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1003), .A2(KEYINPUT118), .A3(new_n1007), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1961), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1044), .A2(new_n1089), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1092), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1090), .A2(new_n1091), .A3(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1100), .A2(new_n591), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1077), .A2(new_n1102), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1081), .A2(new_n1083), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1087), .A2(KEYINPUT125), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1097), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1000), .B1(new_n1013), .B2(KEYINPUT45), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1088), .A2(G2078), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1043), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1091), .A2(new_n1110), .ZN(new_n1111));
  AND4_X1   g686(.A1(G301), .A2(new_n1105), .A3(new_n1107), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n591), .B2(new_n1100), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(G1996), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1015), .A2(new_n1013), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT58), .B(G1341), .Z(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n565), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT59), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1122), .A3(new_n565), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1956), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1060), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT57), .B1(new_n576), .B2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(G299), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1126), .A2(new_n1128), .A3(new_n1134), .A4(new_n1131), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1133), .A2(KEYINPUT61), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1132), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1131), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1124), .A2(new_n1136), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1348), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1143));
  INV_X1    g718(.A(G2067), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1015), .A2(new_n1144), .A3(new_n1013), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n639), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1143), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT60), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n639), .A2(new_n1147), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1141), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n639), .A3(new_n1132), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT119), .Z(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1158), .B2(new_n1131), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1113), .A2(KEYINPUT54), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1105), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(G171), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1162), .B(KEYINPUT54), .C1(new_n1100), .C2(new_n591), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(new_n1083), .A3(new_n1080), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1071), .B(new_n1104), .C1(new_n1160), .C2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1043), .B1(new_n1002), .B2(new_n996), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n722), .B(new_n724), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT109), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n768), .B(new_n1144), .ZN(new_n1169));
  INV_X1    g744(.A(G1996), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n796), .B(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(G290), .B(G1986), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1166), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1165), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1166), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n722), .A2(new_n724), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT126), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1169), .A2(new_n1171), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n769), .A2(new_n1144), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1177), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT46), .Z(new_n1184));
  AOI21_X1  g759(.A(new_n1177), .B1(new_n1169), .B2(new_n797), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT47), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1173), .A2(new_n1166), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1166), .A2(new_n726), .A3(new_n727), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT48), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1182), .B(new_n1187), .C1(new_n1188), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1176), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(G319), .ZN(new_n1194));
  OR2_X1    g768(.A1(G229), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g769(.A(new_n1195), .ZN(new_n1196));
  OAI21_X1  g770(.A(new_n692), .B1(new_n673), .B2(new_n672), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n916), .B2(new_n917), .ZN(new_n1198));
  AND4_X1   g772(.A1(KEYINPUT127), .A2(new_n987), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n978), .B2(new_n986), .ZN(new_n1200));
  AOI21_X1  g774(.A(KEYINPUT127), .B1(new_n1200), .B2(new_n1198), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n1199), .A2(new_n1201), .ZN(G308));
  NAND3_X1  g776(.A1(new_n987), .A2(new_n1198), .A3(new_n1196), .ZN(new_n1203));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g779(.A1(new_n1200), .A2(KEYINPUT127), .A3(new_n1198), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1206), .ZN(G225));
endmodule


