//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT72), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n195), .A2(G227), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n194), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(G128), .A3(new_n200), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT10), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT74), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G104), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(KEYINPUT73), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT73), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G107), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n213), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(G104), .B1(new_n217), .B2(new_n219), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT74), .B(G101), .C1(new_n225), .C2(new_n216), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT73), .B(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n214), .B2(G104), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n215), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n232), .A3(new_n223), .ZN(new_n233));
  AND4_X1   g047(.A1(KEYINPUT75), .A2(new_n224), .A3(new_n226), .A4(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(G101), .B1(new_n225), .B2(new_n216), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n227), .A2(new_n228), .B1(new_n231), .B2(new_n215), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n235), .A2(new_n213), .B1(new_n236), .B2(new_n223), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT75), .B1(new_n237), .B2(new_n226), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n212), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G131), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(KEYINPUT65), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G134), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n248), .B2(G137), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(G137), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n241), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n242), .A2(G134), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n243), .B2(new_n246), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n248), .A2(G137), .ZN(new_n255));
  INV_X1    g069(.A(new_n246), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(new_n244), .ZN(new_n257));
  INV_X1    g071(.A(new_n241), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n236), .A2(new_n223), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n229), .A2(new_n232), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G101), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n207), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n205), .A2(KEYINPUT0), .A3(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n224), .A2(new_n209), .A3(new_n226), .A4(new_n233), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n264), .A2(new_n273), .B1(new_n274), .B2(new_n211), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n239), .A2(new_n261), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n261), .B1(new_n239), .B2(new_n275), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n198), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n197), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n224), .A2(new_n226), .A3(new_n233), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n237), .A2(KEYINPUT75), .A3(new_n226), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n210), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n274), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n260), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT12), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(KEYINPUT12), .A3(new_n260), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n280), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n279), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n276), .A2(new_n197), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n288), .B(new_n261), .C1(new_n285), .C2(new_n274), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT12), .B1(new_n286), .B2(new_n260), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n294), .B(new_n292), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n192), .B(new_n190), .C1(new_n293), .C2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n192), .A2(new_n190), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n280), .A2(new_n278), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n276), .B1(new_n296), .B2(new_n295), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(new_n198), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n303), .B2(G469), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n191), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT16), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(G125), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n310), .B1(new_n314), .B2(new_n308), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n202), .ZN(new_n316));
  OAI211_X1 g130(.A(G146), .B(new_n310), .C1(new_n314), .C2(new_n308), .ZN(new_n317));
  NOR2_X1   g131(.A1(G237), .A2(G953), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n318), .A2(G143), .A3(G214), .ZN(new_n319));
  AOI21_X1  g133(.A(G143), .B1(new_n318), .B2(G214), .ZN(new_n320));
  OAI211_X1 g134(.A(KEYINPUT17), .B(G131), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G131), .B1(new_n319), .B2(new_n320), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT17), .ZN(new_n324));
  INV_X1    g138(.A(G237), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n195), .A3(G214), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n199), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n318), .A2(G143), .A3(G214), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n240), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n323), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT86), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT86), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n323), .A2(new_n329), .A3(new_n332), .A4(new_n324), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n322), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n327), .A2(new_n328), .ZN(new_n335));
  NAND2_X1  g149(.A1(KEYINPUT18), .A2(G131), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n335), .B(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n311), .A2(new_n313), .A3(new_n202), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT70), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n314), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT81), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(G146), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n334), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G113), .B(G122), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT85), .B(G104), .ZN(new_n348));
  XOR2_X1   g162(.A(new_n347), .B(new_n348), .Z(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n345), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n323), .A2(new_n329), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(KEYINPUT19), .A3(new_n342), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n356), .A2(KEYINPUT19), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(KEYINPUT19), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n357), .A2(new_n311), .A3(new_n313), .A4(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n202), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT83), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n355), .A2(new_n362), .A3(new_n202), .A4(new_n359), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n317), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n354), .B1(new_n364), .B2(KEYINPUT84), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n361), .A2(new_n366), .A3(new_n317), .A4(new_n363), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n353), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n352), .B1(new_n368), .B2(new_n349), .ZN(new_n369));
  NOR2_X1   g183(.A1(G475), .A2(G902), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n307), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n346), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n334), .A2(new_n345), .A3(KEYINPUT88), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n373), .A2(KEYINPUT89), .A3(new_n350), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n352), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n349), .B1(new_n346), .B2(new_n372), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT89), .B1(new_n377), .B2(new_n374), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n190), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n306), .A2(new_n371), .B1(new_n379), .B2(G475), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n199), .A2(G128), .ZN(new_n381));
  INV_X1    g195(.A(G128), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G143), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n384), .A2(KEYINPUT93), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(KEYINPUT93), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT92), .ZN(new_n388));
  INV_X1    g202(.A(new_n381), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(KEYINPUT13), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n199), .A2(G128), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n381), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n248), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n393), .A2(KEYINPUT92), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n248), .A2(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G122), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G116), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G116), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G122), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(KEYINPUT91), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT91), .B1(new_n400), .B2(new_n402), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n404), .A2(new_n405), .A3(new_n227), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n400), .A2(new_n402), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT91), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n220), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n396), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n227), .B1(new_n404), .B2(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n387), .A2(new_n248), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n385), .A2(G134), .A3(new_n386), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n400), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n418), .A2(new_n419), .A3(G107), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n418), .B2(G107), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n412), .B(new_n415), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n411), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n189), .A2(G217), .A3(new_n195), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n424), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n411), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G478), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n429), .A2(KEYINPUT15), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n428), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n364), .A2(KEYINPUT84), .ZN(new_n433));
  INV_X1    g247(.A(new_n354), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n367), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n345), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n351), .B1(new_n436), .B2(new_n350), .ZN(new_n437));
  INV_X1    g251(.A(new_n370), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT87), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n369), .A2(new_n307), .A3(new_n370), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(KEYINPUT20), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n380), .A2(new_n432), .A3(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n305), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n401), .A2(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n401), .A2(G119), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT2), .B(G113), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n445), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT30), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT66), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n454), .A2(KEYINPUT66), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n254), .A2(new_n257), .A3(new_n240), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n240), .B1(new_n243), .B2(new_n250), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n209), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n252), .A2(new_n259), .B1(new_n271), .B2(new_n270), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n455), .B(new_n456), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n260), .A2(new_n272), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n458), .B1(new_n206), .B2(new_n208), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n457), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n463), .A2(KEYINPUT66), .A3(new_n465), .A4(new_n454), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n453), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n460), .A2(new_n461), .A3(new_n452), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n318), .A2(G210), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT27), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT26), .B(G101), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n467), .A2(new_n468), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n474), .B2(KEYINPUT31), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n466), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n452), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n463), .A2(new_n453), .A3(new_n465), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n472), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT31), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT28), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n478), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n460), .A2(new_n461), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT28), .B1(new_n484), .B2(new_n453), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n473), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n479), .A2(new_n480), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G472), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n475), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT32), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n475), .A2(new_n487), .A3(new_n491), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n494));
  NOR4_X1   g308(.A1(new_n483), .A2(new_n485), .A3(new_n494), .A4(new_n473), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT67), .B1(new_n495), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT67), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n478), .A2(new_n481), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n482), .A2(new_n478), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n472), .B(new_n498), .C1(new_n499), .C2(new_n481), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n497), .B(new_n190), .C1(new_n500), .C2(new_n494), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n473), .B1(new_n467), .B2(new_n468), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n502), .A3(new_n494), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G472), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n493), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n507));
  INV_X1    g321(.A(G234), .ZN(new_n508));
  OAI21_X1  g322(.A(G217), .B1(new_n508), .B2(G902), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT68), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT23), .B1(new_n382), .B2(G119), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT69), .B1(new_n382), .B2(G119), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G119), .B(G128), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT24), .B(G110), .Z(new_n515));
  OAI22_X1  g329(.A1(new_n513), .A2(G110), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n317), .A3(new_n339), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n513), .A2(G110), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n316), .A2(new_n317), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT22), .B(G137), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n187), .A2(new_n508), .A3(G953), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n522), .B(new_n523), .Z(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n517), .A2(new_n520), .A3(new_n524), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n528), .B2(G902), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n510), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n509), .A2(new_n190), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n506), .A2(new_n507), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n490), .A2(new_n492), .B1(new_n504), .B2(G472), .ZN(new_n538));
  INV_X1    g352(.A(new_n536), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT71), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(G952), .B(new_n195), .C1(new_n508), .C2(new_n325), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT95), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(G902), .B(G953), .C1(new_n508), .C2(new_n325), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT96), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT21), .B(G898), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G214), .B1(G237), .B2(G902), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n272), .A2(G125), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n210), .B2(G125), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n195), .A2(G224), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT7), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n552), .B(new_n554), .Z(new_n555));
  NAND2_X1  g369(.A1(new_n446), .A2(KEYINPUT5), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n556), .B(G113), .C1(KEYINPUT5), .C2(new_n444), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n557), .A2(new_n449), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n234), .B2(new_n238), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G122), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n262), .A2(new_n263), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n452), .A2(new_n267), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT78), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n283), .A2(new_n284), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(new_n567), .B2(new_n558), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n560), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n555), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n560), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n557), .A2(new_n449), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n283), .B2(new_n284), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n573), .A2(new_n281), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT80), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(new_n572), .C1(new_n574), .C2(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n571), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT6), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n559), .A2(new_n564), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n560), .B(KEYINPUT77), .Z(new_n584));
  AOI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n569), .B1(new_n568), .B2(new_n560), .ZN(new_n586));
  INV_X1    g400(.A(new_n560), .ZN(new_n587));
  NOR4_X1   g401(.A1(new_n574), .A2(KEYINPUT78), .A3(new_n587), .A4(new_n563), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n585), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n552), .B(new_n553), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n582), .B(new_n584), .C1(new_n574), .C2(new_n563), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT79), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT79), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n583), .A2(new_n593), .A3(new_n582), .A4(new_n584), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n589), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(G210), .B1(G237), .B2(G902), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n581), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n581), .B2(new_n596), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n549), .B(new_n550), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n443), .A2(new_n541), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  OAI21_X1  g417(.A(new_n550), .B1(new_n598), .B2(new_n599), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(KEYINPUT97), .B(new_n550), .C1(new_n598), .C2(new_n599), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n380), .A2(new_n441), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n425), .A2(new_n427), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n427), .B2(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n425), .B(new_n427), .C1(KEYINPUT98), .C2(new_n611), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(G478), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n429), .A2(new_n190), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n428), .B2(new_n429), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n299), .A2(new_n304), .ZN(new_n620));
  INV_X1    g434(.A(new_n191), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n475), .A2(new_n487), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n489), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n539), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n608), .A2(new_n549), .A3(new_n619), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  NAND3_X1  g443(.A1(new_n380), .A2(new_n431), .A3(new_n441), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n608), .A2(new_n549), .A3(new_n626), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n530), .A2(new_n532), .ZN(new_n635));
  INV_X1    g449(.A(new_n510), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n525), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n521), .B(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n534), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n624), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n443), .A2(new_n601), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT99), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT37), .B(G110), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  NOR2_X1   g462(.A1(new_n538), .A2(new_n643), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n649), .A2(new_n305), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n608), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT100), .B(G900), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n546), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n543), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n380), .A2(new_n431), .A3(new_n441), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n382), .ZN(G30));
  XNOR2_X1  g474(.A(new_n657), .B(KEYINPUT39), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n305), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n477), .A2(new_n478), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n472), .ZN(new_n665));
  AOI21_X1  g479(.A(G902), .B1(new_n499), .B2(new_n473), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n493), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(KEYINPUT102), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n380), .A2(new_n441), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n671), .A2(new_n550), .A3(new_n431), .A4(new_n643), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT103), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n581), .A2(new_n596), .ZN(new_n674));
  INV_X1    g488(.A(new_n597), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n581), .A2(new_n596), .A3(new_n597), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n670), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n672), .A2(KEYINPUT103), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n663), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT104), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  INV_X1    g498(.A(new_n657), .ZN(new_n685));
  AOI211_X1 g499(.A(new_n685), .B(new_n618), .C1(new_n380), .C2(new_n441), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n608), .A2(new_n650), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT105), .B(G146), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G48));
  AOI21_X1  g503(.A(KEYINPUT97), .B1(new_n678), .B2(new_n550), .ZN(new_n690));
  INV_X1    g504(.A(new_n607), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n549), .B(new_n619), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n190), .B1(new_n293), .B2(new_n298), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n694), .A2(new_n621), .A3(new_n299), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n539), .B1(new_n493), .B2(new_n505), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT106), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n698), .B(new_n700), .ZN(G15));
  OAI211_X1 g515(.A(new_n549), .B(new_n631), .C1(new_n690), .C2(new_n691), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n697), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n401), .ZN(G18));
  OAI21_X1  g518(.A(new_n695), .B1(new_n690), .B2(new_n691), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n608), .A2(new_n707), .A3(new_n695), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n649), .A2(new_n549), .A3(new_n442), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NAND3_X1  g526(.A1(new_n694), .A2(new_n621), .A3(new_n299), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT108), .B(G472), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n622), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n489), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n535), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n637), .A2(KEYINPUT110), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n533), .B2(new_n535), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n714), .B1(new_n622), .B2(new_n715), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n718), .A2(new_n723), .A3(new_n549), .A4(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n713), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n609), .A2(new_n432), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n608), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NOR3_X1   g544(.A1(new_n717), .A2(new_n643), .A3(new_n724), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n686), .A2(new_n731), .ZN(new_n732));
  AOI211_X1 g546(.A(KEYINPUT107), .B(new_n713), .C1(new_n606), .C2(new_n607), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n707), .B1(new_n608), .B2(new_n695), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(new_n550), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n598), .A2(new_n599), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n686), .A2(new_n305), .A3(new_n738), .A4(new_n696), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT42), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n305), .A2(new_n738), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT111), .A3(new_n696), .A4(new_n686), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n723), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n538), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n742), .A2(KEYINPUT42), .A3(new_n686), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT112), .B(G131), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G33));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n658), .B(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n305), .A2(new_n738), .A3(new_n696), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(new_n618), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n609), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n624), .A2(new_n642), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT44), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT116), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n303), .A2(KEYINPUT45), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n192), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n303), .A2(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n300), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT114), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT46), .B1(new_n766), .B2(new_n767), .ZN(new_n770));
  INV_X1    g584(.A(new_n299), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n191), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n661), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n759), .A2(KEYINPUT44), .A3(new_n760), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n738), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(KEYINPUT115), .A3(new_n738), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n762), .A2(new_n775), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  NOR3_X1   g597(.A1(new_n779), .A2(new_n506), .A3(new_n536), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n686), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT117), .B(G140), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G42));
  NAND2_X1  g603(.A1(new_n694), .A2(new_n299), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT49), .Z(new_n791));
  INV_X1    g605(.A(new_n670), .ZN(new_n792));
  INV_X1    g606(.A(new_n679), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n757), .A2(new_n745), .A3(new_n737), .A4(new_n191), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n791), .A2(new_n792), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT118), .Z(new_n796));
  XNOR2_X1  g610(.A(new_n757), .B(KEYINPUT43), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n543), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n779), .A2(new_n713), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n746), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT48), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n717), .A2(new_n724), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n544), .A2(new_n759), .A3(new_n723), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n709), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n195), .A2(G952), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n536), .A2(new_n792), .A3(new_n544), .A4(new_n799), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n805), .B1(new_n806), .B2(new_n619), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n801), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n798), .A2(new_n723), .A3(new_n802), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n679), .A2(new_n550), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n695), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n803), .A2(KEYINPUT50), .A3(new_n695), .A4(new_n811), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n798), .A2(new_n799), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n671), .A2(new_n756), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n816), .A2(new_n731), .B1(new_n806), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n815), .A2(KEYINPUT51), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n810), .A2(new_n779), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n769), .A2(new_n772), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n191), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n790), .A2(new_n621), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n808), .B1(new_n819), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n815), .A2(new_n818), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT121), .B1(new_n785), .B2(new_n786), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n823), .A2(new_n831), .A3(new_n824), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n830), .B(new_n832), .C1(new_n621), .C2(new_n790), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n829), .B1(new_n833), .B2(new_n820), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n828), .B1(new_n834), .B2(KEYINPUT51), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n836));
  INV_X1    g650(.A(new_n659), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n657), .B(KEYINPUT119), .Z(new_n838));
  NAND3_X1  g652(.A1(new_n637), .A2(new_n641), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n493), .B2(new_n668), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n305), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n608), .A2(new_n841), .A3(new_n728), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n687), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n735), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n735), .A2(new_n837), .A3(new_n843), .A4(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n630), .B1(new_n609), .B2(new_n618), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n626), .A2(new_n601), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n729), .A2(new_n602), .A3(new_n645), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n697), .B1(new_n692), .B2(new_n702), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n671), .A2(new_n431), .A3(new_n685), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n854), .A2(new_n649), .B1(new_n686), .B2(new_n731), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n305), .A2(new_n738), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n855), .A2(new_n856), .B1(new_n752), .B2(new_n753), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n744), .B2(new_n747), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n853), .A2(new_n858), .A3(new_n711), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n848), .B2(new_n859), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n659), .B1(new_n709), .B2(new_n732), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(new_n864), .B2(new_n843), .ZN(new_n865));
  INV_X1    g679(.A(new_n847), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n859), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n859), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT54), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n836), .B1(new_n863), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n862), .B1(new_n860), .B2(new_n861), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n869), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(KEYINPUT120), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n835), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n796), .B1(new_n876), .B2(new_n877), .ZN(G75));
  AOI21_X1  g692(.A(new_n190), .B1(new_n869), .B2(new_n870), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(G210), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n589), .A2(new_n595), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n590), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(KEYINPUT123), .A2(KEYINPUT56), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n880), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n884), .B1(new_n880), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n195), .A2(G952), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G51));
  INV_X1    g703(.A(new_n766), .ZN(new_n890));
  OAI211_X1 g704(.A(G902), .B(new_n890), .C1(new_n860), .C2(new_n861), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT124), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n300), .B(KEYINPUT57), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n873), .A2(new_n874), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n298), .B2(new_n293), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n888), .B1(new_n892), .B2(new_n895), .ZN(G54));
  INV_X1    g710(.A(new_n888), .ZN(new_n897));
  AND2_X1   g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n879), .A2(new_n369), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n899), .B2(KEYINPUT125), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n879), .A2(new_n898), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(new_n369), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n900), .B1(new_n903), .B2(new_n899), .ZN(G60));
  AND2_X1   g718(.A1(new_n613), .A2(new_n614), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n616), .B(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n873), .A2(new_n874), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n897), .ZN(new_n909));
  INV_X1    g723(.A(new_n906), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n872), .A2(new_n875), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n909), .B1(new_n911), .B2(new_n905), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT60), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n639), .B(new_n915), .C1(new_n860), .C2(new_n861), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n869), .B2(new_n870), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n916), .B(new_n897), .C1(new_n917), .C2(new_n529), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT61), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n918), .B(new_n920), .ZN(G66));
  NAND2_X1  g735(.A1(G224), .A2(G953), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n547), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n853), .A2(new_n711), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n195), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n881), .B1(G898), .B2(new_n195), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  AOI21_X1  g741(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n355), .A2(new_n359), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n476), .B(new_n929), .Z(new_n930));
  AND2_X1   g744(.A1(new_n864), .A2(new_n687), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n683), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n742), .A2(new_n541), .A3(new_n661), .A4(new_n849), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n782), .A2(new_n787), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n683), .A2(new_n937), .A3(new_n931), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n933), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n930), .B1(new_n939), .B2(new_n195), .ZN(new_n940));
  NAND2_X1  g754(.A1(G900), .A2(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n930), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n782), .A2(new_n787), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n608), .A2(new_n728), .A3(new_n746), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n754), .B1(new_n774), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n744), .B2(new_n747), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n943), .A2(new_n931), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n942), .B1(new_n947), .B2(new_n195), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n928), .B1(new_n940), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n928), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n943), .A2(new_n931), .A3(new_n946), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n930), .B(new_n941), .C1(new_n951), .C2(G953), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n935), .B1(KEYINPUT62), .B2(new_n932), .ZN(new_n953));
  AOI21_X1  g767(.A(G953), .B1(new_n953), .B2(new_n938), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n950), .B(new_n952), .C1(new_n954), .C2(new_n930), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n949), .A2(new_n955), .ZN(G72));
  NAND4_X1  g770(.A1(new_n933), .A2(new_n936), .A3(new_n924), .A4(new_n938), .ZN(new_n957));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  AOI21_X1  g773(.A(new_n665), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n664), .A2(new_n472), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n943), .A2(new_n924), .A3(new_n931), .A4(new_n946), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n959), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n665), .A3(new_n959), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n869), .B2(new_n870), .ZN(new_n967));
  NOR4_X1   g781(.A1(new_n960), .A2(new_n964), .A3(new_n888), .A4(new_n967), .ZN(G57));
endmodule


