//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n207), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n207), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT0), .Z(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  AOI211_X1 g0023(.A(new_n215), .B(new_n218), .C1(new_n221), .C2(new_n223), .ZN(G361));
  XOR2_X1   g0024(.A(G250), .B(G257), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G264), .B(G270), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n228), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G58), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G351));
  AND2_X1   g0043(.A1(KEYINPUT3), .A2(G33), .ZN(new_n244));
  NOR2_X1   g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  OAI211_X1 g0045(.A(G244), .B(G1698), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  OAI211_X1 g0047(.A(G238), .B(new_n247), .C1(new_n244), .C2(new_n245), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G116), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n252), .A2(G274), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G45), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n252), .A2(G250), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G169), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G97), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT19), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n220), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G97), .A2(G107), .ZN(new_n269));
  INV_X1    g0069(.A(G87), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n220), .B(G68), .C1(new_n244), .C2(new_n245), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n220), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G97), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n267), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n272), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n219), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT83), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT15), .B(G87), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n220), .A3(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G1), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n284), .A2(new_n279), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n282), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n280), .A2(new_n281), .A3(new_n285), .A4(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n261), .B1(new_n253), .B2(new_n250), .ZN(new_n292));
  INV_X1    g0092(.A(G179), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n265), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n280), .A2(new_n285), .A3(new_n290), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT83), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n263), .A2(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n288), .A2(G87), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n280), .A2(new_n285), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(G190), .B2(new_n292), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n295), .A2(new_n297), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G283), .ZN(new_n303));
  OAI211_X1 g0103(.A(G250), .B(G1698), .C1(new_n244), .C2(new_n245), .ZN(new_n304));
  OAI211_X1 g0104(.A(G244), .B(new_n247), .C1(new_n244), .C2(new_n245), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT4), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n286), .ZN(new_n309));
  NAND2_X1  g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  AOI21_X1  g0110(.A(G1698), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT4), .B1(new_n311), .B2(G244), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n253), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(KEYINPUT5), .A2(G41), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT5), .A2(G41), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n256), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(G257), .A3(new_n252), .ZN(new_n318));
  AND2_X1   g0118(.A1(G33), .A2(G41), .ZN(new_n319));
  OAI21_X1  g0119(.A(G274), .B1(new_n319), .B2(new_n219), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT81), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(KEYINPUT5), .A2(G41), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n259), .B1(new_n323), .B2(new_n314), .ZN(new_n324));
  INV_X1    g0124(.A(G274), .ZN(new_n325));
  AND2_X1   g0125(.A1(G1), .A2(G13), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n251), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT81), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n318), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT82), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n321), .B1(new_n317), .B2(new_n320), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n324), .A2(KEYINPUT81), .A3(new_n327), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT82), .B1(new_n334), .B2(new_n318), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n293), .B(new_n313), .C1(new_n331), .C2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n244), .A2(new_n245), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n337), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n220), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT77), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT77), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT7), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n220), .B2(new_n337), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n309), .A2(KEYINPUT7), .A3(new_n220), .A4(new_n310), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT78), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(G107), .B(new_n338), .C1(new_n344), .C2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT6), .ZN(new_n349));
  INV_X1    g0149(.A(G107), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n275), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n351), .B2(new_n269), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(KEYINPUT6), .A3(G97), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT70), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(new_n220), .A3(new_n286), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n354), .A2(G20), .B1(G77), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n279), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n283), .A2(G1), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G20), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G97), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n288), .B2(G97), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT5), .B(G41), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n256), .B1(new_n326), .B2(new_n251), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n332), .A2(new_n333), .B1(new_n368), .B2(G257), .ZN(new_n369));
  AOI21_X1  g0169(.A(G169), .B1(new_n313), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n336), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n365), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n360), .B2(new_n279), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n313), .A2(new_n369), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G190), .ZN(new_n376));
  INV_X1    g0176(.A(new_n313), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n329), .A2(new_n330), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n369), .A2(KEYINPUT82), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n374), .B(new_n376), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n302), .A2(new_n372), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT21), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n279), .B1(new_n220), .B2(G116), .ZN(new_n385));
  AOI21_X1  g0185(.A(G20), .B1(G33), .B2(G283), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n286), .A2(G97), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT85), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT85), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n389), .A2(KEYINPUT86), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n387), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT85), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G116), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n278), .A2(new_n219), .B1(G20), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n390), .A2(KEYINPUT86), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n390), .A2(KEYINPUT86), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n284), .A2(new_n396), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n288), .B2(G116), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n392), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G169), .ZN(new_n406));
  OAI211_X1 g0206(.A(G264), .B(G1698), .C1(new_n244), .C2(new_n245), .ZN(new_n407));
  OAI211_X1 g0207(.A(G257), .B(new_n247), .C1(new_n244), .C2(new_n245), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n309), .A2(G303), .A3(new_n310), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT84), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT84), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n407), .A2(new_n408), .A3(new_n412), .A4(new_n409), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n252), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n368), .A2(G270), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n334), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n384), .B1(new_n406), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n411), .A2(new_n413), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n253), .ZN(new_n420));
  INV_X1    g0220(.A(new_n416), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(G190), .ZN(new_n422));
  OAI21_X1  g0222(.A(G200), .B1(new_n414), .B2(new_n416), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n278), .A2(new_n219), .ZN(new_n424));
  INV_X1    g0224(.A(new_n287), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n363), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n402), .B1(new_n426), .B2(new_n396), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n398), .A2(new_n399), .ZN(new_n428));
  INV_X1    g0228(.A(new_n400), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n422), .A2(new_n423), .A3(new_n401), .A4(new_n430), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n414), .A2(new_n416), .A3(new_n293), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n405), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n420), .A2(new_n421), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n434), .A2(KEYINPUT21), .A3(G169), .A4(new_n405), .ZN(new_n435));
  AND4_X1   g0235(.A1(new_n418), .A2(new_n431), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n383), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(G232), .B(G1698), .C1(new_n244), .C2(new_n245), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT71), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n309), .A2(new_n310), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT71), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(G232), .A4(G1698), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(G226), .A3(new_n247), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n439), .A2(new_n442), .A3(new_n266), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n253), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT69), .ZN(new_n446));
  NOR2_X1   g0246(.A1(G41), .A2(G45), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n447), .B2(G1), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n258), .B(KEYINPUT69), .C1(G41), .C2(G45), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(G238), .A3(new_n252), .A4(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n447), .A2(G1), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n327), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n445), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT13), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT13), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n445), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT72), .A3(G200), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n457), .B1(new_n445), .B2(new_n454), .ZN(new_n461));
  AOI211_X1 g0261(.A(KEYINPUT13), .B(new_n453), .C1(new_n444), .C2(new_n253), .ZN(new_n462));
  OAI21_X1  g0262(.A(G200), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT72), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n461), .A2(new_n462), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n202), .B1(new_n356), .B2(new_n357), .ZN(new_n468));
  INV_X1    g0268(.A(G77), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n274), .A2(new_n469), .B1(new_n220), .B2(G68), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n279), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT11), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT12), .B1(new_n363), .B2(G68), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT12), .ZN(new_n475));
  INV_X1    g0275(.A(G68), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n284), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n284), .A2(new_n279), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n220), .A2(G1), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n476), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n474), .A2(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(KEYINPUT11), .B(new_n279), .C1(new_n468), .C2(new_n470), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT73), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n473), .A2(new_n481), .A3(KEYINPUT73), .A4(new_n482), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n467), .A2(G190), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n466), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT74), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n485), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n485), .B2(new_n486), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT14), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n459), .B2(G169), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(G169), .C1(new_n461), .C2(new_n462), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n456), .A2(G179), .A3(new_n458), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT75), .ZN(new_n500));
  XNOR2_X1  g0300(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n424), .A2(new_n363), .ZN(new_n502));
  OAI21_X1  g0302(.A(G50), .B1(new_n220), .B2(G1), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(G50), .B2(new_n363), .ZN(new_n504));
  XNOR2_X1  g0304(.A(KEYINPUT8), .B(G58), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n274), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n506), .A2(new_n507), .B1(G20), .B2(new_n203), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n358), .A2(G150), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n504), .B1(new_n510), .B2(new_n279), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT9), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n311), .A2(G222), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n440), .A2(G223), .A3(G1698), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n514), .B(new_n515), .C1(new_n469), .C2(new_n440), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n253), .ZN(new_n517));
  INV_X1    g0317(.A(new_n452), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n448), .A2(new_n252), .A3(new_n449), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(G226), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(G200), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n513), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT10), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT10), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n513), .A2(new_n523), .A3(new_n527), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(new_n264), .ZN(new_n530));
  INV_X1    g0330(.A(new_n511), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(G179), .C2(new_n521), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n311), .A2(G232), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n440), .A2(G238), .A3(G1698), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n350), .C2(new_n440), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n253), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n518), .B1(new_n519), .B2(G244), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n264), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n506), .A2(new_n358), .ZN(new_n540));
  OAI221_X1 g0340(.A(new_n540), .B1(new_n220), .B2(new_n469), .C1(new_n274), .C2(new_n282), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n279), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n479), .A2(new_n469), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n478), .A2(new_n543), .B1(new_n469), .B2(new_n284), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n539), .B(new_n545), .C1(G179), .C2(new_n538), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n538), .A2(G200), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n536), .A2(G190), .A3(new_n537), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n547), .A2(new_n542), .A3(new_n544), .A4(new_n548), .ZN(new_n549));
  AND4_X1   g0349(.A1(new_n529), .A2(new_n532), .A3(new_n546), .A4(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n505), .A2(new_n479), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n502), .B1(KEYINPUT79), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g0352(.A1(new_n551), .A2(KEYINPUT79), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n553), .B1(new_n284), .B2(new_n505), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n358), .A2(G159), .ZN(new_n556));
  INV_X1    g0356(.A(G58), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n476), .ZN(new_n558));
  OAI21_X1  g0358(.A(G20), .B1(new_n558), .B2(new_n201), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT7), .B1(new_n337), .B2(new_n220), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT76), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n476), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n343), .A2(new_n337), .A3(new_n220), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n309), .A2(new_n220), .A3(new_n310), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n339), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT76), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n560), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n424), .B1(new_n568), .B2(KEYINPUT16), .ZN(new_n569));
  OAI211_X1 g0369(.A(G68), .B(new_n338), .C1(new_n344), .C2(new_n347), .ZN(new_n570));
  INV_X1    g0370(.A(new_n560), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT16), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n555), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n448), .A2(G232), .A3(new_n252), .A4(new_n449), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G223), .A2(G1698), .ZN(new_n576));
  INV_X1    g0376(.A(G226), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(G1698), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n440), .B1(G33), .B2(G87), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n452), .B(new_n575), .C1(new_n579), .C2(new_n252), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n293), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(G169), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT18), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT76), .ZN(new_n584));
  OAI21_X1  g0384(.A(G68), .B1(new_n566), .B2(KEYINPUT76), .ZN(new_n585));
  OAI211_X1 g0385(.A(KEYINPUT16), .B(new_n571), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n279), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n554), .B1(new_n587), .B2(new_n572), .ZN(new_n588));
  INV_X1    g0388(.A(new_n582), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT18), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n580), .A2(new_n381), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G190), .B2(new_n580), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n594), .B(new_n554), .C1(new_n587), .C2(new_n572), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT17), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n574), .A2(KEYINPUT17), .A3(new_n594), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(KEYINPUT80), .B1(new_n592), .B2(new_n599), .ZN(new_n600));
  OR3_X1    g0400(.A1(new_n592), .A2(new_n599), .A3(KEYINPUT80), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n550), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n501), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT24), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n220), .B(G87), .C1(new_n244), .C2(new_n245), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT22), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT22), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n440), .A2(new_n608), .A3(new_n220), .A4(G87), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n350), .A2(KEYINPUT23), .A3(G20), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT23), .B1(new_n350), .B2(G20), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n611), .A2(new_n612), .B1(G20), .B2(new_n249), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n605), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n607), .B2(new_n609), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT24), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n279), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT87), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(KEYINPUT25), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n220), .A2(G107), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(KEYINPUT25), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n619), .A2(new_n362), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n362), .A2(new_n620), .ZN(new_n623));
  OAI221_X1 g0423(.A(new_n622), .B1(new_n621), .B2(new_n623), .C1(new_n426), .C2(new_n350), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(G257), .B(G1698), .C1(new_n244), .C2(new_n245), .ZN(new_n626));
  OAI211_X1 g0426(.A(G250), .B(new_n247), .C1(new_n244), .C2(new_n245), .ZN(new_n627));
  NAND2_X1  g0427(.A1(G33), .A2(G294), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n253), .B1(new_n368), .B2(G264), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n334), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(G190), .ZN(new_n632));
  AOI21_X1  g0432(.A(G200), .B1(new_n630), .B2(new_n334), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n617), .B(new_n625), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n279), .B1(new_n615), .B2(KEYINPUT24), .ZN(new_n635));
  AOI211_X1 g0435(.A(new_n605), .B(new_n613), .C1(new_n607), .C2(new_n609), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n625), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n630), .A2(new_n293), .A3(new_n334), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n631), .A2(new_n264), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT88), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n634), .B2(new_n640), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n437), .B(new_n604), .C1(new_n642), .C2(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n546), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT14), .B1(new_n467), .B2(new_n264), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n496), .A3(new_n495), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n488), .A2(new_n646), .B1(new_n492), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n599), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n529), .B1(new_n650), .B2(new_n592), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(new_n532), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n263), .A2(new_n653), .A3(new_n264), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT89), .B1(new_n292), .B2(G169), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n296), .A4(new_n294), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n263), .A2(KEYINPUT90), .A3(G200), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n292), .B2(new_n381), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n292), .A2(G190), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n280), .A2(new_n285), .A3(new_n299), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n657), .A2(new_n659), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(new_n634), .A3(new_n372), .A4(new_n382), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n640), .A2(new_n435), .A3(new_n418), .A4(new_n433), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n656), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n656), .A2(new_n662), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n372), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT91), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT91), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n671), .B(new_n667), .C1(new_n372), .C2(new_n668), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n336), .A2(new_n366), .A3(new_n371), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(KEYINPUT26), .A3(new_n302), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n666), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n652), .B1(new_n604), .B2(new_n676), .ZN(G369));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n435), .A2(new_n433), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n418), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n362), .A2(new_n220), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT92), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n405), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT93), .B1(new_n680), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n679), .A2(new_n418), .A3(new_n431), .A4(new_n688), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n435), .A2(new_n433), .ZN(new_n692));
  INV_X1    g0492(.A(new_n418), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n689), .B(KEYINPUT93), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT94), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT93), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n688), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT94), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n691), .A4(new_n694), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n678), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n644), .A2(new_n642), .ZN(new_n703));
  INV_X1    g0503(.A(new_n637), .ZN(new_n704));
  INV_X1    g0504(.A(new_n687), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n640), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n687), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n705), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n644), .A2(new_n642), .B1(new_n637), .B2(new_n687), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n698), .A2(new_n687), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n711), .A3(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n216), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n271), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n720), .B(KEYINPUT95), .C1(new_n222), .C2(new_n718), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(KEYINPUT95), .B2(new_n720), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  INV_X1    g0523(.A(KEYINPUT96), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n292), .A2(new_n630), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n334), .A2(G179), .A3(new_n415), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n420), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n375), .A2(KEYINPUT30), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n313), .A2(new_n369), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n313), .B1(new_n331), .B2(new_n335), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n631), .A2(new_n293), .A3(new_n263), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n434), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n731), .A2(new_n730), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n432), .A2(new_n736), .A3(KEYINPUT96), .A4(new_n725), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n729), .A2(new_n732), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n739));
  AOI21_X1  g0539(.A(KEYINPUT31), .B1(new_n738), .B2(new_n687), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n703), .A2(new_n383), .A3(new_n436), .A4(new_n705), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n678), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT97), .ZN(new_n745));
  INV_X1    g0545(.A(new_n656), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n372), .A2(new_n382), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n634), .A2(new_n656), .A3(new_n662), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n418), .A2(new_n435), .A3(new_n640), .A4(new_n433), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n670), .A2(new_n674), .A3(new_n672), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n745), .B(new_n687), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n372), .A2(new_n382), .ZN(new_n754));
  INV_X1    g0554(.A(new_n748), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n754), .A2(new_n755), .A3(new_n750), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n672), .A2(new_n674), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n370), .B1(new_n380), .B2(new_n293), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(new_n366), .A3(new_n656), .A4(new_n662), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n671), .B1(new_n759), .B2(new_n667), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n656), .B(new_n756), .C1(new_n757), .C2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT97), .B1(new_n761), .B2(new_n705), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n744), .B1(new_n753), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT26), .B1(new_n673), .B2(new_n302), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n372), .A2(new_n668), .A3(new_n667), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n705), .B1(new_n666), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n744), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n743), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n723), .B1(new_n770), .B2(G1), .ZN(G364));
  NOR2_X1   g0571(.A1(new_n283), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n258), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n717), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n702), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n696), .A2(new_n678), .A3(new_n701), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n696), .A2(new_n701), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n220), .A2(new_n293), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(G317), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(KEYINPUT33), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G190), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G179), .A2(G200), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n220), .B1(new_n792), .B2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n791), .A2(G326), .B1(G294), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT102), .Z(new_n796));
  NOR2_X1   g0596(.A1(new_n220), .A2(new_n790), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(G179), .A3(new_n381), .ZN(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n783), .A2(new_n790), .A3(new_n381), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n381), .A2(G179), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n440), .B(new_n802), .C1(G303), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT101), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n220), .B2(G190), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n790), .A2(KEYINPUT101), .A3(G20), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n808), .A2(new_n809), .A3(new_n792), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G283), .A2(new_n811), .B1(new_n813), .B2(G329), .ZN(new_n814));
  AND4_X1   g0614(.A1(new_n789), .A2(new_n796), .A3(new_n806), .A4(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT103), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(KEYINPUT103), .ZN(new_n817));
  INV_X1    g0617(.A(new_n798), .ZN(new_n818));
  INV_X1    g0618(.A(new_n800), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(G58), .B1(new_n819), .B2(G77), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT100), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n820), .A2(new_n821), .B1(new_n350), .B2(new_n810), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G50), .A2(new_n791), .B1(new_n785), .B2(G68), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n794), .A2(G97), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n337), .B1(new_n805), .B2(G87), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n813), .A2(G159), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(KEYINPUT32), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n823), .B(new_n829), .C1(KEYINPUT32), .C2(new_n828), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n816), .A2(new_n817), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n219), .B1(G20), .B2(new_n264), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT99), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT99), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n781), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n716), .A2(new_n440), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n242), .A2(G45), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT98), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(new_n255), .C2(new_n223), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n216), .A2(G355), .A3(new_n440), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(G116), .B2(new_n216), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n837), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n782), .A2(new_n836), .A3(new_n775), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n778), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G396));
  NAND2_X1  g0648(.A1(new_n687), .A2(new_n545), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n549), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n546), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n646), .A2(new_n705), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n753), .B2(new_n762), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n546), .A2(new_n705), .A3(new_n549), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n751), .B2(new_n752), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n743), .ZN(new_n859));
  INV_X1    g0659(.A(new_n775), .ZN(new_n860));
  INV_X1    g0660(.A(new_n743), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n854), .A2(new_n861), .A3(new_n857), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT106), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n818), .A2(G294), .B1(new_n805), .B2(G107), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n811), .A2(G87), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n440), .B1(new_n819), .B2(G116), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n785), .ZN(new_n869));
  INV_X1    g0669(.A(G283), .ZN(new_n870));
  INV_X1    g0670(.A(G303), .ZN(new_n871));
  INV_X1    g0671(.A(new_n791), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n825), .B1(new_n869), .B2(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n868), .B(new_n873), .C1(G311), .C2(new_n813), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n440), .B1(new_n793), .B2(new_n557), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n811), .A2(G68), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n202), .B2(new_n804), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT105), .Z(new_n878));
  AOI211_X1 g0678(.A(new_n875), .B(new_n878), .C1(G132), .C2(new_n813), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n818), .A2(G143), .B1(new_n819), .B2(G159), .ZN(new_n880));
  AOI22_X1  g0680(.A1(G137), .A2(new_n791), .B1(new_n785), .B2(G150), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT34), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n874), .B1(new_n879), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n835), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n835), .A2(new_n779), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n887), .A2(new_n888), .B1(G77), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n853), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n780), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n775), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n863), .A2(new_n864), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n864), .B1(new_n863), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(G384));
  OR2_X1    g0697(.A1(new_n354), .A2(KEYINPUT35), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n354), .A2(KEYINPUT35), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n898), .A2(G116), .A3(new_n221), .A4(new_n899), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT36), .Z(new_n901));
  OR3_X1    g0701(.A1(new_n558), .A2(new_n222), .A3(new_n469), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n202), .A2(G68), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n258), .B(G13), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n571), .B1(new_n584), .B2(new_n585), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT16), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n555), .B1(new_n569), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n685), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n592), .B2(new_n599), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n595), .B1(new_n910), .B2(new_n685), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n582), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n588), .A2(new_n589), .ZN(new_n916));
  INV_X1    g0716(.A(new_n685), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n588), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT37), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n595), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n912), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT108), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n498), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n648), .A2(KEYINPUT108), .A3(new_n492), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n466), .A2(new_n487), .B1(new_n492), .B2(new_n687), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n485), .A2(new_n486), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n459), .B2(new_n790), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n465), .B2(new_n460), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n492), .B(new_n687), .C1(new_n934), .C2(new_n648), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n853), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n738), .A2(new_n687), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT31), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n705), .B1(new_n942), .B2(new_n643), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n437), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT110), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT110), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n742), .A2(new_n946), .A3(new_n939), .A4(new_n940), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n926), .A2(new_n936), .A3(new_n945), .A4(new_n947), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n945), .A2(new_n936), .A3(new_n947), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n595), .B1(new_n574), .B2(new_n582), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n574), .A2(new_n685), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT37), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(KEYINPUT109), .A3(new_n920), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n951), .B1(new_n592), .B2(new_n599), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT109), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n955), .B(KEYINPUT37), .C1(new_n950), .C2(new_n951), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n923), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n906), .B1(new_n958), .B2(new_n925), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n906), .A2(new_n948), .B1(new_n949), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n603), .A2(new_n945), .A3(new_n947), .ZN(new_n962));
  OAI21_X1  g0762(.A(G330), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  INV_X1    g0764(.A(new_n852), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT107), .B1(new_n856), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT107), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n967), .B(new_n852), .C1(new_n676), .C2(new_n855), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n931), .A2(new_n935), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n926), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n687), .B1(new_n928), .B2(new_n929), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n923), .B2(new_n957), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n972), .B(new_n973), .C1(new_n975), .C2(KEYINPUT39), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n592), .A2(new_n685), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n971), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n763), .A2(new_n603), .A3(new_n769), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n652), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n978), .B(new_n980), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n964), .A2(new_n981), .B1(new_n258), .B2(new_n772), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n964), .A2(new_n981), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n905), .B1(new_n982), .B2(new_n983), .ZN(G367));
  NAND2_X1  g0784(.A1(new_n707), .A2(new_n382), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n687), .B1(new_n985), .B2(new_n372), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n705), .A2(new_n374), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n747), .A2(new_n987), .B1(new_n372), .B2(new_n705), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n712), .A2(new_n713), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n986), .B1(new_n989), .B2(KEYINPUT42), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT111), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n687), .A2(new_n300), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n663), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n656), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n989), .A2(KEYINPUT42), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n990), .B2(KEYINPUT111), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n991), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT112), .ZN(new_n999));
  INV_X1    g0799(.A(new_n710), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n988), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n991), .A2(new_n997), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n994), .B(KEYINPUT43), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n999), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1002), .B1(new_n999), .B2(new_n1005), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n717), .B(KEYINPUT41), .Z(new_n1009));
  INV_X1    g0809(.A(new_n713), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n706), .A2(new_n708), .A3(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(new_n714), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n702), .B2(KEYINPUT113), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n702), .A2(KEYINPUT113), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n770), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT114), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n988), .B1(new_n714), .B2(new_n711), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT44), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n714), .A2(new_n988), .A3(new_n711), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(new_n710), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT113), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1025), .B(new_n678), .C1(new_n696), .C2(new_n701), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1013), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT114), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n770), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1017), .A2(new_n1024), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1009), .B1(new_n1030), .B2(new_n770), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1008), .B1(new_n1031), .B2(new_n774), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n440), .B1(new_n804), .B2(new_n557), .ZN(new_n1033));
  INV_X1    g0833(.A(G159), .ZN(new_n1034));
  INV_X1    g0834(.A(G143), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n869), .A2(new_n1034), .B1(new_n872), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1033), .B(new_n1036), .C1(G50), .C2(new_n819), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n794), .A2(G68), .ZN(new_n1038));
  INV_X1    g0838(.A(G150), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1038), .B1(new_n1039), .B2(new_n798), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n813), .A2(G137), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n811), .A2(G77), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1037), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n337), .B1(new_n800), .B2(new_n870), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G294), .B2(new_n785), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n275), .B2(new_n810), .C1(new_n786), .C2(new_n812), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G311), .A2(new_n791), .B1(new_n818), .B2(G303), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT115), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT46), .B1(new_n805), .B2(G116), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G107), .B2(new_n794), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1048), .A2(KEYINPUT115), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1044), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT117), .Z(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT47), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(KEYINPUT47), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n835), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n228), .A2(new_n838), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n781), .B(new_n835), .C1(new_n716), .C2(new_n289), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n860), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n781), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1059), .B(new_n1062), .C1(new_n1063), .C2(new_n994), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1032), .A2(new_n1064), .ZN(G387));
  NAND2_X1  g0865(.A1(new_n1027), .A2(new_n770), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n717), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n706), .A2(new_n708), .A3(new_n781), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n233), .A2(G45), .A3(new_n337), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT50), .B1(new_n505), .B2(G50), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n255), .C1(new_n476), .C2(new_n469), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n505), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n337), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n719), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n716), .B1(new_n1070), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n837), .B1(new_n350), .B2(new_n216), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n775), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n440), .B1(new_n813), .B2(G326), .ZN(new_n1079));
  INV_X1    g0879(.A(G294), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n804), .A2(new_n1080), .B1(new_n793), .B2(new_n870), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n818), .A2(G317), .B1(new_n819), .B2(G303), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n801), .B2(new_n869), .C1(new_n799), .C2(new_n872), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT48), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1084), .B2(new_n1083), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT49), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1079), .B1(new_n396), .B2(new_n810), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n794), .A2(new_n289), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n869), .B2(new_n505), .C1(new_n1034), .C2(new_n872), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n440), .B1(new_n800), .B2(new_n476), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n798), .A2(new_n202), .B1(new_n804), .B2(new_n469), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G97), .C2(new_n811), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT118), .B(G150), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n812), .B2(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1088), .A2(new_n1089), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1078), .B1(new_n1097), .B2(new_n835), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1027), .A2(new_n774), .B1(new_n1069), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1068), .A2(new_n1099), .ZN(G393));
  AND2_X1   g0900(.A1(new_n238), .A2(new_n838), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n837), .B1(new_n275), .B2(new_n216), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n775), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n872), .A2(new_n1039), .B1(new_n1034), .B2(new_n798), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT51), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n793), .A2(new_n469), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n440), .B1(new_n800), .B2(new_n505), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G50), .C2(new_n785), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1105), .A2(new_n866), .A3(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n812), .A2(new_n1035), .B1(new_n804), .B2(new_n476), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT119), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G317), .A2(new_n791), .B1(new_n818), .B2(G311), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT52), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n869), .A2(new_n871), .B1(new_n793), .B2(new_n396), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n337), .B1(new_n804), .B2(new_n870), .C1(new_n1080), .C2(new_n800), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n350), .A2(new_n810), .B1(new_n812), .B2(new_n799), .ZN(new_n1116));
  OR3_X1    g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1109), .A2(new_n1111), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1103), .B1(new_n1118), .B2(new_n835), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n988), .B2(new_n1063), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1023), .B(new_n1000), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n773), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n718), .B1(new_n1121), .B2(new_n1066), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1030), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(G390));
  NAND4_X1  g0925(.A1(new_n603), .A2(G330), .A3(new_n945), .A4(new_n947), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n979), .A2(new_n652), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n705), .B(new_n851), .C1(new_n666), .C2(new_n766), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n852), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT120), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT120), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1129), .A2(new_n1132), .A3(new_n852), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n678), .B(new_n853), .C1(new_n741), .C2(new_n742), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1131), .A2(new_n1133), .B1(new_n1134), .B2(new_n970), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n970), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n945), .A2(G330), .A3(new_n947), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n853), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n945), .A2(new_n936), .A3(G330), .A4(new_n947), .ZN(new_n1140));
  OAI211_X1 g0940(.A(G330), .B(new_n892), .C1(new_n941), .C2(new_n944), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1136), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n969), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1128), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n973), .B1(new_n975), .B2(KEYINPUT39), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1136), .B1(new_n966), .B2(new_n968), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n972), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1131), .A2(new_n970), .A3(new_n1133), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n975), .A2(new_n972), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1134), .A2(new_n970), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1149), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1140), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1146), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1140), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1135), .A2(new_n1138), .B1(new_n1143), .B2(new_n969), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(new_n1127), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1149), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1156), .A2(new_n1163), .A3(new_n717), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1147), .A2(new_n779), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n775), .B1(new_n506), .B2(new_n890), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n791), .A2(G128), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1034), .B2(new_n793), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n804), .A2(new_n1095), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(KEYINPUT53), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT54), .B(G143), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n440), .B1(new_n800), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G132), .B2(new_n818), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1170), .A2(KEYINPUT53), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G137), .B2(new_n785), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G50), .A2(new_n811), .B1(new_n813), .B2(G125), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1171), .A2(new_n1174), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n798), .A2(new_n396), .B1(new_n800), .B2(new_n275), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n440), .B(new_n1179), .C1(G87), .C2(new_n805), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n876), .C1(new_n1080), .C2(new_n812), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1106), .B1(new_n785), .B2(G107), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n870), .B2(new_n872), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1178), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1167), .B1(new_n1184), .B2(new_n835), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1165), .A2(new_n774), .B1(new_n1166), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1164), .A2(new_n1186), .ZN(G378));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1127), .B1(new_n1165), .B2(new_n1161), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n949), .A2(new_n959), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n945), .A2(new_n936), .A3(new_n947), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n924), .A2(new_n925), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n906), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1193), .A3(G330), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n529), .A2(new_n532), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n685), .A2(new_n511), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1194), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1190), .A2(new_n1193), .A3(G330), .A4(new_n1204), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1206), .A2(new_n978), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n978), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1188), .B1(new_n1189), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n971), .A2(new_n976), .A3(new_n977), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1204), .B1(new_n960), .B2(G330), .ZN(new_n1213));
  AND4_X1   g1013(.A1(G330), .A2(new_n1190), .A3(new_n1193), .A4(new_n1204), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1206), .A2(new_n978), .A3(new_n1207), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1188), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1163), .A2(new_n1128), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n718), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1211), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1205), .A2(new_n779), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n440), .A2(G41), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1223), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(G107), .B2(new_n818), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n811), .A2(G58), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n819), .A2(new_n289), .B1(new_n805), .B2(G77), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1038), .B1(new_n869), .B2(new_n275), .C1(new_n396), .C2(new_n872), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G283), .C2(new_n813), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1224), .B1(new_n1230), .B2(KEYINPUT58), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT121), .Z(new_n1232));
  NOR2_X1   g1032(.A1(new_n804), .A2(new_n1172), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G128), .B2(new_n818), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n785), .A2(G132), .B1(G150), .B2(new_n794), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n819), .A2(G137), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n791), .A2(G125), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT59), .ZN(new_n1239));
  AOI211_X1 g1039(.A(G33), .B(G41), .C1(new_n813), .C2(G124), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1034), .B2(new_n810), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1238), .B2(KEYINPUT59), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1230), .A2(KEYINPUT58), .B1(new_n1239), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n888), .B1(new_n1232), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT122), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n860), .B(new_n1245), .C1(new_n202), .C2(new_n889), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1221), .A2(new_n774), .B1(new_n1222), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1220), .A2(new_n1247), .ZN(G375));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1145), .A2(new_n1249), .A3(new_n774), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT123), .B1(new_n1160), .B2(new_n773), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n775), .B1(G68), .B2(new_n890), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G294), .A2(new_n791), .B1(new_n819), .B2(G107), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n396), .B2(new_n869), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT124), .Z(new_n1255));
  OAI21_X1  g1055(.A(new_n337), .B1(new_n804), .B2(new_n275), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G283), .B2(new_n818), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n813), .A2(G303), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(new_n1043), .A3(new_n1090), .A4(new_n1258), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n791), .A2(G132), .B1(G50), .B2(new_n794), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n869), .B2(new_n1172), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n819), .A2(G150), .B1(new_n805), .B2(G159), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n337), .B1(new_n818), .B2(G137), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n813), .A2(G128), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1226), .A4(new_n1264), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n1255), .A2(new_n1259), .B1(new_n1261), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1252), .B1(new_n1266), .B2(new_n835), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n970), .B2(new_n780), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1250), .A2(new_n1251), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1009), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1160), .A2(new_n1127), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1146), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(G381));
  NAND2_X1  g1074(.A1(new_n1246), .A2(new_n1222), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1210), .B2(new_n773), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1211), .B2(new_n1219), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1164), .A2(new_n1186), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n895), .A2(new_n896), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1124), .A3(new_n1281), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(G387), .A2(G381), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1279), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1284), .B2(new_n1283), .ZN(G407));
  NAND2_X1  g1086(.A1(new_n686), .A2(G213), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(KEYINPUT126), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1279), .A2(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(KEYINPUT127), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G407), .A3(G213), .ZN(G409));
  NAND3_X1  g1092(.A1(new_n1218), .A2(new_n1271), .A3(new_n1221), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1278), .A2(new_n1247), .A3(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1289), .B(new_n1294), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1160), .A2(new_n1127), .A3(KEYINPUT60), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n717), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT60), .B1(new_n1160), .B2(new_n1127), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1272), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1281), .B1(new_n1299), .B2(new_n1269), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1298), .A2(new_n1272), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1270), .B(G384), .C1(new_n1301), .C2(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(KEYINPUT62), .B1(new_n1295), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1288), .A2(G2897), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1300), .A2(new_n1302), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G375), .A2(G378), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1276), .A2(G378), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1288), .B1(new_n1311), .B2(new_n1293), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1303), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1310), .A2(new_n1312), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1304), .A2(new_n1309), .A3(new_n1315), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1032), .A2(new_n1064), .A3(G390), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G390), .B1(new_n1032), .B2(new_n1064), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n847), .B1(new_n1068), .B2(new_n1099), .ZN(new_n1319));
  OAI22_X1  g1119(.A1(new_n1317), .A2(new_n1318), .B1(new_n1280), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G387), .A2(new_n1124), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1280), .A2(new_n1319), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1032), .A2(new_n1064), .A3(G390), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1320), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1316), .A2(new_n1325), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1320), .A2(new_n1324), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1295), .B2(new_n1303), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1310), .A2(new_n1312), .A3(KEYINPUT63), .A4(new_n1314), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1327), .A2(new_n1329), .A3(new_n1330), .A4(new_n1309), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(G405));
  NAND3_X1  g1132(.A1(new_n1310), .A2(new_n1279), .A3(new_n1303), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1303), .B1(new_n1310), .B2(new_n1279), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1334), .A2(new_n1325), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1310), .A2(new_n1279), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1314), .ZN(new_n1338));
  AOI22_X1  g1138(.A1(new_n1338), .A2(new_n1333), .B1(new_n1324), .B2(new_n1320), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1336), .A2(new_n1339), .ZN(G402));
endmodule


