//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT82), .A2(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT82), .A2(G107), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(G104), .C1(new_n190), .C2(new_n191), .ZN(new_n192));
  OAI211_X1 g006(.A(KEYINPUT81), .B(KEYINPUT3), .C1(new_n187), .C2(G107), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT81), .B1(new_n196), .B2(KEYINPUT3), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n188), .B(new_n192), .C1(new_n194), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT83), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n193), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n204), .A2(KEYINPUT83), .A3(new_n188), .A4(new_n192), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(G101), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n204), .A2(new_n207), .A3(new_n188), .A4(new_n192), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(KEYINPUT4), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G116), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G119), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n213));
  INV_X1    g027(.A(G119), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G116), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(KEYINPUT68), .A3(G119), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT67), .ZN(new_n218));
  XOR2_X1   g032(.A(KEYINPUT2), .B(G113), .Z(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n200), .A2(new_n222), .A3(G101), .A4(new_n205), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n210), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n211), .A2(KEYINPUT5), .A3(G119), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n228), .A2(KEYINPUT87), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(KEYINPUT87), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G113), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n225), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT82), .B(G107), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n196), .B1(new_n233), .B2(G104), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n208), .A2(new_n235), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n224), .A2(new_n239), .A3(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(KEYINPUT6), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g060(.A(G128), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G146), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(KEYINPUT64), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n252), .A3(new_n248), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n249), .B1(new_n253), .B2(KEYINPUT65), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n247), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n248), .B1(new_n250), .B2(new_n252), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(new_n245), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n246), .A3(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G125), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT0), .B(G128), .Z(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n254), .B2(new_n256), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n259), .A2(KEYINPUT0), .A3(G128), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n268), .A2(KEYINPUT88), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(KEYINPUT88), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT89), .B(G224), .Z(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n274), .B(new_n263), .C1(new_n269), .C2(new_n270), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n238), .A2(new_n279), .A3(new_n240), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n243), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G210), .B1(G237), .B2(G902), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(KEYINPUT7), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n263), .B(new_n284), .C1(new_n269), .C2(new_n270), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n242), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n231), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n226), .A2(KEYINPUT90), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT90), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n217), .A2(new_n289), .A3(KEYINPUT5), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n236), .B1(new_n291), .B2(new_n225), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n208), .A2(new_n235), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(new_n232), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n239), .B(KEYINPUT8), .Z(new_n295));
  NOR3_X1   g109(.A1(new_n292), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n283), .B1(new_n262), .B2(new_n268), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT91), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT91), .B(new_n283), .C1(new_n262), .C2(new_n268), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n286), .B2(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n281), .A2(new_n282), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n282), .B(KEYINPUT93), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n281), .A2(new_n302), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT92), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n281), .A2(new_n302), .A3(KEYINPUT92), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n303), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT94), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT94), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n281), .A2(KEYINPUT92), .A3(new_n302), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT92), .B1(new_n281), .B2(new_n302), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n314), .A2(new_n315), .A3(new_n304), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n313), .B(new_n310), .C1(new_n316), .C2(new_n303), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT9), .B(G234), .Z(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G221), .B1(new_n320), .B2(G902), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n266), .A2(new_n267), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n210), .A2(new_n324), .A3(new_n223), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT84), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT84), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n210), .A2(new_n327), .A3(new_n324), .A4(new_n223), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT11), .ZN(new_n330));
  INV_X1    g144(.A(G134), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(G137), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(G137), .ZN(new_n333));
  INV_X1    g147(.A(G137), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT11), .A3(G134), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G131), .ZN(new_n337));
  INV_X1    g151(.A(G131), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n332), .A2(new_n335), .A3(new_n338), .A4(new_n333), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n342));
  INV_X1    g156(.A(G128), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(new_n259), .ZN(new_n345));
  NOR4_X1   g159(.A1(new_n258), .A2(KEYINPUT1), .A3(new_n343), .A4(new_n245), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n347), .A2(new_n236), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n260), .B1(new_n259), .B2(new_n344), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT85), .B1(new_n293), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n342), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT65), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT64), .B(G143), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n354), .B2(new_n248), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n255), .B1(new_n355), .B2(new_n249), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n346), .B1(new_n356), .B2(new_n247), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n357), .A2(new_n342), .A3(new_n236), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n329), .A2(new_n341), .A3(new_n352), .A4(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G110), .B(G140), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n273), .A2(G227), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n361), .B(new_n362), .Z(new_n363));
  AND2_X1   g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n329), .A2(new_n352), .A3(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n340), .ZN(new_n366));
  OAI22_X1  g180(.A1(new_n349), .A2(new_n351), .B1(new_n261), .B2(new_n293), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT12), .A3(new_n340), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT12), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n348), .B1(new_n347), .B2(new_n236), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n293), .A2(new_n350), .A3(KEYINPUT85), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n370), .A2(new_n371), .B1(new_n357), .B2(new_n236), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n369), .B1(new_n372), .B2(new_n341), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n360), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n363), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n364), .A2(new_n366), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G469), .B1(new_n377), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(G902), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT86), .B(G469), .Z(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n363), .B1(new_n366), .B2(new_n360), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n360), .A2(new_n374), .A3(new_n363), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n379), .B(new_n381), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n322), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G478), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT15), .ZN(new_n387));
  INV_X1    g201(.A(G122), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G116), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT98), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(G116), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT98), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(KEYINPUT14), .C1(new_n388), .C2(G116), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT99), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n391), .A2(KEYINPUT99), .A3(new_n392), .A4(new_n394), .ZN(new_n398));
  INV_X1    g212(.A(new_n389), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(new_n398), .C1(KEYINPUT14), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G107), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n399), .A2(new_n392), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n233), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n343), .A2(G143), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n354), .B2(new_n343), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(G134), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n402), .B(new_n233), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n405), .A2(G134), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n354), .A2(KEYINPUT13), .A3(new_n343), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT13), .ZN(new_n411));
  OAI21_X1  g225(.A(G134), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n319), .A2(G217), .A3(new_n273), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n387), .B1(new_n419), .B2(G902), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n418), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(new_n379), .C1(KEYINPUT15), .C2(new_n386), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G237), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n273), .A3(G214), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n426), .A2(G143), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n354), .A2(new_n426), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(new_n338), .ZN(new_n431));
  XNOR2_X1  g245(.A(G125), .B(G140), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(new_n248), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n428), .A3(G131), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n431), .B(new_n433), .C1(new_n430), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(KEYINPUT16), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT16), .ZN(new_n437));
  INV_X1    g251(.A(G140), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(G125), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT75), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT75), .A4(G125), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(G146), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n441), .A3(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n248), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n429), .A2(new_n338), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n434), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n434), .A2(new_n450), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n435), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n187), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(KEYINPUT96), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n435), .B(new_n459), .C1(new_n448), .C2(new_n453), .ZN(new_n460));
  AOI21_X1  g274(.A(G902), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT97), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G475), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n273), .A2(G952), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(G234), .B2(G237), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n379), .B(new_n273), .C1(G234), .C2(G237), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT21), .B(G898), .Z(new_n469));
  OAI21_X1  g283(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT100), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n432), .A2(KEYINPUT95), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT19), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n474), .A2(new_n248), .B1(new_n449), .B2(new_n434), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT77), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n443), .B(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n435), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n457), .ZN(new_n480));
  AOI21_X1  g294(.A(G475), .B1(new_n480), .B2(new_n460), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n379), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT20), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n484), .A3(new_n379), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n424), .A2(new_n463), .A3(new_n471), .A4(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT101), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n318), .A2(new_n385), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT80), .ZN(new_n490));
  NOR2_X1   g304(.A1(G472), .A2(G902), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT31), .ZN(new_n492));
  INV_X1    g306(.A(new_n333), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n331), .A2(G137), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n339), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n261), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n266), .A2(new_n340), .A3(new_n267), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n220), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT66), .B1(new_n261), .B2(new_n497), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n504), .B(new_n496), .C1(new_n257), .C2(new_n260), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n499), .B(KEYINPUT30), .C1(new_n357), .C2(new_n496), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT69), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n498), .A2(KEYINPUT69), .A3(KEYINPUT30), .A4(new_n499), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n502), .A2(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n501), .B1(new_n511), .B2(new_n221), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n425), .A2(new_n273), .A3(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n207), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n514), .B(new_n515), .Z(new_n516));
  AOI21_X1  g330(.A(new_n492), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n506), .A2(new_n502), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n509), .A2(new_n510), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(new_n221), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(new_n492), .A3(new_n500), .A4(new_n516), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n506), .A2(new_n221), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n501), .A2(KEYINPUT28), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n500), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n516), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n491), .B1(new_n517), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT32), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n520), .A2(new_n500), .A3(new_n516), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT31), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n521), .A3(new_n528), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n491), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(KEYINPUT70), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n538), .A3(new_n531), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G472), .ZN(new_n541));
  INV_X1    g355(.A(new_n512), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT29), .B1(new_n542), .B2(new_n527), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n527), .B2(new_n526), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n498), .A2(new_n499), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n221), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n524), .B1(new_n546), .B2(new_n500), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n547), .A2(KEYINPUT71), .ZN(new_n548));
  INV_X1    g362(.A(new_n525), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT71), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n516), .A2(KEYINPUT29), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n541), .B1(new_n544), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n540), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G110), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n343), .A2(G119), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(KEYINPUT23), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n343), .A2(G119), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT23), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n559), .B2(new_n560), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n559), .B1(new_n563), .B2(KEYINPUT73), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(KEYINPUT73), .B2(new_n559), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT24), .B(G110), .ZN(new_n569));
  OAI221_X1 g383(.A(new_n448), .B1(new_n558), .B2(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n558), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n569), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n571), .A2(new_n572), .B1(new_n248), .B2(new_n432), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n477), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT22), .B(G137), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n575), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G234), .ZN(new_n580));
  OAI21_X1  g394(.A(G217), .B1(new_n580), .B2(G902), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT72), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT79), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n379), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT78), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT25), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n579), .A2(new_n587), .A3(new_n588), .A4(new_n379), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n582), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n585), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n490), .B1(new_n557), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n555), .B1(new_n537), .B2(new_n539), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n597), .A2(KEYINPUT80), .A3(new_n594), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n489), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n378), .A2(new_n384), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n535), .A2(new_n379), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n602), .A2(G472), .B1(new_n491), .B2(new_n535), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n601), .A2(new_n603), .A3(new_n321), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n595), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n282), .B1(new_n281), .B2(new_n302), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n310), .B1(new_n303), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n421), .A2(KEYINPUT33), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n421), .A2(KEYINPUT33), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(G478), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(G478), .A2(G902), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n421), .A2(new_n386), .A3(new_n379), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n463), .A2(new_n486), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n471), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n608), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n187), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n623));
  INV_X1    g437(.A(new_n485), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n484), .B1(new_n481), .B2(new_n379), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n483), .A2(KEYINPUT103), .A3(new_n485), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n462), .A2(G475), .B1(new_n420), .B2(new_n422), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n471), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT104), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n608), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n578), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT105), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n575), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n583), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n593), .A2(new_n640), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n318), .A2(new_n604), .A3(new_n488), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT37), .B(G110), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n467), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n466), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n628), .A2(new_n629), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT106), .ZN(new_n649));
  INV_X1    g463(.A(new_n607), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n641), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n557), .A2(new_n649), .A3(new_n385), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XNOR2_X1  g468(.A(new_n647), .B(KEYINPUT39), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n385), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n616), .A2(new_n423), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n512), .A2(new_n527), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n546), .A2(new_n500), .A3(new_n527), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n663));
  AOI21_X1  g477(.A(G902), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n540), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n309), .B(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n668), .A2(new_n641), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n659), .A2(new_n310), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n354), .ZN(G45));
  NAND3_X1  g487(.A1(new_n615), .A2(new_n616), .A3(new_n647), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n557), .A2(new_n652), .A3(new_n385), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  AOI21_X1  g491(.A(new_n594), .B1(new_n540), .B2(new_n556), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g495(.A(KEYINPUT109), .B(new_n379), .C1(new_n382), .C2(new_n383), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(G469), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n321), .A4(new_n384), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(G469), .ZN(new_n686));
  INV_X1    g500(.A(new_n360), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n358), .B1(new_n326), .B2(new_n328), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n341), .B1(new_n688), .B2(new_n352), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n376), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n360), .A2(new_n374), .A3(new_n363), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT109), .B1(new_n692), .B2(new_n379), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n321), .B(new_n384), .C1(new_n686), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT110), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n678), .A2(new_n650), .A3(new_n685), .A4(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n617), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT41), .B(G113), .Z(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT111), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n697), .B(new_n699), .ZN(G15));
  NOR2_X1   g514(.A1(new_n696), .A2(new_n631), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n211), .ZN(G18));
  NOR2_X1   g516(.A1(new_n597), .A2(new_n651), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n488), .A3(new_n685), .A4(new_n695), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND3_X1  g519(.A1(new_n650), .A2(new_n616), .A3(new_n423), .ZN(new_n706));
  INV_X1    g520(.A(new_n471), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n491), .ZN(new_n709));
  INV_X1    g523(.A(new_n521), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n527), .B2(new_n551), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n711), .B2(new_n534), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n541), .B1(new_n535), .B2(new_n379), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n594), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n695), .A2(new_n708), .A3(new_n685), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  NOR3_X1   g530(.A1(new_n674), .A2(new_n712), .A3(new_n713), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n695), .A2(new_n685), .A3(new_n652), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  NAND2_X1  g533(.A1(new_n532), .A2(new_n536), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n595), .B1(new_n720), .B2(new_n555), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n721), .A2(new_n722), .A3(new_n674), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n321), .A2(new_n601), .A3(new_n310), .A4(new_n309), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n678), .A2(new_n675), .A3(new_n724), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(KEYINPUT112), .A3(new_n722), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT112), .B1(new_n726), .B2(new_n722), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  AND2_X1   g545(.A1(new_n678), .A2(new_n724), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n649), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND2_X1  g548(.A1(new_n377), .A2(KEYINPUT45), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n737), .B(G469), .C1(KEYINPUT45), .C2(new_n377), .ZN(new_n738));
  NAND2_X1  g552(.A1(G469), .A2(G902), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT46), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  INV_X1    g555(.A(new_n384), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n322), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n616), .A2(new_n614), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT43), .B1(new_n616), .B2(new_n614), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n641), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n750), .A2(new_n603), .A3(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n744), .A2(new_n655), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n309), .A2(new_n310), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n334), .ZN(G39));
  XNOR2_X1  g574(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n743), .B2(new_n322), .ZN(new_n763));
  INV_X1    g577(.A(new_n741), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n384), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n321), .A3(new_n761), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n557), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n595), .A2(new_n756), .A3(new_n674), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  NAND3_X1  g585(.A1(new_n683), .A2(new_n322), .A3(new_n384), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n763), .A2(new_n767), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n714), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n749), .A2(new_n465), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT120), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n749), .A2(new_n777), .A3(new_n465), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n757), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n695), .A2(new_n685), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n779), .A2(new_n311), .A3(new_n670), .A4(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(KEYINPUT50), .Z(new_n783));
  AND2_X1   g597(.A1(new_n781), .A2(new_n757), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n595), .A3(new_n465), .A4(new_n668), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n616), .A3(new_n615), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n776), .A2(new_n778), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n788), .A2(new_n713), .A3(new_n751), .A4(new_n712), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n780), .A2(new_n783), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n779), .A2(new_n650), .A3(new_n781), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT121), .Z(new_n795));
  INV_X1    g609(.A(new_n616), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n785), .A2(new_n796), .A3(new_n614), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n795), .A2(new_n464), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n780), .A2(new_n783), .A3(KEYINPUT51), .A4(new_n790), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n793), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n695), .A2(new_n650), .A3(new_n685), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n557), .A2(new_n595), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n557), .A2(new_n488), .A3(new_n652), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n803), .A2(new_n632), .B1(new_n781), .B2(new_n804), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n685), .A2(new_n695), .A3(new_n708), .A4(new_n714), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n803), .B2(new_n618), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n616), .A2(new_n424), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n318), .A2(new_n471), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT116), .B1(new_n318), .B2(new_n618), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n811), .B(new_n617), .C1(new_n312), .C2(new_n317), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n605), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n557), .A2(new_n490), .A3(new_n595), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT80), .B1(new_n597), .B2(new_n594), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n642), .B1(new_n818), .B2(new_n489), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n805), .A2(new_n807), .A3(new_n815), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n706), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n647), .B(KEYINPUT117), .Z(new_n822));
  AOI211_X1 g636(.A(new_n322), .B(new_n822), .C1(new_n378), .C2(new_n384), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n667), .A2(new_n821), .A3(new_n823), .A4(new_n751), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n641), .B1(new_n540), .B2(new_n666), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(KEYINPUT118), .A3(new_n821), .A4(new_n823), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n653), .A2(new_n718), .A3(new_n676), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT52), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n820), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n424), .A2(new_n463), .A3(new_n647), .ZN(new_n836));
  INV_X1    g650(.A(new_n628), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n597), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n641), .B(new_n724), .C1(new_n838), .C2(new_n717), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n730), .A2(new_n733), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT53), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n815), .A2(new_n819), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n704), .B1(new_n696), .B2(new_n631), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n715), .B1(new_n696), .B2(new_n617), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT52), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(new_n829), .B2(new_n830), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n842), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n730), .A2(new_n733), .A3(new_n839), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT54), .B1(new_n841), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n848), .B2(new_n849), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n833), .A2(new_n834), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n805), .A2(new_n807), .A3(KEYINPUT119), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n843), .B2(new_n844), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n733), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n726), .A2(new_n722), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n727), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n860), .B1(new_n864), .B2(new_n725), .ZN(new_n865));
  AND4_X1   g679(.A1(KEYINPUT53), .A2(new_n815), .A3(new_n819), .A4(new_n839), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n855), .A2(new_n859), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n853), .A2(new_n854), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n788), .A2(new_n721), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT48), .Z(new_n870));
  NAND4_X1  g684(.A1(new_n800), .A2(new_n852), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n683), .A2(new_n384), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n873), .A2(KEYINPUT49), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n873), .A2(KEYINPUT49), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT115), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n595), .A2(new_n321), .A3(new_n310), .A4(new_n745), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n874), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n878), .A2(new_n877), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n668), .A3(new_n670), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n872), .A2(new_n881), .ZN(G75));
  OR3_X1    g696(.A1(new_n273), .A2(KEYINPUT123), .A3(G952), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT123), .B1(new_n273), .B2(G952), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT124), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n379), .B1(new_n853), .B2(new_n867), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT56), .B1(new_n887), .B2(G210), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n243), .A2(new_n280), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n278), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n890), .B(new_n891), .Z(new_n892));
  OAI21_X1  g706(.A(new_n886), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n304), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(G51));
  XOR2_X1   g710(.A(new_n739), .B(KEYINPUT57), .Z(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n855), .A2(new_n859), .A3(new_n865), .A4(new_n866), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT54), .B1(new_n841), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n898), .B1(new_n900), .B2(new_n868), .ZN(new_n901));
  INV_X1    g715(.A(new_n692), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT125), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n853), .A2(new_n854), .A3(new_n867), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n854), .B1(new_n853), .B2(new_n867), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n692), .ZN(new_n908));
  INV_X1    g722(.A(new_n738), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n887), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n903), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n885), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n887), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n480), .A2(new_n460), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n885), .B1(new_n916), .B2(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(new_n609), .A2(new_n610), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n612), .B(KEYINPUT59), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n919), .B(new_n921), .C1(new_n904), .C2(new_n905), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n852), .B2(new_n868), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n922), .B(new_n886), .C1(new_n923), .C2(new_n919), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT60), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n853), .B2(new_n867), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(new_n579), .ZN(new_n929));
  INV_X1    g743(.A(new_n886), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n928), .B2(new_n639), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G66));
  NAND2_X1  g748(.A1(new_n272), .A2(new_n469), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(G953), .ZN(new_n936));
  INV_X1    g750(.A(new_n820), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n889), .B1(G898), .B2(new_n273), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  AOI21_X1  g754(.A(new_n759), .B1(new_n768), .B2(new_n769), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n730), .A2(new_n733), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n744), .A2(new_n655), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n721), .A2(new_n706), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n941), .A2(new_n273), .A3(new_n945), .A4(new_n830), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n511), .B(new_n474), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n946), .B(new_n948), .C1(new_n645), .C2(new_n273), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n950));
  INV_X1    g764(.A(new_n759), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n672), .A2(new_n830), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  INV_X1    g767(.A(new_n818), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n796), .A2(new_n614), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n757), .B1(new_n955), .B2(new_n808), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n954), .A2(new_n656), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n951), .A2(new_n953), .A3(new_n770), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n273), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n947), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n949), .A2(new_n950), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n273), .B1(G227), .B2(G900), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n949), .A2(new_n950), .A3(new_n960), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(G72));
  NOR2_X1   g780(.A1(new_n542), .A2(new_n516), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n830), .A2(new_n941), .A3(new_n937), .A4(new_n945), .ZN(new_n968));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n958), .B2(new_n820), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n660), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n912), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n841), .A2(new_n851), .ZN(new_n976));
  NOR4_X1   g790(.A1(new_n976), .A2(new_n660), .A3(new_n971), .A4(new_n967), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n975), .A2(new_n977), .ZN(G57));
endmodule


