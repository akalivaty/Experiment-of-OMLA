//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT3), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT65), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n477), .A2(KEYINPUT65), .A3(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n473), .B1(new_n479), .B2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n468), .A2(new_n471), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n468), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n471), .A2(G112), .ZN(new_n486));
  OR3_X1    g061(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(G2104), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n483), .B(new_n485), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n465), .A2(G126), .A3(new_n467), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n471), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n464), .A2(G2105), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n499), .A2(G102), .ZN(new_n500));
  OR3_X1    g075(.A1(new_n498), .A2(KEYINPUT69), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT4), .A2(G138), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n474), .A2(G138), .A3(new_n471), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n484), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT69), .B1(new_n498), .B2(new_n500), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT70), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n515), .B1(new_n520), .B2(KEYINPUT5), .ZN(new_n521));
  AOI211_X1 g096(.A(new_n513), .B(new_n514), .C1(new_n517), .C2(new_n519), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(new_n509), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT72), .B(G88), .Z(new_n525));
  OAI21_X1  g100(.A(new_n512), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n523), .A2(G62), .ZN(new_n528));
  NAND2_X1  g103(.A1(G75), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(G166));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(G63), .ZN(new_n533));
  NAND3_X1  g108(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT73), .B(G89), .Z(new_n537));
  NAND3_X1  g112(.A1(new_n523), .A2(new_n509), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n511), .A2(G51), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n532), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g119(.A1(new_n535), .A2(new_n542), .A3(KEYINPUT74), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(G168));
  AOI22_X1  g121(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT75), .Z(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n527), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n511), .A2(G52), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n524), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G171));
  NAND2_X1  g128(.A1(new_n511), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n524), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT71), .B1(new_n516), .B2(KEYINPUT5), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT70), .B(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n558), .B2(new_n514), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n520), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(new_n560), .A3(G56), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n556), .B1(new_n567), .B2(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT77), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(new_n511), .A2(G53), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n523), .A2(G91), .A3(new_n509), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n521), .B2(new_n522), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT78), .ZN(new_n582));
  XNOR2_X1  g157(.A(KEYINPUT79), .B(G65), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G78), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT80), .B1(new_n586), .B2(G651), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  AOI211_X1 g163(.A(new_n588), .B(new_n527), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n579), .B1(new_n587), .B2(new_n589), .ZN(G299));
  INV_X1    g165(.A(G171), .ZN(G301));
  NOR2_X1   g166(.A1(new_n544), .A2(new_n545), .ZN(G286));
  INV_X1    g167(.A(G166), .ZN(G303));
  OAI21_X1  g168(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n511), .A2(G49), .ZN(new_n595));
  INV_X1    g170(.A(G87), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n594), .B(new_n595), .C1(new_n596), .C2(new_n524), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT81), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G288));
  NAND3_X1  g174(.A1(new_n523), .A2(G86), .A3(new_n509), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT82), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n559), .A2(new_n560), .ZN(new_n606));
  INV_X1    g181(.A(G61), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n604), .A2(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(new_n511), .A2(G47), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  OAI221_X1 g188(.A(new_n611), .B1(new_n524), .B2(new_n612), .C1(new_n613), .C2(new_n527), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(G290));
  XNOR2_X1  g193(.A(KEYINPUT85), .B(G66), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n581), .A2(new_n582), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(G79), .A2(G543), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT84), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n527), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n559), .A2(new_n560), .A3(G92), .A4(new_n509), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT10), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n511), .A2(G54), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  NOR3_X1   g203(.A1(new_n624), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G171), .B2(new_n631), .ZN(G284));
  OAI21_X1  g208(.A(new_n632), .B1(G171), .B2(new_n631), .ZN(G321));
  NAND2_X1  g209(.A1(G299), .A2(new_n631), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G168), .B2(new_n631), .ZN(G297));
  XOR2_X1   g211(.A(G297), .B(KEYINPUT86), .Z(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n629), .B1(new_n638), .B2(G860), .ZN(G148));
  INV_X1    g214(.A(new_n566), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n640), .A2(G651), .A3(new_n564), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(new_n554), .C1(new_n555), .C2(new_n524), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(new_n631), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n630), .A2(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n631), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g221(.A1(new_n482), .A2(G123), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT87), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n484), .A2(G135), .ZN(new_n649));
  NOR2_X1   g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n474), .A2(new_n499), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT13), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n657), .ZN(G156));
  NOR2_X1   g233(.A1(KEYINPUT89), .A2(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT90), .B(G2438), .Z(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT15), .B(G2435), .Z(new_n663));
  AOI21_X1  g238(.A(new_n659), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(KEYINPUT89), .B2(KEYINPUT14), .ZN(new_n666));
  XOR2_X1   g241(.A(G2451), .B(G2454), .Z(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(G2443), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT88), .B(KEYINPUT16), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2446), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1341), .B(G1348), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT91), .Z(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(G14), .C1(new_n673), .C2(new_n672), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT92), .ZN(new_n679));
  XOR2_X1   g254(.A(G2067), .B(G2678), .Z(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT17), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT18), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(KEYINPUT18), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n687), .B(new_n689), .Z(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n692), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n696), .A2(KEYINPUT20), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n698), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n700), .A2(new_n692), .A3(new_n695), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n699), .B(new_n701), .C1(KEYINPUT20), .C2(new_n696), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1986), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1981), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1991), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n704), .B(new_n707), .ZN(G229));
  AOI22_X1  g283(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(new_n471), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT97), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n484), .A2(G139), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n499), .A2(G103), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT25), .Z(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G33), .B(new_n715), .S(G29), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G2072), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G35), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n717), .B1(G2090), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G5), .A2(G16), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G171), .B2(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G1961), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n568), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(G19), .ZN(new_n729));
  INV_X1    g304(.A(G1341), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n723), .A2(new_n726), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT98), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT26), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n499), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n482), .A2(G129), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G32), .B(new_n739), .S(G29), .Z(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT99), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G11), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT101), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n718), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n482), .A2(G128), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n484), .A2(G140), .ZN(new_n750));
  NOR2_X1   g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(new_n471), .B2(G116), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G29), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(KEYINPUT96), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(KEYINPUT96), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n748), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  INV_X1    g333(.A(G2078), .ZN(new_n759));
  NOR2_X1   g334(.A1(G164), .A2(new_n718), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G27), .B2(new_n718), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT30), .B(G28), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(new_n718), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT24), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n765), .A2(G34), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(G34), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n718), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G160), .B2(new_n718), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n764), .B1(new_n652), .B2(new_n718), .C1(G2084), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G2084), .B2(new_n769), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n762), .B(new_n771), .C1(new_n759), .C2(new_n761), .ZN(new_n772));
  NOR2_X1   g347(.A1(G4), .A2(G16), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n629), .B2(G16), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT95), .B(G1348), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n744), .A2(new_n746), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n727), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n727), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G1966), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT100), .Z(new_n782));
  OAI22_X1  g357(.A1(new_n725), .A2(G1961), .B1(new_n780), .B2(G1966), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n778), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G299), .ZN(new_n785));
  OAI21_X1  g360(.A(KEYINPUT23), .B1(new_n785), .B2(new_n727), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n727), .A2(G20), .ZN(new_n787));
  MUX2_X1   g362(.A(KEYINPUT23), .B(new_n786), .S(new_n787), .Z(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G1956), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G1956), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n784), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2090), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n721), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT102), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n482), .A2(G119), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n484), .A2(G131), .ZN(new_n796));
  NOR2_X1   g371(.A1(G95), .A2(G2105), .ZN(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G25), .B(new_n799), .S(G29), .Z(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT35), .B(G1991), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n800), .B(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n614), .B(KEYINPUT83), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(new_n727), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n727), .B2(G24), .ZN(new_n806));
  INV_X1    g381(.A(G1986), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n727), .A2(G23), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n597), .B(KEYINPUT93), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n809), .B1(new_n811), .B2(new_n727), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT33), .B(G1976), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n727), .A2(G6), .ZN(new_n815));
  INV_X1    g390(.A(G305), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n727), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n727), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n727), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT94), .B(G1971), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n814), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n808), .B1(new_n824), .B2(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n806), .A2(new_n807), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n825), .B(new_n826), .C1(KEYINPUT34), .C2(new_n824), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT36), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n791), .A2(new_n794), .A3(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  INV_X1    g405(.A(KEYINPUT104), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n559), .A2(new_n560), .A3(G67), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT103), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(new_n832), .B2(new_n834), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n836), .A2(new_n837), .A3(new_n527), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n523), .A2(G93), .A3(new_n509), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n511), .A2(G55), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n831), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n837), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n843), .A2(G651), .A3(new_n835), .ZN(new_n844));
  INV_X1    g419(.A(new_n841), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT104), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n629), .A2(G559), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n568), .B1(new_n842), .B2(new_n846), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n838), .A2(new_n841), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n642), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n853), .B(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n850), .B1(new_n858), .B2(G860), .ZN(G145));
  XNOR2_X1  g434(.A(new_n715), .B(KEYINPUT105), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n652), .ZN(new_n861));
  XNOR2_X1  g436(.A(G160), .B(G162), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n498), .A2(new_n500), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n505), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n482), .A2(G130), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n484), .A2(G142), .ZN(new_n867));
  NOR2_X1   g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n865), .B(new_n870), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n655), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n739), .B(new_n753), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n799), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n872), .B(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n863), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n863), .A2(new_n875), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g455(.A1(new_n848), .A2(new_n631), .ZN(new_n881));
  NOR2_X1   g456(.A1(G290), .A2(G166), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n804), .A2(G303), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n816), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(G290), .A2(G166), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n804), .A2(G303), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(G305), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n811), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(new_n887), .A3(new_n810), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT42), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n857), .B(new_n644), .ZN(new_n893));
  NAND2_X1  g468(.A1(G299), .A2(new_n630), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n629), .B(new_n579), .C1(new_n587), .C2(new_n589), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n894), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n894), .B2(new_n895), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT106), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n894), .A2(new_n898), .A3(new_n895), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n897), .B1(new_n893), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n892), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n881), .B1(new_n907), .B2(new_n631), .ZN(G295));
  OAI21_X1  g483(.A(new_n881), .B1(new_n907), .B2(new_n631), .ZN(G331));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n902), .A2(new_n903), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n896), .A2(KEYINPUT41), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n894), .A2(new_n898), .A3(new_n895), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n911), .B1(new_n914), .B2(KEYINPUT106), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n838), .A2(new_n831), .A3(new_n841), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT104), .B1(new_n844), .B2(new_n845), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n642), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n568), .B1(new_n841), .B2(new_n838), .ZN(new_n919));
  AOI21_X1  g494(.A(G168), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n854), .A2(new_n856), .A3(G286), .ZN(new_n921));
  OAI21_X1  g496(.A(G301), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(G286), .B1(new_n854), .B2(new_n856), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(G168), .A3(new_n919), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(G171), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT107), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n884), .A2(new_n887), .A3(new_n810), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n810), .B1(new_n884), .B2(new_n887), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n894), .A3(new_n895), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n923), .A2(new_n924), .A3(G171), .ZN(new_n932));
  AOI21_X1  g507(.A(G171), .B1(new_n923), .B2(new_n924), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n905), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n927), .A2(new_n930), .A3(new_n931), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n922), .A2(new_n914), .A3(new_n925), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n934), .B2(new_n896), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n939), .B2(new_n891), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n910), .B1(new_n941), .B2(KEYINPUT43), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n927), .A2(new_n931), .A3(new_n936), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n891), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n945), .A2(new_n946), .A3(new_n877), .A4(new_n937), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n943), .B1(new_n942), .B2(new_n947), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n937), .A2(new_n940), .A3(new_n946), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n877), .A3(new_n937), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(KEYINPUT43), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n948), .A2(new_n949), .B1(KEYINPUT44), .B2(new_n952), .ZN(G397));
  XNOR2_X1  g528(.A(KEYINPUT109), .B(G1384), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n864), .B2(new_n505), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(KEYINPUT45), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n477), .A2(KEYINPUT65), .A3(G2105), .ZN(new_n958));
  OAI211_X1 g533(.A(G40), .B(new_n472), .C1(new_n958), .C2(new_n478), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G2067), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n753), .B(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n739), .B(G1996), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT110), .Z(new_n967));
  NOR2_X1   g542(.A1(new_n799), .A2(new_n801), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n753), .A2(G2067), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n961), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT125), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n961), .A2(G1996), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT126), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT46), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n973), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n960), .B1(new_n739), .B2(new_n964), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n976), .B(new_n977), .C1(new_n974), .C2(KEYINPUT46), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n799), .B(new_n802), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n967), .B1(new_n961), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n804), .A2(new_n807), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n961), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT48), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n972), .B(new_n979), .C1(new_n981), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT112), .B1(new_n600), .B2(new_n602), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n600), .A2(KEYINPUT112), .A3(new_n602), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(new_n609), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(G1981), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  INV_X1    g568(.A(new_n989), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(new_n987), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n995), .B2(new_n609), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT113), .B1(G305), .B2(G1981), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n992), .B(KEYINPUT114), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n816), .A2(new_n993), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n990), .A2(G1981), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(KEYINPUT113), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1002), .A2(KEYINPUT114), .A3(new_n1003), .A4(new_n992), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n864), .B2(new_n505), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(G8), .B1(new_n1006), .B2(new_n959), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n999), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n811), .B2(G1976), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1010), .B(new_n1011), .C1(G1976), .C2(new_n598), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G166), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(KEYINPUT111), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1017), .A2(KEYINPUT111), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1016), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n507), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n959), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n955), .A2(KEYINPUT45), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1971), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n959), .B1(new_n1006), .B2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n507), .A2(new_n1034), .A3(new_n1024), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(G2090), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1023), .B1(new_n1037), .B2(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n959), .B1(new_n1034), .B2(new_n1005), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1041), .A2(new_n792), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1022), .A2(new_n1042), .A3(new_n1015), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1014), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1030), .B2(G2078), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1047));
  INV_X1    g622(.A(G1961), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1028), .B(KEYINPUT116), .C1(KEYINPUT45), .C2(new_n1005), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1052), .B2(new_n959), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1045), .A2(G2078), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1050), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1046), .A2(new_n1049), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G171), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT124), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n957), .A2(G40), .A3(new_n472), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n477), .A2(G2105), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n1029), .A4(new_n1054), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(G301), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1065), .A3(G171), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1059), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(KEYINPUT54), .C1(G171), .C2(new_n1057), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n1073));
  INV_X1    g648(.A(G2084), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1050), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1075));
  INV_X1    g650(.A(G1966), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1074), .A2(new_n1041), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1073), .B1(new_n1077), .B2(new_n1015), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT51), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(G168), .C1(G2084), .C2(new_n1047), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1077), .A2(G168), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT51), .B(new_n1078), .C1(new_n1082), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AND4_X1   g662(.A1(new_n1044), .A2(new_n1069), .A3(new_n1072), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1036), .B2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g666(.A(KEYINPUT119), .B(G1956), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1091), .A2(new_n1092), .B1(new_n1030), .B2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(G299), .B(KEYINPUT57), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1006), .A2(new_n959), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1047), .A2(new_n1100), .B1(new_n962), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n630), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1097), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1097), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1097), .A2(new_n1107), .A3(KEYINPUT61), .A4(new_n1098), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n629), .A2(KEYINPUT121), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n629), .A2(KEYINPUT121), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1102), .A2(KEYINPUT60), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1112), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1110), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT122), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1099), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1113), .A2(new_n1114), .A3(new_n1122), .A4(new_n1116), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1030), .A2(G1996), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT58), .B(G1341), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1101), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n568), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT59), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1118), .A2(new_n1121), .A3(new_n1123), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1104), .B1(new_n1109), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1014), .A2(new_n1043), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1038), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1084), .A2(new_n1086), .A3(new_n1131), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1088), .A2(new_n1130), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1022), .B1(new_n1042), .B2(new_n1015), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1009), .A2(new_n1139), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1140), .A2(KEYINPUT117), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1077), .A2(new_n1015), .A3(G286), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1140), .B2(KEYINPUT117), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT63), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1014), .A2(new_n1145), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1044), .A2(new_n1146), .B1(new_n1043), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(G1976), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1009), .A2(new_n1149), .A3(new_n598), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1000), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(KEYINPUT115), .A3(new_n1000), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(new_n1008), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1144), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT118), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1144), .A2(new_n1148), .A3(new_n1155), .A4(KEYINPUT118), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1138), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n961), .B1(new_n1161), .B2(new_n982), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n981), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n986), .B1(new_n1160), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g739(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n1166));
  INV_X1    g740(.A(new_n950), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g742(.A(G227), .ZN(new_n1169));
  NOR2_X1   g743(.A1(G229), .A2(new_n460), .ZN(new_n1170));
  NAND4_X1  g744(.A1(new_n676), .A2(new_n1169), .A3(new_n879), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g745(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n1168), .A2(KEYINPUT127), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n1174));
  OAI21_X1  g748(.A(new_n1174), .B1(new_n952), .B2(new_n1171), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1175), .ZN(G308));
  NAND2_X1  g750(.A1(new_n1168), .A2(new_n1172), .ZN(G225));
endmodule


