//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT91), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT91), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT92), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n207), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT93), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(KEYINPUT93), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT92), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(new_n204), .B2(new_n206), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G1gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n211), .A2(new_n213), .A3(new_n214), .A4(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n217), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n205), .B(new_n203), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n216), .A2(G1gat), .B1(new_n220), .B2(KEYINPUT16), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT93), .B(new_n212), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT94), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n218), .A2(new_n222), .A3(KEYINPUT94), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G71gat), .A2(G78gat), .ZN(new_n228));
  OR2_X1    g027(.A1(G71gat), .A2(G78gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT9), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G57gat), .ZN(new_n232));
  OR3_X1    g031(.A1(new_n232), .A2(KEYINPUT98), .A3(G64gat), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT98), .B1(new_n232), .B2(G64gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G64gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G57gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n231), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n232), .A2(G64gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT9), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n228), .A3(new_n229), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT21), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(G183gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n247), .A3(new_n244), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n248), .A3(new_n250), .ZN(new_n253));
  XNOR2_X1  g052(.A(G127gat), .B(G155gat), .ZN(new_n254));
  INV_X1    g053(.A(G211gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n252), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n252), .B2(new_n253), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n243), .A2(KEYINPUT21), .ZN(new_n260));
  NAND2_X1  g059(.A1(G231gat), .A2(G233gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n261), .B(KEYINPUT99), .Z(new_n262));
  XNOR2_X1  g061(.A(new_n260), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OR3_X1    g063(.A1(new_n258), .A2(new_n259), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(new_n258), .B2(new_n259), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G43gat), .B(G50gat), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n268), .A2(KEYINPUT15), .ZN(new_n269));
  OR3_X1    g068(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G29gat), .A2(G36gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT89), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n272), .B(new_n274), .C1(KEYINPUT15), .C2(new_n268), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n270), .B2(new_n276), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT17), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT90), .A3(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n283), .A2(KEYINPUT90), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(KEYINPUT90), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G85gat), .A2(G92gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT7), .ZN(new_n290));
  NAND2_X1  g089(.A1(G99gat), .A2(G106gat), .ZN(new_n291));
  INV_X1    g090(.A(G85gat), .ZN(new_n292));
  INV_X1    g091(.A(G92gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(KEYINPUT8), .A2(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G99gat), .B(G106gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT100), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT100), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n290), .A2(new_n299), .A3(new_n296), .A4(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n288), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n303), .B(new_n304), .C1(new_n282), .C2(new_n302), .ZN(new_n305));
  XOR2_X1   g104(.A(G134gat), .B(G162gat), .Z(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G190gat), .B(G218gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(KEYINPUT101), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n307), .B(new_n311), .Z(new_n312));
  NAND2_X1  g111(.A1(new_n267), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G230gat), .ZN(new_n314));
  INV_X1    g113(.A(G233gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT10), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n243), .B1(new_n298), .B2(new_n300), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n297), .A2(new_n242), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n301), .A2(KEYINPUT10), .A3(new_n243), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n318), .A2(new_n319), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n316), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT102), .ZN(new_n327));
  XNOR2_X1  g126(.A(G120gat), .B(G148gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G204gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n327), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT18), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(KEYINPUT96), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n288), .A2(new_n223), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n225), .A2(new_n226), .A3(new_n281), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT95), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n225), .A2(KEYINPUT95), .A3(new_n226), .A4(new_n281), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G229gat), .A2(G233gat), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n336), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n335), .A2(KEYINPUT96), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n342), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n227), .A2(new_n282), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n344), .B(KEYINPUT13), .Z(new_n350));
  AOI22_X1  g149(.A1(new_n345), .A2(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(KEYINPUT18), .A3(new_n344), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT97), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n345), .B2(new_n346), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT11), .B(G169gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G197gat), .ZN(new_n356));
  XOR2_X1   g155(.A(G113gat), .B(G141gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT87), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT12), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n351), .B(new_n352), .C1(new_n354), .C2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n347), .A2(new_n344), .A3(new_n337), .ZN(new_n362));
  INV_X1    g161(.A(new_n336), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n346), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n360), .B1(new_n364), .B2(KEYINPUT97), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n352), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n313), .A2(new_n334), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G197gat), .B(G204gat), .ZN(new_n372));
  INV_X1    g171(.A(G218gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n255), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(KEYINPUT22), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G211gat), .B(G218gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(KEYINPUT29), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT3), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n379), .B2(new_n378), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(G155gat), .B2(G162gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G141gat), .B(G148gat), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT2), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(G155gat), .B2(G162gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G155gat), .B(G162gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n388), .B(new_n383), .C1(new_n384), .C2(new_n386), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n381), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n377), .B(KEYINPUT72), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n394), .A2(G228gat), .A3(G233gat), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n393), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n377), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT80), .B(new_n393), .C1(new_n378), .C2(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G228gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n315), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(G22gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n401), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT31), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G50gat), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n401), .A2(new_n410), .ZN(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n412), .B(new_n415), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n415), .B(KEYINPUT79), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n401), .A2(new_n410), .A3(new_n411), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n411), .B1(new_n401), .B2(new_n410), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT67), .ZN(new_n425));
  NAND2_X1  g224(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G169gat), .A2(G176gat), .ZN(new_n431));
  INV_X1    g230(.A(G169gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n329), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT23), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n425), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G183gat), .A2(G190gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(KEYINPUT24), .ZN(new_n438));
  AND2_X1   g237(.A1(G183gat), .A2(G190gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n441), .B2(KEYINPUT24), .ZN(new_n442));
  AND2_X1   g241(.A1(G169gat), .A2(G176gat), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(KEYINPUT23), .B2(new_n428), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n434), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n433), .A2(new_n446), .A3(new_n426), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT67), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n436), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT25), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n430), .A2(new_n435), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT25), .A4(new_n442), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT25), .ZN(new_n455));
  INV_X1    g254(.A(new_n440), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(KEYINPUT24), .A3(new_n437), .ZN(new_n457));
  INV_X1    g256(.A(new_n438), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT68), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n451), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT26), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n433), .A2(new_n463), .A3(new_n431), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n428), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT69), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT27), .B(G183gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT28), .B1(new_n469), .B2(G190gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT28), .ZN(new_n471));
  INV_X1    g270(.A(G190gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT29), .B1(new_n462), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(G226gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(new_n315), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT73), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n475), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n478), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT73), .ZN(new_n482));
  INV_X1    g281(.A(new_n478), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n451), .A2(new_n461), .B1(new_n467), .B2(new_n474), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n482), .B(new_n483), .C1(new_n484), .C2(KEYINPUT29), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n479), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n395), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n483), .B1(new_n484), .B2(KEYINPUT29), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT74), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n488), .A2(new_n489), .B1(new_n478), .B2(new_n480), .ZN(new_n490));
  INV_X1    g289(.A(new_n377), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT74), .B(new_n483), .C1(new_n484), .C2(KEYINPUT29), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G64gat), .B(G92gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(G36gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT75), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(new_n212), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n494), .A2(new_n499), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n487), .A2(new_n493), .A3(new_n498), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT77), .ZN(new_n505));
  XNOR2_X1  g304(.A(G113gat), .B(G120gat), .ZN(new_n506));
  OAI21_X1  g305(.A(G127gat), .B1(new_n506), .B2(KEYINPUT1), .ZN(new_n507));
  INV_X1    g306(.A(G120gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G113gat), .ZN(new_n509));
  INV_X1    g308(.A(G113gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G120gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT1), .ZN(new_n513));
  INV_X1    g312(.A(G127gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n507), .A2(new_n515), .A3(G134gat), .ZN(new_n516));
  AOI21_X1  g315(.A(G134gat), .B1(new_n507), .B2(new_n515), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n505), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G134gat), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n506), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n514), .B1(new_n512), .B2(new_n513), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n515), .A3(G134gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT77), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n392), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G225gat), .A2(G233gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n392), .A2(new_n522), .A3(new_n523), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n525), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT39), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n504), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n518), .A2(new_n524), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n393), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n526), .A3(new_n528), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT84), .A3(KEYINPUT39), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n404), .A3(new_n397), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT4), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n528), .B(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n527), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n532), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT0), .B(G57gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G85gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G1gat), .B(G29gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n544), .B(new_n545), .Z(new_n546));
  XOR2_X1   g345(.A(new_n546), .B(KEYINPUT83), .Z(new_n547));
  OAI211_X1 g346(.A(new_n531), .B(new_n527), .C1(new_n538), .C2(new_n540), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT85), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT40), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n528), .B(KEYINPUT4), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n526), .A3(new_n537), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n527), .B1(new_n525), .B2(new_n529), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT5), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT5), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n547), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AND4_X1   g359(.A1(new_n500), .A2(new_n503), .A3(new_n551), .A4(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n550), .A2(KEYINPUT40), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n424), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n486), .A2(new_n395), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT37), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT38), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n487), .A2(new_n493), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n499), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT6), .ZN(new_n574));
  INV_X1    g373(.A(new_n558), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n557), .B1(new_n553), .B2(new_n554), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n546), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n560), .B(new_n574), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(KEYINPUT6), .A3(new_n578), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n502), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n565), .B1(new_n573), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n571), .A2(new_n499), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n570), .B1(new_n487), .B2(new_n493), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT38), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR4_X1   g384(.A1(new_n575), .A2(new_n576), .A3(new_n574), .A4(new_n546), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n556), .A2(new_n558), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT6), .B1(new_n587), .B2(new_n546), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n588), .B2(new_n560), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n589), .A2(KEYINPUT86), .A3(new_n572), .A4(new_n502), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n564), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT78), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(new_n587), .B2(new_n546), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n577), .A2(KEYINPUT78), .A3(new_n578), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n588), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n580), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n503), .A2(new_n500), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n424), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n601));
  XNOR2_X1  g400(.A(G15gat), .B(G43gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G71gat), .ZN(new_n603));
  INV_X1    g402(.A(G99gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n522), .A2(new_n523), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n462), .A2(new_n608), .A3(new_n475), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT70), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n480), .A2(new_n607), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT70), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n484), .A2(new_n612), .A3(new_n608), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G227gat), .A2(G233gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT64), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT65), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n614), .A2(KEYINPUT71), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT71), .B1(new_n614), .B2(new_n617), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT32), .B(new_n606), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n614), .A2(new_n616), .ZN(new_n621));
  INV_X1    g420(.A(new_n614), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n617), .A2(KEYINPUT34), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n621), .A2(KEYINPUT34), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(KEYINPUT32), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n614), .A2(new_n617), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT71), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n614), .A2(KEYINPUT71), .A3(new_n617), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n605), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n620), .B(new_n624), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI22_X1  g433(.A1(new_n618), .A2(new_n619), .B1(KEYINPUT32), .B2(new_n625), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n605), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n624), .B1(new_n636), .B2(new_n620), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n601), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n620), .B1(new_n631), .B2(new_n632), .ZN(new_n639));
  INV_X1    g438(.A(new_n624), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(KEYINPUT36), .A3(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n592), .A2(new_n600), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n633), .A3(new_n423), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT35), .B1(new_n599), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n634), .A2(new_n637), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n589), .B1(new_n500), .B2(new_n503), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT35), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .A4(new_n423), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n371), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n597), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n209), .ZN(G1324gat));
  XNOR2_X1  g454(.A(KEYINPUT16), .B(G8gat), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n653), .ZN(new_n659));
  INV_X1    g458(.A(new_n598), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n661), .A2(new_n657), .A3(new_n656), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(KEYINPUT103), .Z(new_n663));
  NOR2_X1   g462(.A1(new_n657), .A2(G8gat), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n658), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(G1325gat));
  AOI21_X1  g464(.A(G15gat), .B1(new_n659), .B2(new_n647), .ZN(new_n666));
  INV_X1    g465(.A(new_n643), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G15gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT104), .Z(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n659), .B2(new_n669), .ZN(G1326gat));
  NOR2_X1   g469(.A1(new_n653), .A2(new_n423), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT43), .B(G22gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  AOI21_X1  g472(.A(new_n312), .B1(new_n644), .B2(new_n651), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n370), .A2(new_n267), .A3(new_n334), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n676), .A2(G29gat), .A3(new_n597), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT105), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT45), .Z(new_n679));
  NOR2_X1   g478(.A1(new_n312), .A2(KEYINPUT44), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n646), .A2(new_n650), .A3(KEYINPUT106), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT106), .B1(new_n646), .B2(new_n650), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n644), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n644), .B(new_n686), .C1(new_n682), .C2(new_n683), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n681), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n675), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n597), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G29gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n696), .ZN(G1328gat));
  NAND2_X1  g496(.A1(new_n693), .A2(new_n660), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G36gat), .ZN(new_n699));
  OR3_X1    g498(.A1(new_n676), .A2(G36gat), .A3(new_n598), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(KEYINPUT108), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n701), .A2(KEYINPUT108), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n699), .B(new_n704), .C1(new_n702), .C2(new_n700), .ZN(G1329gat));
  NAND3_X1  g504(.A1(new_n693), .A2(G43gat), .A3(new_n667), .ZN(new_n706));
  INV_X1    g505(.A(G43gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n647), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n676), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g510(.A(G50gat), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n423), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n675), .B(new_n713), .C1(new_n688), .C2(new_n690), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n676), .B2(new_n423), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT109), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(new_n718), .A3(new_n715), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g520(.A(new_n313), .B1(new_n685), .B2(new_n687), .ZN(new_n722));
  INV_X1    g521(.A(new_n334), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n369), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n597), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(new_n232), .ZN(G1332gat));
  AND2_X1   g526(.A1(new_n722), .A2(new_n724), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n660), .B1(new_n729), .B2(new_n236), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT110), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT111), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n732), .B(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n729), .A3(new_n236), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n725), .B2(new_n708), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n722), .A2(G71gat), .A3(new_n667), .A4(new_n724), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT112), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n744), .A3(new_n741), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n743), .A2(KEYINPUT50), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT50), .B1(new_n743), .B2(new_n745), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n728), .A2(new_n424), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  INV_X1    g549(.A(new_n691), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n267), .A2(new_n369), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n334), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n755), .A2(new_n292), .A3(new_n597), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n641), .A2(new_n633), .A3(new_n423), .ZN(new_n759));
  AOI22_X1  g558(.A1(new_n580), .A2(new_n596), .B1(new_n503), .B2(new_n500), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n649), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n641), .A2(new_n423), .A3(new_n649), .A4(new_n633), .ZN(new_n762));
  INV_X1    g561(.A(new_n589), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n598), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n758), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n646), .A2(new_n650), .A3(KEYINPUT106), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n564), .A2(new_n591), .B1(new_n638), .B2(new_n642), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n600), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n757), .B1(new_n769), .B2(new_n312), .ZN(new_n770));
  INV_X1    g569(.A(new_n312), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n684), .A2(KEYINPUT113), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n752), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n770), .A2(KEYINPUT51), .A3(new_n772), .A4(new_n752), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n694), .A3(new_n334), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n756), .B1(new_n292), .B2(new_n778), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n751), .A2(new_n660), .A3(new_n754), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n598), .A2(G92gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n777), .A2(new_n334), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n773), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n723), .B1(new_n787), .B2(new_n776), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n780), .A2(G92gat), .B1(new_n788), .B2(new_n783), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n789), .B2(new_n782), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n755), .B2(new_n643), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n777), .A2(new_n604), .A3(new_n334), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n708), .B2(new_n792), .ZN(G1338gat));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n424), .B(new_n754), .C1(new_n688), .C2(new_n690), .ZN(new_n795));
  XOR2_X1   g594(.A(KEYINPUT115), .B(G106gat), .Z(new_n796));
  AND2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n723), .A2(G106gat), .A3(new_n423), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n775), .B2(new_n776), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n797), .A2(new_n800), .A3(KEYINPUT53), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n776), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n798), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n795), .A2(new_n796), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n794), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n800), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n802), .A3(new_n805), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n799), .B1(new_n787), .B2(new_n776), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n797), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n811), .A3(KEYINPUT116), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n807), .A2(new_n812), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n320), .A2(new_n316), .A3(new_n321), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n322), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(KEYINPUT54), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n815), .A2(new_n322), .A3(KEYINPUT117), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n322), .A2(new_n818), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n820), .A2(KEYINPUT118), .A3(new_n332), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT118), .B1(new_n820), .B2(new_n332), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n817), .A2(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI221_X1 g624(.A(KEYINPUT55), .B1(new_n821), .B2(new_n822), .C1(new_n817), .C2(new_n819), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n323), .A2(new_n325), .A3(new_n333), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n361), .B2(new_n368), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n349), .A2(new_n350), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n343), .A2(new_n344), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n358), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n360), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n367), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n723), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n312), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n312), .A2(new_n834), .A3(new_n828), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n267), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n313), .A2(new_n334), .A3(new_n369), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n645), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n660), .A2(new_n597), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n370), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(new_n510), .ZN(G1340gat));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n723), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(new_n508), .ZN(G1341gat));
  INV_X1    g646(.A(new_n267), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n514), .A2(KEYINPUT119), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n849), .B(new_n850), .Z(G1342gat));
  NAND4_X1  g650(.A1(new_n841), .A2(new_n519), .A3(new_n771), .A4(new_n842), .ZN(new_n852));
  OR2_X1    g651(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n843), .B2(new_n312), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(KEYINPUT56), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(G1343gat));
  INV_X1    g655(.A(G141gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n424), .B1(new_n838), .B2(new_n839), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT57), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n424), .C1(new_n838), .C2(new_n839), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n643), .A2(new_n842), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n859), .A2(KEYINPUT120), .A3(new_n861), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n857), .B1(new_n868), .B2(new_n369), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n858), .A2(new_n862), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n857), .A3(new_n369), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT58), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n864), .B2(new_n370), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n871), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(G1344gat));
  INV_X1    g676(.A(G148gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n870), .A2(new_n878), .A3(new_n334), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT121), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n334), .A3(new_n861), .ZN(new_n881));
  OAI21_X1  g680(.A(G148gat), .B1(new_n881), .B2(new_n862), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT59), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(KEYINPUT122), .A3(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n723), .B1(new_n866), .B2(new_n867), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(KEYINPUT59), .A3(new_n878), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n880), .B1(new_n887), .B2(new_n889), .ZN(G1345gat));
  AOI21_X1  g689(.A(G155gat), .B1(new_n870), .B2(new_n267), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n267), .A2(G155gat), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT123), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n868), .B2(new_n893), .ZN(G1346gat));
  AOI21_X1  g693(.A(G162gat), .B1(new_n870), .B2(new_n771), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n312), .B1(new_n866), .B2(new_n867), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n694), .A2(new_n598), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n841), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n370), .ZN(new_n900));
  XNOR2_X1  g699(.A(KEYINPUT124), .B(G169gat), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n900), .B(new_n901), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n899), .A2(new_n723), .ZN(new_n903));
  XNOR2_X1  g702(.A(KEYINPUT125), .B(G176gat), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(G1349gat));
  INV_X1    g704(.A(new_n899), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n468), .A3(new_n267), .ZN(new_n907));
  OAI21_X1  g706(.A(G183gat), .B1(new_n899), .B2(new_n848), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n771), .ZN(new_n911));
  NOR2_X1   g710(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n912));
  AND2_X1   g711(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n911), .B2(new_n913), .ZN(G1351gat));
  AND2_X1   g714(.A1(new_n643), .A2(new_n898), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n859), .A2(new_n861), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n370), .ZN(new_n918));
  INV_X1    g717(.A(new_n858), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n916), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(G197gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n921), .B2(new_n370), .ZN(G1352gat));
  INV_X1    g721(.A(new_n920), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n331), .A3(new_n334), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(KEYINPUT126), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n925), .A2(KEYINPUT126), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR4_X1   g727(.A1(new_n881), .A2(new_n694), .A3(new_n598), .A4(new_n667), .ZN(new_n929));
  OAI221_X1 g728(.A(new_n928), .B1(new_n926), .B2(new_n924), .C1(new_n331), .C2(new_n929), .ZN(G1353gat));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  OAI221_X1 g730(.A(G211gat), .B1(new_n931), .B2(KEYINPUT63), .C1(new_n917), .C2(new_n848), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n931), .A2(KEYINPUT63), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n923), .A2(new_n255), .A3(new_n267), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G1354gat));
  NAND3_X1  g736(.A1(new_n923), .A2(new_n373), .A3(new_n771), .ZN(new_n938));
  OAI21_X1  g737(.A(G218gat), .B1(new_n917), .B2(new_n312), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1355gat));
endmodule


