//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  NAND2_X1  g001(.A1(G43gat), .A2(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT90), .B(G50gat), .Z(new_n204));
  OAI211_X1 g003(.A(new_n202), .B(new_n203), .C1(new_n204), .C2(G43gat), .ZN(new_n205));
  OR2_X1    g004(.A1(G43gat), .A2(G50gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n206), .B2(new_n203), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT89), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n213), .A2(KEYINPUT89), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n207), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n225), .A2(G1gat), .ZN(new_n226));
  INV_X1    g025(.A(G8gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n227), .B1(new_n226), .B2(new_n229), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n224), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n223), .A2(KEYINPUT17), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n236), .A3(new_n222), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT91), .B1(new_n231), .B2(new_n232), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n226), .A2(new_n229), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G8gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n230), .A3(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n235), .A2(new_n237), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n234), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n242), .ZN(new_n247));
  INV_X1    g046(.A(new_n237), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n236), .B1(new_n216), .B2(new_n222), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT92), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n245), .A2(new_n251), .A3(KEYINPUT18), .A4(new_n246), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n224), .B(new_n233), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n246), .B(KEYINPUT13), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G113gat), .B(G141gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G169gat), .B(G197gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT12), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n254), .A2(new_n255), .A3(new_n258), .A4(new_n265), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G197gat), .B(G204gat), .ZN(new_n271));
  AND2_X1   g070(.A1(G211gat), .A2(G218gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(KEYINPUT22), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G155gat), .B(G162gat), .ZN(new_n276));
  INV_X1    g075(.A(G148gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(G141gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n278), .B2(KEYINPUT77), .ZN(new_n279));
  XNOR2_X1  g078(.A(G141gat), .B(G148gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(KEYINPUT77), .B2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT78), .B(G155gat), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G162gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT2), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n280), .A2(KEYINPUT2), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n288), .A2(new_n276), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n275), .B1(new_n291), .B2(KEYINPUT29), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n287), .B1(new_n275), .B2(KEYINPUT29), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(new_n289), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(G228gat), .A3(G233gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(KEYINPUT80), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n286), .A2(new_n299), .A3(new_n289), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n293), .ZN(new_n302));
  NAND2_X1  g101(.A1(G228gat), .A2(G233gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n292), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G22gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G78gat), .B(G106gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT31), .B(G50gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT83), .ZN(new_n311));
  INV_X1    g110(.A(G22gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n312), .A3(new_n304), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n306), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n310), .A2(KEYINPUT83), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n315), .B(KEYINPUT84), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n306), .A2(new_n311), .A3(new_n313), .A4(new_n316), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT23), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT66), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(KEYINPUT23), .ZN(new_n325));
  INV_X1    g124(.A(G169gat), .ZN(new_n326));
  INV_X1    g125(.A(G176gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(KEYINPUT67), .B(G190gat), .Z(new_n330));
  INV_X1    g129(.A(G183gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n321), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n322), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT26), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n326), .B2(new_n327), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n338), .B1(new_n322), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT27), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(KEYINPUT68), .ZN(new_n343));
  NAND2_X1  g142(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n331), .A2(KEYINPUT27), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n343), .A2(new_n344), .B1(new_n345), .B2(KEYINPUT68), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n330), .C1(new_n343), .C2(new_n344), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT27), .B(G183gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n330), .A2(KEYINPUT28), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n341), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n337), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT64), .ZN(new_n354));
  OAI221_X1 g153(.A(new_n335), .B1(G183gat), .B2(G190gat), .C1(new_n333), .C2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(new_n354), .B2(new_n333), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT65), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n358), .A2(new_n321), .A3(new_n359), .A4(new_n329), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n353), .B2(new_n360), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n275), .ZN(new_n366));
  INV_X1    g165(.A(new_n275), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n363), .B(new_n367), .C1(new_n362), .C2(new_n364), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G8gat), .B(G36gat), .Z(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT76), .ZN(new_n371));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n373), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n366), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n376), .ZN(new_n377));
  OR3_X1    g176(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n373), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT71), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G113gat), .ZN(new_n384));
  INV_X1    g183(.A(G120gat), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT1), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT70), .B(G113gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n383), .B(new_n386), .C1(new_n385), .C2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n384), .B2(new_n385), .ZN(new_n389));
  INV_X1    g188(.A(new_n381), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n298), .A2(new_n393), .A3(KEYINPUT4), .A4(new_n300), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n392), .A3(new_n290), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n397), .B(KEYINPUT79), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n388), .A2(new_n286), .A3(new_n391), .A4(new_n289), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n394), .A2(new_n396), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n392), .A2(new_n294), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n400), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n392), .A2(new_n294), .A3(KEYINPUT81), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n403), .B(KEYINPUT5), .C1(new_n399), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n400), .A2(KEYINPUT4), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n298), .A2(new_n393), .A3(new_n300), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(KEYINPUT4), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n399), .A4(new_n396), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT0), .ZN(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n409), .A2(new_n419), .A3(new_n414), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n419), .B1(new_n409), .B2(new_n414), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT6), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n380), .A2(new_n427), .A3(KEYINPUT35), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT75), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT32), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n361), .A2(new_n393), .ZN(new_n431));
  INV_X1    g230(.A(G227gat), .ZN(new_n432));
  INV_X1    g231(.A(G233gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n353), .A2(new_n392), .A3(new_n360), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT72), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n431), .A2(KEYINPUT72), .A3(new_n434), .A4(new_n435), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n430), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT33), .B1(new_n438), .B2(new_n439), .ZN(new_n441));
  XOR2_X1   g240(.A(G15gat), .B(G43gat), .Z(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n440), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  AOI221_X4 g245(.A(new_n430), .B1(KEYINPUT33), .B2(new_n444), .C1(new_n438), .C2(new_n439), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n429), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n441), .A2(new_n445), .ZN(new_n449));
  INV_X1    g248(.A(new_n440), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n447), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(KEYINPUT75), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n431), .A2(new_n435), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n432), .B2(new_n433), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n457), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n448), .A2(new_n453), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n460), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(new_n429), .C1(new_n446), .C2(new_n447), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(KEYINPUT87), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT87), .B1(new_n461), .B2(new_n463), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n320), .B(new_n428), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n320), .ZN(new_n468));
  OAI22_X1  g267(.A1(KEYINPUT73), .A2(new_n462), .B1(new_n446), .B2(new_n447), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT73), .B1(new_n458), .B2(new_n459), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n452), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n468), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n424), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n421), .A2(KEYINPUT82), .A3(new_n422), .A4(new_n423), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n426), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n476), .A3(new_n379), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT35), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n399), .B1(new_n412), .B2(new_n396), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n398), .B1(new_n406), .B2(new_n407), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n482), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n419), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n425), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n484), .A2(KEYINPUT40), .A3(new_n419), .A4(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n320), .B1(new_n490), .B2(new_n379), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n366), .A2(new_n368), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n373), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n366), .B2(new_n368), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(KEYINPUT85), .A3(new_n373), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT38), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n495), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n424), .A2(new_n426), .A3(new_n376), .ZN(new_n501));
  NOR4_X1   g300(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT85), .A4(KEYINPUT38), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n480), .B1(new_n491), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n498), .A2(new_n499), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n494), .B2(new_n496), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n380), .A2(new_n489), .A3(new_n488), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT86), .A4(new_n320), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n469), .A2(KEYINPUT36), .A3(new_n471), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n461), .A2(new_n463), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n476), .A2(new_n379), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n468), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n511), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n270), .B1(new_n479), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n476), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT9), .ZN(new_n521));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n523), .B2(new_n522), .ZN(new_n525));
  OR2_X1    g324(.A1(G71gat), .A2(G78gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n522), .B(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n527), .B1(new_n526), .B2(new_n521), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT21), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n536), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G127gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n536), .B(new_n537), .ZN(new_n541));
  INV_X1    g340(.A(G127gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n233), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n525), .A2(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(KEYINPUT21), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n547), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n540), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT95), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G155gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT96), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n553), .B(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n548), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n548), .B2(new_n550), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT97), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n564));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G190gat), .B(G218gat), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT100), .B(G92gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n570), .A2(new_n571), .B1(KEYINPUT8), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT98), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(KEYINPUT7), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT99), .B1(new_n577), .B2(KEYINPUT98), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(new_n579), .A3(KEYINPUT7), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n573), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G99gat), .B(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n578), .A2(new_n580), .ZN(new_n588));
  INV_X1    g387(.A(new_n576), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(new_n584), .A3(new_n573), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n586), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n592), .A2(KEYINPUT101), .A3(new_n584), .A4(new_n573), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n249), .B2(new_n248), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n597), .A2(new_n224), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n569), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n599), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n604), .A2(new_n568), .A3(new_n601), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n567), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n600), .A2(new_n569), .A3(new_n602), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n568), .B1(new_n604), .B2(new_n601), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n566), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n534), .A3(new_n595), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n546), .A2(new_n593), .A3(new_n586), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n546), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n614), .ZN(new_n620));
  INV_X1    g419(.A(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n619), .B2(new_n622), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n560), .A2(new_n611), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n519), .A2(new_n520), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g432(.A1(new_n519), .A2(new_n631), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n634), .A2(new_n380), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(new_n227), .B2(new_n635), .ZN(new_n638));
  MUX2_X1   g437(.A(new_n637), .B(new_n638), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g438(.A(G15gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n465), .A2(new_n466), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n519), .A2(new_n640), .A3(new_n642), .A4(new_n631), .ZN(new_n643));
  INV_X1    g442(.A(new_n515), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n645), .B2(new_n640), .ZN(G1326gat));
  NAND2_X1  g445(.A1(new_n634), .A2(new_n468), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT43), .B(G22gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  AND4_X1   g448(.A1(new_n519), .A2(new_n560), .A3(new_n611), .A4(new_n629), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n211), .A3(new_n520), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT45), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n479), .A2(new_n518), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(KEYINPUT44), .A3(new_n611), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n560), .A2(new_n629), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n270), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT102), .B1(new_n516), .B2(new_n468), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n658), .B(new_n320), .C1(new_n476), .C2(new_n379), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n511), .A2(new_n660), .A3(new_n515), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n610), .B1(new_n479), .B2(new_n661), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n654), .B(new_n656), .C1(new_n662), .C2(KEYINPUT44), .ZN(new_n663));
  OAI21_X1  g462(.A(G29gat), .B1(new_n663), .B2(new_n476), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n652), .A2(new_n664), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n212), .A3(new_n380), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT46), .Z(new_n667));
  OAI21_X1  g466(.A(G36gat), .B1(new_n663), .B2(new_n379), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(G1329gat));
  OAI21_X1  g468(.A(G43gat), .B1(new_n663), .B2(new_n515), .ZN(new_n670));
  INV_X1    g469(.A(G43gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n650), .A2(new_n671), .A3(new_n642), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g473(.A(new_n204), .B1(new_n663), .B2(new_n320), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n320), .A2(new_n204), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n650), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT48), .B1(new_n677), .B2(KEYINPUT103), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1331gat));
  NOR2_X1   g479(.A1(new_n560), .A2(new_n611), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n270), .A3(new_n630), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n479), .B2(new_n661), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n476), .B(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g485(.A(new_n379), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT105), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(G1333gat));
  NAND2_X1  g490(.A1(new_n683), .A2(new_n644), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n641), .A2(G71gat), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n692), .A2(G71gat), .B1(new_n683), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g494(.A1(new_n683), .A2(new_n468), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT106), .B(G78gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1335gat));
  NAND2_X1  g497(.A1(new_n560), .A2(new_n270), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(KEYINPUT107), .Z(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n629), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n654), .B(new_n701), .C1(new_n662), .C2(KEYINPUT44), .ZN(new_n702));
  OAI21_X1  g501(.A(G85gat), .B1(new_n702), .B2(new_n476), .ZN(new_n703));
  INV_X1    g502(.A(new_n700), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT87), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n513), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n468), .B1(new_n706), .B2(new_n464), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n707), .A2(new_n428), .B1(KEYINPUT35), .B2(new_n477), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n511), .A2(new_n660), .A3(new_n515), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n611), .B(new_n704), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT51), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n662), .A2(KEYINPUT51), .A3(new_n704), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n520), .A2(new_n571), .A3(new_n630), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n703), .B1(new_n715), .B2(new_n716), .ZN(G1336gat));
  NAND3_X1  g516(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT108), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n710), .A2(new_n719), .A3(new_n711), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n379), .A2(new_n629), .A3(G92gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT109), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n718), .A2(new_n720), .A3(new_n724), .A4(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(new_n570), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n702), .B2(new_n379), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n723), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT52), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT52), .B1(new_n714), .B2(new_n721), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1337gat));
  OAI21_X1  g531(.A(G99gat), .B1(new_n702), .B2(new_n515), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n641), .A2(G99gat), .A3(new_n629), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT110), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n735), .B2(new_n715), .ZN(G1338gat));
  NOR3_X1   g535(.A1(new_n320), .A2(G106gat), .A3(new_n629), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT111), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n718), .A2(new_n720), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT112), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n718), .A2(new_n720), .A3(new_n741), .A4(new_n738), .ZN(new_n742));
  OAI21_X1  g541(.A(G106gat), .B1(new_n702), .B2(new_n320), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT53), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT53), .B1(new_n714), .B2(new_n737), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1339gat));
  NAND3_X1  g547(.A1(new_n615), .A2(new_n621), .A3(new_n616), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n619), .A2(KEYINPUT54), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT113), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n619), .A2(new_n752), .A3(KEYINPUT54), .A4(new_n749), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n621), .B1(new_n615), .B2(new_n616), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n625), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n751), .A2(KEYINPUT55), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(new_n626), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n751), .A2(new_n753), .A3(new_n756), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(KEYINPUT114), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT114), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT115), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n765), .B(new_n758), .C1(new_n761), .C2(new_n762), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n269), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n246), .B1(new_n245), .B2(new_n251), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n256), .A2(new_n257), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n264), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n268), .B(new_n770), .C1(new_n628), .C2(new_n627), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n611), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  AND4_X1   g571(.A1(new_n268), .A2(new_n606), .A3(new_n770), .A4(new_n609), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n764), .A2(new_n773), .A3(new_n766), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n560), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n631), .A2(new_n270), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(new_n707), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n476), .A2(new_n380), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(G113gat), .B1(new_n781), .B2(new_n270), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT116), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n778), .A2(new_n684), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(new_n472), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n379), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT117), .Z(new_n787));
  NAND2_X1  g586(.A1(new_n269), .A2(new_n387), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(G1340gat));
  OAI21_X1  g588(.A(G120gat), .B1(new_n781), .B2(new_n629), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT118), .Z(new_n791));
  NAND2_X1  g590(.A1(new_n630), .A2(new_n385), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n787), .B2(new_n792), .ZN(G1341gat));
  OAI21_X1  g592(.A(G127gat), .B1(new_n781), .B2(new_n560), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n559), .A2(new_n542), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n786), .B2(new_n795), .ZN(G1342gat));
  INV_X1    g595(.A(G134gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n380), .A2(new_n610), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n785), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n799), .A2(KEYINPUT56), .ZN(new_n800));
  OAI21_X1  g599(.A(G134gat), .B1(new_n781), .B2(new_n610), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(KEYINPUT56), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(G1343gat));
  AND2_X1   g602(.A1(new_n515), .A2(new_n780), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n320), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n759), .A2(new_n760), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n269), .A3(new_n626), .A4(new_n757), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n611), .B1(new_n808), .B2(new_n771), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n559), .B1(new_n774), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n631), .A2(new_n270), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n806), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT119), .Z(new_n814));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n778), .B2(new_n468), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n804), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(G141gat), .B1(new_n816), .B2(new_n270), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n644), .A2(new_n320), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n784), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n380), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n270), .A2(G141gat), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n817), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT58), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n817), .B(new_n826), .C1(new_n821), .C2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1344gat));
  OAI211_X1 g627(.A(new_n773), .B(new_n758), .C1(new_n761), .C2(new_n762), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n560), .B1(new_n830), .B2(new_n809), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n320), .B1(new_n831), .B2(new_n777), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT120), .B1(new_n832), .B2(KEYINPUT57), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n834));
  INV_X1    g633(.A(new_n771), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n760), .A2(new_n759), .B1(new_n267), .B2(new_n268), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n758), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n829), .B1(new_n837), .B2(new_n611), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n812), .B1(new_n838), .B2(new_n560), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n834), .B(new_n805), .C1(new_n839), .C2(new_n320), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n778), .A2(new_n806), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n844), .A2(new_n630), .A3(new_n804), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT59), .B1(new_n845), .B2(new_n277), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n277), .A2(KEYINPUT59), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n816), .B2(new_n629), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n820), .A2(new_n277), .A3(new_n630), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1345gat));
  OAI21_X1  g650(.A(new_n282), .B1(new_n816), .B2(new_n560), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n820), .A2(new_n283), .A3(new_n559), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1346gat));
  OAI21_X1  g653(.A(G162gat), .B1(new_n816), .B2(new_n610), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n798), .A2(new_n284), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n819), .B2(new_n856), .ZN(G1347gat));
  NAND2_X1  g656(.A1(new_n778), .A2(new_n476), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT121), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n379), .B1(new_n858), .B2(KEYINPUT121), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n469), .A2(new_n471), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n861), .A2(new_n862), .A3(new_n468), .ZN(new_n863));
  AOI21_X1  g662(.A(G169gat), .B1(new_n863), .B2(new_n269), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n684), .A2(new_n379), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n779), .A2(KEYINPUT122), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT122), .B1(new_n779), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n270), .A2(new_n326), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n864), .B1(new_n868), .B2(new_n869), .ZN(G1348gat));
  NAND3_X1  g669(.A1(new_n863), .A2(new_n327), .A3(new_n630), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n866), .A2(new_n867), .A3(new_n629), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n327), .B2(new_n872), .ZN(G1349gat));
  NOR3_X1   g672(.A1(new_n866), .A2(new_n867), .A3(new_n560), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n331), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n559), .A2(new_n350), .ZN(new_n876));
  NOR4_X1   g675(.A1(new_n861), .A2(new_n862), .A3(new_n468), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT60), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n861), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n879), .A2(new_n350), .A3(new_n472), .A4(new_n559), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n880), .B(new_n881), .C1(new_n874), .C2(new_n331), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n882), .ZN(G1350gat));
  NAND3_X1  g682(.A1(new_n863), .A2(new_n330), .A3(new_n611), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n611), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(G190gat), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n885), .B2(G190gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(G1351gat));
  AND3_X1   g688(.A1(new_n859), .A2(new_n818), .A3(new_n860), .ZN(new_n890));
  AOI21_X1  g689(.A(G197gat), .B1(new_n890), .B2(new_n269), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n844), .B(KEYINPUT123), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n865), .A2(new_n515), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n269), .A2(G197gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(G1352gat));
  NAND4_X1  g696(.A1(new_n892), .A2(KEYINPUT125), .A3(new_n630), .A4(new_n894), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n844), .A2(KEYINPUT123), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n900), .B1(new_n842), .B2(new_n843), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n630), .B(new_n894), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n898), .A2(new_n904), .A3(G204gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n629), .A2(G204gat), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n859), .A2(new_n860), .A3(new_n818), .A4(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT62), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n907), .B2(KEYINPUT62), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n907), .A2(KEYINPUT62), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n905), .A2(new_n911), .A3(new_n912), .ZN(G1353gat));
  NOR2_X1   g712(.A1(new_n560), .A2(G211gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n890), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n893), .A2(new_n560), .ZN(new_n917));
  INV_X1    g716(.A(new_n806), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n776), .B2(new_n777), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n916), .B(new_n917), .C1(new_n919), .C2(new_n841), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n920), .A2(G211gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n919), .B2(new_n841), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT126), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT63), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AND4_X1   g723(.A1(KEYINPUT63), .A2(new_n923), .A3(G211gat), .A4(new_n920), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT127), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n915), .B(new_n928), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1354gat));
  AOI21_X1  g729(.A(G218gat), .B1(new_n890), .B2(new_n611), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n611), .A2(G218gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n895), .B2(new_n932), .ZN(G1355gat));
endmodule


