

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759;

  AND2_X1 U366 ( .A1(n582), .A2(n581), .ZN(n351) );
  NOR2_X1 U367 ( .A1(n701), .A2(n564), .ZN(n682) );
  XNOR2_X1 U368 ( .A(KEYINPUT99), .B(n522), .ZN(n561) );
  AND2_X1 U369 ( .A1(n539), .A2(n704), .ZN(n343) );
  XNOR2_X1 U370 ( .A(n744), .B(G146), .ZN(n495) );
  XNOR2_X1 U371 ( .A(n472), .B(G134), .ZN(n489) );
  XNOR2_X1 U372 ( .A(G119), .B(G110), .ZN(n500) );
  XNOR2_X1 U373 ( .A(KEYINPUT85), .B(G110), .ZN(n424) );
  OR2_X1 U374 ( .A1(n687), .A2(KEYINPUT34), .ZN(n403) );
  AND2_X2 U375 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X2 U376 ( .A(n661), .B(n430), .ZN(n636) );
  XNOR2_X2 U377 ( .A(n387), .B(n494), .ZN(n661) );
  NOR2_X1 U378 ( .A1(n701), .A2(n700), .ZN(n601) );
  XNOR2_X2 U379 ( .A(n344), .B(KEYINPUT0), .ZN(n593) );
  XNOR2_X1 U380 ( .A(n400), .B(n401), .ZN(n505) );
  NAND2_X1 U381 ( .A1(n535), .A2(n343), .ZN(n520) );
  AND2_X2 U382 ( .A1(n399), .A2(n586), .ZN(n733) );
  NAND2_X2 U383 ( .A1(n654), .A2(n414), .ZN(n730) );
  XNOR2_X2 U384 ( .A(G107), .B(G104), .ZN(n423) );
  XNOR2_X2 U385 ( .A(G101), .B(KEYINPUT73), .ZN(n422) );
  XNOR2_X2 U386 ( .A(n495), .B(n389), .ZN(n620) );
  NOR2_X1 U387 ( .A1(n608), .A2(n549), .ZN(n521) );
  INV_X4 U388 ( .A(G953), .ZN(n466) );
  NOR2_X1 U389 ( .A1(n380), .A2(n379), .ZN(n378) );
  NAND2_X1 U390 ( .A1(n724), .A2(KEYINPUT2), .ZN(n380) );
  AND2_X1 U391 ( .A1(n611), .A2(n383), .ZN(n368) );
  XNOR2_X1 U392 ( .A(n351), .B(KEYINPUT48), .ZN(n399) );
  NOR2_X1 U393 ( .A1(n758), .A2(n759), .ZN(n558) );
  NAND2_X1 U394 ( .A1(n416), .A2(n532), .ZN(n415) );
  NOR2_X1 U395 ( .A1(n607), .A2(n609), .ZN(n610) );
  AND2_X1 U396 ( .A1(n583), .A2(n545), .ZN(n548) );
  XNOR2_X1 U397 ( .A(n555), .B(n554), .ZN(n713) );
  XNOR2_X1 U398 ( .A(n398), .B(KEYINPUT74), .ZN(n542) );
  XNOR2_X1 U399 ( .A(n393), .B(n592), .ZN(n687) );
  NAND2_X1 U400 ( .A1(n601), .A2(n590), .ZN(n393) );
  NAND2_X2 U401 ( .A1(n409), .A2(n407), .ZN(n551) );
  XNOR2_X1 U402 ( .A(n531), .B(n492), .ZN(n608) );
  XNOR2_X1 U403 ( .A(n491), .B(n490), .ZN(n531) );
  XNOR2_X1 U404 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U405 ( .A(n489), .B(n488), .ZN(n744) );
  NAND2_X1 U406 ( .A1(n448), .A2(n353), .ZN(n344) );
  XNOR2_X2 U407 ( .A(n559), .B(n360), .ZN(n448) );
  NAND2_X2 U408 ( .A1(n527), .A2(n438), .ZN(n559) );
  XNOR2_X1 U409 ( .A(n423), .B(n422), .ZN(n386) );
  NAND2_X1 U410 ( .A1(n384), .A2(n415), .ZN(n345) );
  NAND2_X1 U411 ( .A1(n384), .A2(n415), .ZN(n588) );
  AND2_X1 U412 ( .A1(n385), .A2(n417), .ZN(n384) );
  BUF_X1 U413 ( .A(n494), .Z(n346) );
  XNOR2_X1 U414 ( .A(n386), .B(n424), .ZN(n494) );
  NAND2_X1 U415 ( .A1(n345), .A2(n587), .ZN(n347) );
  XNOR2_X2 U416 ( .A(n513), .B(n512), .ZN(n587) );
  BUF_X1 U417 ( .A(n559), .Z(n348) );
  BUF_X1 U418 ( .A(n530), .Z(n349) );
  BUF_X1 U419 ( .A(n593), .Z(n602) );
  XNOR2_X1 U420 ( .A(n636), .B(n639), .ZN(n640) );
  NAND2_X1 U421 ( .A1(n365), .A2(n362), .ZN(n616) );
  NAND2_X1 U422 ( .A1(n356), .A2(n363), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n365) );
  NAND2_X1 U424 ( .A1(n477), .A2(n618), .ZN(n374) );
  INV_X1 U425 ( .A(n379), .ZN(n376) );
  AND2_X1 U426 ( .A1(n394), .A2(G210), .ZN(n484) );
  XOR2_X1 U427 ( .A(KEYINPUT5), .B(G101), .Z(n486) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n452) );
  XOR2_X1 U429 ( .A(G122), .B(G104), .Z(n450) );
  XNOR2_X1 U430 ( .A(G140), .B(KEYINPUT10), .ZN(n456) );
  XOR2_X1 U431 ( .A(KEYINPUT4), .B(G131), .Z(n488) );
  INV_X1 U432 ( .A(n523), .ZN(n529) );
  NAND2_X1 U433 ( .A1(n645), .A2(n506), .ZN(n491) );
  XNOR2_X1 U434 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U435 ( .A(G128), .B(KEYINPUT23), .Z(n498) );
  NAND2_X1 U436 ( .A1(n497), .A2(G221), .ZN(n401) );
  AND2_X1 U437 ( .A1(n399), .A2(n359), .ZN(n414) );
  OR2_X1 U438 ( .A1(n620), .A2(n408), .ZN(n407) );
  NAND2_X1 U439 ( .A1(G469), .A2(n506), .ZN(n408) );
  INV_X1 U440 ( .A(KEYINPUT78), .ZN(n366) );
  INV_X1 U441 ( .A(KEYINPUT80), .ZN(n364) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n439) );
  INV_X1 U443 ( .A(G237), .ZN(n431) );
  NAND2_X1 U444 ( .A1(n617), .A2(KEYINPUT64), .ZN(n379) );
  BUF_X1 U445 ( .A(n687), .Z(n698) );
  XNOR2_X1 U446 ( .A(n382), .B(KEYINPUT104), .ZN(n694) );
  NOR2_X1 U447 ( .A1(n690), .A2(n689), .ZN(n382) );
  NAND2_X1 U448 ( .A1(n538), .A2(n539), .ZN(n397) );
  NAND2_X1 U449 ( .A1(n496), .A2(G902), .ZN(n410) );
  XNOR2_X1 U450 ( .A(n495), .B(n395), .ZN(n645) );
  XNOR2_X1 U451 ( .A(n487), .B(n396), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n486), .B(G137), .ZN(n396) );
  BUF_X1 U453 ( .A(n654), .Z(n732) );
  XOR2_X1 U454 ( .A(KEYINPUT9), .B(G122), .Z(n471) );
  XNOR2_X1 U455 ( .A(G116), .B(G107), .ZN(n470) );
  NOR2_X1 U456 ( .A1(G953), .A2(G237), .ZN(n394) );
  XNOR2_X1 U457 ( .A(G113), .B(G143), .ZN(n449) );
  XNOR2_X1 U458 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n427) );
  NAND2_X1 U459 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U460 ( .A1(n570), .A2(n690), .ZN(n544) );
  AND2_X1 U461 ( .A1(n406), .A2(n596), .ZN(n405) );
  AND2_X1 U462 ( .A1(n418), .A2(n533), .ZN(n417) );
  NAND2_X1 U463 ( .A1(n707), .A2(n532), .ZN(n418) );
  XNOR2_X1 U464 ( .A(n465), .B(n464), .ZN(n572) );
  XNOR2_X1 U465 ( .A(n463), .B(KEYINPUT13), .ZN(n464) );
  INV_X1 U466 ( .A(G475), .ZN(n463) );
  XOR2_X1 U467 ( .A(KEYINPUT62), .B(n645), .Z(n646) );
  XNOR2_X1 U468 ( .A(n485), .B(n421), .ZN(n387) );
  XNOR2_X1 U469 ( .A(KEYINPUT16), .B(G122), .ZN(n421) );
  XNOR2_X1 U470 ( .A(n501), .B(n498), .ZN(n400) );
  NAND2_X1 U471 ( .A1(n380), .A2(n357), .ZN(n371) );
  XNOR2_X1 U472 ( .A(n391), .B(n503), .ZN(n390) );
  XNOR2_X1 U473 ( .A(n493), .B(G140), .ZN(n391) );
  NOR2_X1 U474 ( .A1(n466), .A2(G952), .ZN(n648) );
  BUF_X1 U475 ( .A(n612), .Z(n652) );
  BUF_X1 U476 ( .A(n531), .Z(n600) );
  XOR2_X1 U477 ( .A(KEYINPUT76), .B(KEYINPUT8), .Z(n350) );
  XNOR2_X1 U478 ( .A(n350), .B(n467), .ZN(n497) );
  XOR2_X1 U479 ( .A(n625), .B(n624), .Z(n352) );
  XOR2_X1 U480 ( .A(n447), .B(n446), .Z(n353) );
  XOR2_X1 U481 ( .A(n526), .B(n525), .Z(n354) );
  AND2_X1 U482 ( .A1(n606), .A2(n693), .ZN(n355) );
  AND2_X1 U483 ( .A1(n614), .A2(n613), .ZN(n356) );
  AND2_X1 U484 ( .A1(n730), .A2(n618), .ZN(n357) );
  AND2_X1 U485 ( .A1(n608), .A2(n511), .ZN(n358) );
  AND2_X1 U486 ( .A1(n586), .A2(n727), .ZN(n359) );
  XOR2_X1 U487 ( .A(KEYINPUT69), .B(KEYINPUT19), .Z(n360) );
  XNOR2_X1 U488 ( .A(KEYINPUT68), .B(KEYINPUT22), .ZN(n361) );
  XNOR2_X1 U489 ( .A(n347), .B(n364), .ZN(n363) );
  NAND2_X1 U490 ( .A1(n368), .A2(n369), .ZN(n367) );
  XNOR2_X1 U491 ( .A(n589), .B(n370), .ZN(n369) );
  INV_X1 U492 ( .A(KEYINPUT65), .ZN(n370) );
  NAND2_X2 U493 ( .A1(n372), .A2(n371), .ZN(n644) );
  NOR2_X2 U494 ( .A1(n378), .A2(n373), .ZN(n372) );
  NAND2_X1 U495 ( .A1(n375), .A2(n374), .ZN(n373) );
  NAND2_X1 U496 ( .A1(n377), .A2(n376), .ZN(n375) );
  INV_X1 U497 ( .A(n730), .ZN(n377) );
  INV_X1 U498 ( .A(n607), .ZN(n420) );
  NAND2_X1 U499 ( .A1(n530), .A2(n529), .ZN(n607) );
  NOR2_X1 U500 ( .A1(n756), .A2(n355), .ZN(n383) );
  NAND2_X1 U501 ( .A1(n381), .A2(n687), .ZN(n402) );
  NAND2_X1 U502 ( .A1(n388), .A2(n594), .ZN(n381) );
  NAND2_X1 U503 ( .A1(n404), .A2(n405), .ZN(n597) );
  NAND2_X1 U504 ( .A1(n588), .A2(n587), .ZN(n615) );
  NAND2_X1 U505 ( .A1(n420), .A2(n419), .ZN(n385) );
  XNOR2_X2 U506 ( .A(n413), .B(n412), .ZN(n485) );
  NAND2_X1 U507 ( .A1(n349), .A2(n358), .ZN(n513) );
  XNOR2_X1 U508 ( .A(n483), .B(n361), .ZN(n530) );
  INV_X1 U509 ( .A(n602), .ZN(n388) );
  NAND2_X1 U510 ( .A1(n388), .A2(n605), .ZN(n666) );
  XNOR2_X1 U511 ( .A(n346), .B(n390), .ZN(n389) );
  XNOR2_X2 U512 ( .A(n551), .B(KEYINPUT1), .ZN(n701) );
  NAND2_X1 U513 ( .A1(n394), .A2(G214), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n700), .A2(n397), .ZN(n398) );
  OR2_X1 U515 ( .A1(n700), .A2(n551), .ZN(n604) );
  NOR2_X2 U516 ( .A1(n593), .A2(n482), .ZN(n483) );
  XNOR2_X2 U517 ( .A(G143), .B(G128), .ZN(n472) );
  NAND2_X1 U518 ( .A1(n402), .A2(n403), .ZN(n404) );
  NAND2_X1 U519 ( .A1(n602), .A2(KEYINPUT34), .ZN(n406) );
  NAND2_X1 U520 ( .A1(n620), .A2(n496), .ZN(n411) );
  XNOR2_X2 U521 ( .A(G119), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X2 U522 ( .A(G116), .B(G113), .ZN(n413) );
  XNOR2_X2 U523 ( .A(n434), .B(n433), .ZN(n527) );
  NAND2_X1 U524 ( .A1(n654), .A2(n733), .ZN(n724) );
  XNOR2_X2 U525 ( .A(n616), .B(KEYINPUT45), .ZN(n654) );
  INV_X1 U526 ( .A(n420), .ZN(n416) );
  AND2_X1 U527 ( .A1(n600), .A2(KEYINPUT67), .ZN(n419) );
  INV_X1 U528 ( .A(n757), .ZN(n579) );
  AND2_X1 U529 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U530 ( .A(KEYINPUT24), .ZN(n499) );
  INV_X1 U531 ( .A(n502), .ZN(n457) );
  INV_X1 U532 ( .A(KEYINPUT34), .ZN(n594) );
  INV_X1 U533 ( .A(n703), .ZN(n533) );
  NAND2_X1 U534 ( .A1(n466), .A2(G224), .ZN(n425) );
  XNOR2_X1 U535 ( .A(n425), .B(KEYINPUT4), .ZN(n426) );
  XNOR2_X1 U536 ( .A(n472), .B(n426), .ZN(n429) );
  XNOR2_X2 U537 ( .A(G146), .B(G125), .ZN(n455) );
  XNOR2_X1 U538 ( .A(n455), .B(n427), .ZN(n428) );
  XNOR2_X1 U539 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U540 ( .A(KEYINPUT15), .B(G902), .ZN(n477) );
  INV_X1 U541 ( .A(n477), .ZN(n617) );
  OR2_X2 U542 ( .A1(n636), .A2(n617), .ZN(n434) );
  INV_X1 U543 ( .A(G902), .ZN(n506) );
  NAND2_X1 U544 ( .A1(n506), .A2(n431), .ZN(n435) );
  NAND2_X1 U545 ( .A1(n435), .A2(G210), .ZN(n432) );
  XNOR2_X1 U546 ( .A(n432), .B(KEYINPUT75), .ZN(n433) );
  NAND2_X1 U547 ( .A1(n435), .A2(G214), .ZN(n437) );
  INV_X1 U548 ( .A(KEYINPUT86), .ZN(n436) );
  XNOR2_X1 U549 ( .A(n437), .B(n436), .ZN(n689) );
  INV_X1 U550 ( .A(n689), .ZN(n438) );
  XOR2_X1 U551 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n440) );
  XNOR2_X1 U552 ( .A(n440), .B(n439), .ZN(n443) );
  NAND2_X1 U553 ( .A1(G902), .A2(n443), .ZN(n515) );
  INV_X1 U554 ( .A(n515), .ZN(n441) );
  NOR2_X1 U555 ( .A1(G898), .A2(n466), .ZN(n662) );
  NAND2_X1 U556 ( .A1(n441), .A2(n662), .ZN(n442) );
  XOR2_X1 U557 ( .A(KEYINPUT89), .B(n442), .Z(n445) );
  NAND2_X1 U558 ( .A1(n443), .A2(G952), .ZN(n444) );
  XOR2_X1 U559 ( .A(KEYINPUT88), .B(n444), .Z(n718) );
  NAND2_X1 U560 ( .A1(n466), .A2(n718), .ZN(n517) );
  NAND2_X1 U561 ( .A1(n445), .A2(n517), .ZN(n447) );
  INV_X1 U562 ( .A(KEYINPUT90), .ZN(n446) );
  XNOR2_X1 U563 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U564 ( .A(G131), .B(KEYINPUT93), .ZN(n451) );
  XNOR2_X1 U565 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U566 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n456), .B(n455), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n458), .B(n457), .ZN(n462) );
  XOR2_X1 U569 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n460) );
  XNOR2_X1 U570 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U571 ( .A(n462), .B(n461), .ZN(n631) );
  NOR2_X1 U572 ( .A1(G902), .A2(n631), .ZN(n465) );
  XOR2_X1 U573 ( .A(KEYINPUT95), .B(KEYINPUT7), .Z(n469) );
  NAND2_X1 U574 ( .A1(G234), .A2(n466), .ZN(n467) );
  NAND2_X1 U575 ( .A1(G217), .A2(n497), .ZN(n468) );
  XNOR2_X1 U576 ( .A(n469), .B(n468), .ZN(n475) );
  XNOR2_X1 U577 ( .A(n471), .B(n470), .ZN(n473) );
  XNOR2_X1 U578 ( .A(n473), .B(n489), .ZN(n474) );
  XNOR2_X1 U579 ( .A(n475), .B(n474), .ZN(n625) );
  NAND2_X1 U580 ( .A1(n625), .A2(n506), .ZN(n476) );
  XNOR2_X1 U581 ( .A(n476), .B(G478), .ZN(n566) );
  INV_X1 U582 ( .A(n566), .ZN(n571) );
  AND2_X1 U583 ( .A1(n572), .A2(n571), .ZN(n691) );
  NAND2_X1 U584 ( .A1(G234), .A2(n477), .ZN(n478) );
  XNOR2_X1 U585 ( .A(KEYINPUT20), .B(n478), .ZN(n507) );
  NAND2_X1 U586 ( .A1(n507), .A2(G221), .ZN(n480) );
  INV_X1 U587 ( .A(KEYINPUT21), .ZN(n479) );
  XNOR2_X1 U588 ( .A(n480), .B(n479), .ZN(n704) );
  XNOR2_X1 U589 ( .A(n704), .B(KEYINPUT91), .ZN(n534) );
  INV_X1 U590 ( .A(n534), .ZN(n481) );
  NAND2_X1 U591 ( .A1(n691), .A2(n481), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n485), .B(n484), .ZN(n487) );
  INV_X1 U593 ( .A(G472), .ZN(n490) );
  INV_X1 U594 ( .A(KEYINPUT6), .ZN(n492) );
  NAND2_X1 U595 ( .A1(G227), .A2(n466), .ZN(n493) );
  XOR2_X1 U596 ( .A(G137), .B(KEYINPUT71), .Z(n503) );
  INV_X1 U597 ( .A(G469), .ZN(n496) );
  INV_X1 U598 ( .A(n701), .ZN(n523) );
  XNOR2_X1 U599 ( .A(n503), .B(n502), .ZN(n743) );
  INV_X1 U600 ( .A(n743), .ZN(n504) );
  XNOR2_X1 U601 ( .A(n505), .B(n504), .ZN(n626) );
  NAND2_X1 U602 ( .A1(n626), .A2(n506), .ZN(n510) );
  NAND2_X1 U603 ( .A1(n507), .A2(G217), .ZN(n508) );
  XNOR2_X1 U604 ( .A(n508), .B(KEYINPUT25), .ZN(n509) );
  XNOR2_X2 U605 ( .A(n510), .B(n509), .ZN(n535) );
  INV_X1 U606 ( .A(n535), .ZN(n703) );
  NOR2_X1 U607 ( .A1(n529), .A2(n703), .ZN(n511) );
  XNOR2_X1 U608 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n512) );
  XNOR2_X1 U609 ( .A(n587), .B(G119), .ZN(G21) );
  XOR2_X1 U610 ( .A(KEYINPUT100), .B(KEYINPUT43), .Z(n526) );
  INV_X1 U611 ( .A(n572), .ZN(n514) );
  NAND2_X1 U612 ( .A1(n514), .A2(n571), .ZN(n677) );
  INV_X1 U613 ( .A(n677), .ZN(n545) );
  NOR2_X1 U614 ( .A1(G900), .A2(n515), .ZN(n516) );
  NAND2_X1 U615 ( .A1(G953), .A2(n516), .ZN(n518) );
  NAND2_X1 U616 ( .A1(n518), .A2(n517), .ZN(n539) );
  XNOR2_X1 U617 ( .A(n520), .B(KEYINPUT72), .ZN(n549) );
  NAND2_X1 U618 ( .A1(n545), .A2(n521), .ZN(n522) );
  NOR2_X1 U619 ( .A1(n689), .A2(n523), .ZN(n524) );
  NAND2_X1 U620 ( .A1(n561), .A2(n524), .ZN(n525) );
  BUF_X1 U621 ( .A(n527), .Z(n528) );
  INV_X1 U622 ( .A(n528), .ZN(n575) );
  NAND2_X1 U623 ( .A1(n354), .A2(n575), .ZN(n585) );
  XNOR2_X1 U624 ( .A(n585), .B(G140), .ZN(G42) );
  INV_X1 U625 ( .A(KEYINPUT67), .ZN(n532) );
  XNOR2_X1 U626 ( .A(n345), .B(G110), .ZN(G12) );
  NOR2_X1 U627 ( .A1(n535), .A2(n534), .ZN(n537) );
  INV_X1 U628 ( .A(KEYINPUT70), .ZN(n536) );
  XNOR2_X1 U629 ( .A(n537), .B(n536), .ZN(n700) );
  INV_X1 U630 ( .A(n551), .ZN(n538) );
  NOR2_X1 U631 ( .A1(n689), .A2(n600), .ZN(n540) );
  XNOR2_X1 U632 ( .A(KEYINPUT30), .B(n540), .ZN(n541) );
  NAND2_X1 U633 ( .A1(n542), .A2(n541), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n528), .B(KEYINPUT38), .ZN(n690) );
  INV_X1 U635 ( .A(KEYINPUT39), .ZN(n543) );
  XNOR2_X1 U636 ( .A(n544), .B(n543), .ZN(n583) );
  XOR2_X1 U637 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n546) );
  XNOR2_X1 U638 ( .A(KEYINPUT102), .B(n546), .ZN(n547) );
  XNOR2_X1 U639 ( .A(n548), .B(n547), .ZN(n758) );
  XNOR2_X1 U640 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n557) );
  NOR2_X1 U641 ( .A1(n549), .A2(n600), .ZN(n550) );
  XOR2_X1 U642 ( .A(KEYINPUT28), .B(n550), .Z(n552) );
  NOR2_X1 U643 ( .A1(n552), .A2(n551), .ZN(n565) );
  NAND2_X1 U644 ( .A1(n694), .A2(n691), .ZN(n555) );
  XOR2_X1 U645 ( .A(KEYINPUT41), .B(KEYINPUT105), .Z(n553) );
  XNOR2_X1 U646 ( .A(KEYINPUT106), .B(n553), .ZN(n554) );
  NAND2_X1 U647 ( .A1(n565), .A2(n713), .ZN(n556) );
  XNOR2_X1 U648 ( .A(n557), .B(n556), .ZN(n759) );
  XNOR2_X1 U649 ( .A(n558), .B(KEYINPUT46), .ZN(n582) );
  INV_X1 U650 ( .A(n348), .ZN(n560) );
  NAND2_X1 U651 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U652 ( .A(n562), .B(KEYINPUT36), .ZN(n563) );
  XOR2_X1 U653 ( .A(KEYINPUT81), .B(n563), .Z(n564) );
  NAND2_X1 U654 ( .A1(n565), .A2(n448), .ZN(n675) );
  NAND2_X1 U655 ( .A1(n572), .A2(n566), .ZN(n680) );
  NAND2_X1 U656 ( .A1(n677), .A2(n680), .ZN(n693) );
  INV_X1 U657 ( .A(n693), .ZN(n567) );
  NOR2_X1 U658 ( .A1(n675), .A2(n567), .ZN(n568) );
  XOR2_X1 U659 ( .A(KEYINPUT47), .B(n568), .Z(n569) );
  NOR2_X1 U660 ( .A1(n682), .A2(n569), .ZN(n580) );
  INV_X1 U661 ( .A(n570), .ZN(n577) );
  NOR2_X1 U662 ( .A1(n572), .A2(n571), .ZN(n574) );
  INV_X1 U663 ( .A(KEYINPUT98), .ZN(n573) );
  XNOR2_X1 U664 ( .A(n574), .B(n573), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n595), .A2(n575), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U667 ( .A(n578), .B(KEYINPUT101), .ZN(n757) );
  INV_X1 U668 ( .A(n680), .ZN(n584) );
  NAND2_X1 U669 ( .A1(n583), .A2(n584), .ZN(n686) );
  AND2_X1 U670 ( .A1(n585), .A2(n686), .ZN(n586) );
  NAND2_X1 U671 ( .A1(n615), .A2(KEYINPUT44), .ZN(n589) );
  INV_X1 U672 ( .A(n608), .ZN(n590) );
  INV_X1 U673 ( .A(KEYINPUT97), .ZN(n591) );
  XNOR2_X1 U674 ( .A(n591), .B(KEYINPUT33), .ZN(n592) );
  INV_X1 U675 ( .A(n595), .ZN(n596) );
  XNOR2_X2 U676 ( .A(n597), .B(KEYINPUT35), .ZN(n612) );
  NAND2_X1 U677 ( .A1(n612), .A2(KEYINPUT44), .ZN(n599) );
  INV_X1 U678 ( .A(KEYINPUT79), .ZN(n598) );
  XNOR2_X1 U679 ( .A(n599), .B(n598), .ZN(n611) );
  INV_X1 U680 ( .A(n600), .ZN(n707) );
  NAND2_X1 U681 ( .A1(n601), .A2(n707), .ZN(n710) );
  NOR2_X1 U682 ( .A1(n710), .A2(n602), .ZN(n603) );
  XNOR2_X1 U683 ( .A(n603), .B(KEYINPUT31), .ZN(n679) );
  NOR2_X1 U684 ( .A1(n604), .A2(n707), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n679), .A2(n666), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n608), .A2(n703), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT96), .ZN(n756) );
  INV_X1 U688 ( .A(n652), .ZN(n614) );
  INV_X1 U689 ( .A(KEYINPUT44), .ZN(n613) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n727) );
  INV_X1 U691 ( .A(KEYINPUT64), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n644), .A2(G469), .ZN(n622) );
  XOR2_X1 U693 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n619) );
  XNOR2_X1 U694 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n623), .A2(n648), .ZN(G54) );
  NAND2_X1 U697 ( .A1(n644), .A2(G478), .ZN(n624) );
  NOR2_X1 U698 ( .A1(n352), .A2(n648), .ZN(G63) );
  NAND2_X1 U699 ( .A1(n644), .A2(G217), .ZN(n628) );
  XOR2_X1 U700 ( .A(KEYINPUT120), .B(n626), .Z(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n629), .A2(n648), .ZN(G66) );
  NAND2_X1 U703 ( .A1(n644), .A2(G475), .ZN(n633) );
  XOR2_X1 U704 ( .A(KEYINPUT84), .B(KEYINPUT59), .Z(n630) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(n634) );
  NOR2_X2 U706 ( .A1(n634), .A2(n648), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n635), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U708 ( .A1(n644), .A2(G210), .ZN(n641) );
  XOR2_X1 U709 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n638) );
  XNOR2_X1 U710 ( .A(KEYINPUT55), .B(KEYINPUT83), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X2 U713 ( .A1(n642), .A2(n648), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U715 ( .A1(n644), .A2(G472), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n649) );
  NOR2_X2 U717 ( .A1(n649), .A2(n648), .ZN(n651) );
  XOR2_X1 U718 ( .A(KEYINPUT82), .B(KEYINPUT63), .Z(n650) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(G57) );
  XNOR2_X1 U720 ( .A(G122), .B(KEYINPUT126), .ZN(n653) );
  XOR2_X1 U721 ( .A(n653), .B(n652), .Z(G24) );
  NAND2_X1 U722 ( .A1(n732), .A2(n466), .ZN(n655) );
  XOR2_X1 U723 ( .A(KEYINPUT121), .B(n655), .Z(n659) );
  NAND2_X1 U724 ( .A1(G953), .A2(G224), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT61), .B(n656), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n657), .A2(G898), .ZN(n658) );
  NAND2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT122), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n661), .A2(n662), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n664), .B(n663), .ZN(G69) );
  NOR2_X1 U731 ( .A1(n677), .A2(n666), .ZN(n665) );
  XOR2_X1 U732 ( .A(G104), .B(n665), .Z(G6) );
  NOR2_X1 U733 ( .A1(n666), .A2(n680), .ZN(n670) );
  XOR2_X1 U734 ( .A(KEYINPUT109), .B(KEYINPUT26), .Z(n668) );
  XNOR2_X1 U735 ( .A(G107), .B(KEYINPUT27), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(G9) );
  NOR2_X1 U738 ( .A1(n675), .A2(n680), .ZN(n674) );
  XOR2_X1 U739 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n672) );
  XNOR2_X1 U740 ( .A(G128), .B(KEYINPUT29), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n674), .B(n673), .ZN(G30) );
  NOR2_X1 U743 ( .A1(n675), .A2(n677), .ZN(n676) );
  XOR2_X1 U744 ( .A(G146), .B(n676), .Z(G48) );
  NOR2_X1 U745 ( .A1(n677), .A2(n679), .ZN(n678) );
  XOR2_X1 U746 ( .A(G113), .B(n678), .Z(G15) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U748 ( .A(G116), .B(n681), .Z(G18) );
  XNOR2_X1 U749 ( .A(n682), .B(KEYINPUT112), .ZN(n683) );
  XNOR2_X1 U750 ( .A(n683), .B(KEYINPUT37), .ZN(n684) );
  XNOR2_X1 U751 ( .A(G125), .B(n684), .ZN(G27) );
  XOR2_X1 U752 ( .A(G134), .B(KEYINPUT113), .Z(n685) );
  XNOR2_X1 U753 ( .A(n686), .B(n685), .ZN(G36) );
  NAND2_X1 U754 ( .A1(n698), .A2(n713), .ZN(n688) );
  XNOR2_X1 U755 ( .A(KEYINPUT116), .B(n688), .ZN(n722) );
  NAND2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U760 ( .A(KEYINPUT114), .B(n697), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n716) );
  NAND2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U763 ( .A(n702), .B(KEYINPUT50), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U765 ( .A(KEYINPUT49), .B(n705), .Z(n706) );
  NOR2_X1 U766 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U767 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U768 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U769 ( .A(KEYINPUT51), .B(n712), .Z(n714) );
  NAND2_X1 U770 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U771 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U772 ( .A(n717), .B(KEYINPUT52), .ZN(n719) );
  NAND2_X1 U773 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U774 ( .A(KEYINPUT115), .B(n720), .Z(n721) );
  NAND2_X1 U775 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U776 ( .A(n723), .B(KEYINPUT117), .ZN(n739) );
  INV_X1 U777 ( .A(KEYINPUT77), .ZN(n726) );
  NAND2_X1 U778 ( .A1(n724), .A2(n726), .ZN(n725) );
  NAND2_X1 U779 ( .A1(n725), .A2(KEYINPUT2), .ZN(n729) );
  NAND2_X1 U780 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U781 ( .A1(n731), .A2(n730), .ZN(n737) );
  INV_X1 U782 ( .A(n732), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(KEYINPUT77), .ZN(n736) );
  NAND2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U787 ( .A(KEYINPUT118), .B(n740), .ZN(n741) );
  NOR2_X1 U788 ( .A1(n741), .A2(G953), .ZN(n742) );
  XNOR2_X1 U789 ( .A(n742), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U790 ( .A(n744), .B(n743), .ZN(n748) );
  INV_X1 U791 ( .A(n733), .ZN(n745) );
  XOR2_X1 U792 ( .A(n748), .B(n745), .Z(n746) );
  NOR2_X1 U793 ( .A1(G953), .A2(n746), .ZN(n747) );
  XNOR2_X1 U794 ( .A(n747), .B(KEYINPUT123), .ZN(n754) );
  XNOR2_X1 U795 ( .A(n748), .B(G227), .ZN(n749) );
  XNOR2_X1 U796 ( .A(n749), .B(KEYINPUT124), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n750), .A2(G900), .ZN(n751) );
  XOR2_X1 U798 ( .A(KEYINPUT125), .B(n751), .Z(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(G953), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n754), .A2(n753), .ZN(G72) );
  XOR2_X1 U801 ( .A(G101), .B(KEYINPUT108), .Z(n755) );
  XNOR2_X1 U802 ( .A(n756), .B(n755), .ZN(G3) );
  XOR2_X1 U803 ( .A(G143), .B(n757), .Z(G45) );
  XOR2_X1 U804 ( .A(G131), .B(n758), .Z(G33) );
  XOR2_X1 U805 ( .A(G137), .B(n759), .Z(G39) );
endmodule

