//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1130;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n458), .A2(new_n460), .A3(G137), .ZN(new_n461));
  NAND2_X1  g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n458), .A2(new_n460), .A3(G125), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n458), .A2(new_n460), .A3(KEYINPUT67), .A4(G125), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n469), .B2(G2105), .ZN(G160));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n474), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n457), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G102), .ZN(new_n485));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n471), .B2(G126), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n485), .B1(new_n488), .B2(new_n475), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n458), .A2(new_n460), .A3(G138), .A4(new_n475), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n471), .A2(KEYINPUT4), .A3(G138), .A4(new_n475), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n483), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n485), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n458), .A2(new_n460), .A3(G126), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n486), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n499), .A2(KEYINPUT68), .A3(new_n492), .A4(new_n493), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT70), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n512), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(KEYINPUT69), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(KEYINPUT69), .ZN(new_n527));
  OAI221_X1 g102(.A(new_n521), .B1(new_n522), .B2(new_n510), .C1(new_n526), .C2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n510), .A2(new_n530), .B1(new_n512), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n516), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G171));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT71), .B(G43), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n510), .A2(new_n536), .B1(new_n512), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n516), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  INV_X1    g122(.A(G78), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT72), .B1(new_n548), .B2(new_n502), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n550), .A2(G78), .A3(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n503), .A2(new_n505), .A3(G65), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(G651), .A3(new_n557), .ZN(new_n558));
  OAI211_X1 g133(.A(G53), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(new_n510), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G91), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n558), .A2(new_n560), .A3(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n561), .A2(G87), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n503), .A2(new_n505), .ZN(new_n571));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT74), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n576), .A3(G651), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n575), .A2(new_n577), .B1(G86), .B2(new_n561), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT75), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(new_n561), .A2(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI221_X1 g159(.A(new_n582), .B1(new_n583), .B2(new_n512), .C1(new_n516), .C2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n512), .B(KEYINPUT76), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G54), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n506), .A2(new_n509), .A3(G92), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n506), .A2(G66), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT77), .Z(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n588), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n586), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n586), .B1(new_n595), .B2(G868), .ZN(G321));
  MUX2_X1   g172(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g173(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n595), .B1(new_n600), .B2(G860), .ZN(G148));
  NOR2_X1   g176(.A1(new_n541), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n600), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n471), .A2(new_n484), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n473), .A2(G123), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n477), .A2(G135), .ZN(new_n612));
  NOR2_X1   g187(.A1(G99), .A2(G2105), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2096), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n610), .A2(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(G2451), .B(G2454), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT16), .ZN(new_n619));
  XOR2_X1   g194(.A(G2443), .B(G2446), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G1341), .B(G1348), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT15), .B(G2435), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n623), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G14), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(G401));
  XOR2_X1   g206(.A(G2084), .B(G2090), .Z(new_n632));
  XOR2_X1   g207(.A(G2072), .B(G2078), .Z(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n633), .B(new_n634), .Z(new_n635));
  XOR2_X1   g210(.A(G2067), .B(G2678), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n632), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n633), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n638), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n635), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n641), .A2(new_n636), .A3(new_n632), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n637), .A2(new_n639), .A3(new_n632), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT79), .B(KEYINPUT18), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n640), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2096), .B(G2100), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G227));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n650));
  XOR2_X1   g225(.A(G1956), .B(G2474), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT81), .ZN(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT82), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n650), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n652), .A2(new_n654), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n655), .A3(new_n657), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n655), .A2(new_n650), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(new_n659), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n658), .B(new_n661), .C1(new_n663), .C2(new_n657), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1981), .B(G1991), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G1996), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT83), .B(G1986), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n664), .B(new_n670), .ZN(G229));
  NAND2_X1  g246(.A1(new_n473), .A2(G119), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n477), .A2(G131), .ZN(new_n673));
  NOR2_X1   g248(.A1(G95), .A2(G2105), .ZN(new_n674));
  OAI21_X1  g249(.A(G2104), .B1(new_n475), .B2(G107), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n672), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  MUX2_X1   g251(.A(G25), .B(new_n676), .S(G29), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT35), .B(G1991), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(G1986), .ZN(new_n680));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n681), .A2(G24), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(G290), .B2(G16), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n679), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(G23), .ZN(new_n685));
  INV_X1    g260(.A(G288), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n681), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT33), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1976), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n681), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n681), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT85), .B(G1971), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G6), .B(G305), .S(G16), .Z(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT32), .B(G1981), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT84), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n689), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n684), .B1(new_n698), .B2(KEYINPUT34), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(KEYINPUT34), .B2(new_n698), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n680), .B2(new_n683), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT36), .Z(new_n702));
  NOR2_X1   g277(.A1(G27), .A2(G29), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G164), .B2(G29), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT92), .B(G2078), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G33), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(new_n475), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n484), .A2(G103), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT88), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT25), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n710), .B(new_n713), .C1(G139), .C2(new_n477), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n708), .B1(new_n714), .B2(new_n707), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2072), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT31), .B(G11), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n615), .A2(new_n707), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT91), .B(G28), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT30), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(G29), .ZN(new_n721));
  NOR2_X1   g296(.A1(G5), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G171), .B2(G16), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n718), .B(new_n721), .C1(new_n723), .C2(G1961), .ZN(new_n724));
  OR2_X1    g299(.A1(G29), .A2(G32), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n477), .A2(G141), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n473), .A2(G129), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n484), .A2(G105), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n707), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n724), .B1(G1961), .B2(new_n723), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n681), .A2(G19), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n541), .B2(new_n681), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G1341), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(new_n734), .ZN(new_n739));
  NAND2_X1  g314(.A1(G168), .A2(G16), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G16), .B2(G21), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n738), .B(new_n739), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NOR4_X1   g318(.A1(new_n716), .A2(new_n717), .A3(new_n735), .A4(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G1341), .B2(new_n737), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n595), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G4), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1348), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  NAND2_X1  g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n750), .A2(new_n707), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G160), .B2(new_n707), .ZN(new_n753));
  OAI22_X1  g328(.A1(new_n747), .A2(new_n748), .B1(G2084), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(G299), .A2(G16), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(KEYINPUT23), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n681), .A2(G20), .ZN(new_n757));
  MUX2_X1   g332(.A(KEYINPUT23), .B(new_n756), .S(new_n757), .Z(new_n758));
  AOI211_X1 g333(.A(new_n749), .B(new_n754), .C1(G1956), .C2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(G1956), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n741), .A2(new_n742), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n753), .A2(G2084), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT89), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n473), .A2(G128), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n477), .A2(G140), .ZN(new_n766));
  NOR2_X1   g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(new_n475), .B2(G116), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT86), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n707), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT87), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n707), .A2(G35), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G162), .B2(new_n707), .ZN(new_n778));
  MUX2_X1   g353(.A(new_n777), .B(new_n778), .S(KEYINPUT93), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2090), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n745), .A2(new_n764), .A3(new_n776), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n702), .A2(new_n706), .A3(new_n782), .ZN(G150));
  INV_X1    g358(.A(G150), .ZN(G311));
  INV_X1    g359(.A(G93), .ZN(new_n785));
  INV_X1    g360(.A(G55), .ZN(new_n786));
  OAI22_X1  g361(.A1(new_n510), .A2(new_n785), .B1(new_n512), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n506), .A2(G67), .ZN(new_n788));
  NAND2_X1  g363(.A1(G80), .A2(G543), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n516), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G860), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT37), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n595), .A2(G559), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n541), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n797), .B2(new_n791), .ZN(new_n799));
  INV_X1    g374(.A(new_n791), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n800), .A2(KEYINPUT94), .A3(new_n541), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n796), .B(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n793), .B1(new_n803), .B2(G860), .ZN(G145));
  AOI22_X1  g379(.A1(G130), .A2(new_n473), .B1(new_n477), .B2(G142), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n475), .A2(G118), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n457), .B1(new_n806), .B2(KEYINPUT95), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n807), .B1(KEYINPUT95), .B2(new_n806), .C1(G106), .C2(G2105), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(new_n676), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT96), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(new_n608), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n489), .A2(new_n494), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n769), .B(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(new_n732), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(new_n714), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n615), .B(G160), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(new_n481), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n812), .A2(new_n816), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n823), .A2(new_n818), .A3(new_n817), .ZN(new_n824));
  AOI21_X1  g399(.A(G37), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n823), .A2(new_n817), .A3(new_n821), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g403(.A(new_n802), .B(new_n603), .Z(new_n829));
  OR2_X1    g404(.A1(new_n595), .A2(G299), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n595), .A2(G299), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(new_n835), .A3(new_n831), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n595), .A2(new_n835), .A3(G299), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n838), .A2(KEYINPUT41), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n834), .B1(new_n840), .B2(new_n829), .ZN(new_n841));
  XNOR2_X1  g416(.A(G166), .B(KEYINPUT100), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n686), .ZN(new_n843));
  XOR2_X1   g418(.A(G305), .B(G290), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT42), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n841), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G868), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G868), .B2(new_n800), .ZN(new_n849));
  MUX2_X1   g424(.A(new_n848), .B(new_n849), .S(KEYINPUT101), .Z(G295));
  MUX2_X1   g425(.A(new_n848), .B(new_n849), .S(KEYINPUT101), .Z(G331));
  INV_X1    g426(.A(KEYINPUT44), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(G301), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(G286), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n802), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n799), .A2(new_n855), .A3(new_n801), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(G301), .A2(new_n853), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n833), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n860), .B1(new_n857), .B2(new_n858), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n864), .B1(new_n867), .B2(new_n840), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n868), .B2(new_n845), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n870));
  INV_X1    g445(.A(new_n845), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(new_n864), .C1(new_n867), .C2(new_n840), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT103), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n869), .A2(new_n875), .A3(new_n870), .A4(new_n872), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n852), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n832), .B1(new_n867), .B2(new_n839), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n838), .B(KEYINPUT41), .C1(new_n865), .C2(new_n866), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n869), .B1(new_n880), .B2(new_n845), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT43), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n877), .A2(KEYINPUT104), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT104), .B1(new_n877), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n881), .A2(KEYINPUT43), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n870), .B1(new_n869), .B2(new_n872), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI22_X1  g462(.A1(new_n883), .A2(new_n884), .B1(KEYINPUT44), .B2(new_n887), .ZN(G397));
  INV_X1    g463(.A(KEYINPUT123), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT53), .ZN(new_n890));
  INV_X1    g465(.A(G1384), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n495), .A2(new_n500), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT45), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G40), .ZN(new_n895));
  AOI211_X1 g470(.A(new_n895), .B(new_n463), .C1(new_n469), .C2(G2105), .ZN(new_n896));
  OAI211_X1 g471(.A(KEYINPUT45), .B(new_n891), .C1(new_n489), .C2(new_n494), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n890), .B1(new_n899), .B2(G2078), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n469), .A2(G2105), .ZN(new_n901));
  INV_X1    g476(.A(new_n463), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(G40), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(new_n892), .B2(KEYINPUT50), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n891), .B1(new_n489), .B2(new_n494), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n905), .A2(KEYINPUT50), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  XOR2_X1   g483(.A(KEYINPUT121), .B(G1961), .Z(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND4_X1   g485(.A1(KEYINPUT45), .A2(new_n495), .A3(new_n500), .A4(new_n891), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n905), .A2(new_n893), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n896), .ZN(new_n913));
  NOR4_X1   g488(.A1(new_n911), .A2(new_n913), .A3(new_n890), .A4(G2078), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT122), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n910), .A2(KEYINPUT122), .A3(new_n914), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n900), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(G171), .B(KEYINPUT54), .Z(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1976), .ZN(new_n922));
  OAI221_X1 g497(.A(G8), .B1(G288), .B2(new_n922), .C1(new_n903), .C2(new_n905), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT52), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n903), .A2(new_n905), .ZN(new_n927));
  INV_X1    g502(.A(G8), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n686), .A2(G1976), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n929), .A2(KEYINPUT107), .A3(KEYINPUT52), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(G288), .A2(new_n925), .A3(new_n922), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n926), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n934));
  INV_X1    g509(.A(G1981), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n578), .A2(new_n935), .A3(new_n580), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n935), .B1(new_n578), .B2(new_n580), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n938), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(KEYINPUT49), .A3(new_n936), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n941), .A3(new_n929), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n933), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1971), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n899), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G2090), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n904), .A2(new_n946), .A3(new_n906), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n928), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT55), .ZN(new_n949));
  NAND3_X1  g524(.A1(G303), .A2(new_n949), .A3(G8), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT55), .B1(G166), .B2(new_n928), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n943), .B1(new_n948), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n903), .B1(KEYINPUT50), .B2(new_n905), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n495), .A2(new_n500), .A3(new_n958), .A4(new_n891), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n946), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n945), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n952), .B1(new_n961), .B2(new_n928), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n913), .A2(new_n890), .A3(G2078), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n920), .B1(new_n963), .B2(new_n897), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n964), .B(new_n900), .C1(new_n909), .C2(new_n908), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n956), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n892), .A2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(G2084), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n896), .A4(new_n906), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n742), .B1(new_n911), .B2(new_n913), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT119), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT119), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(G168), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT120), .ZN(new_n976));
  AND2_X1   g551(.A1(KEYINPUT51), .A2(G8), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n975), .B2(new_n977), .ZN(new_n979));
  AOI211_X1 g554(.A(new_n928), .B(G286), .C1(new_n969), .C2(new_n970), .ZN(new_n980));
  NOR2_X1   g555(.A1(G168), .A2(new_n928), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n980), .A2(KEYINPUT51), .A3(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  AOI211_X1 g558(.A(new_n928), .B(G168), .C1(new_n973), .C2(new_n974), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n921), .B(new_n966), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(KEYINPUT57), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n558), .A2(new_n560), .A3(new_n562), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(KEYINPUT57), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT56), .B(G2072), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n894), .A2(new_n898), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1956), .B1(new_n957), .B2(new_n959), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1956), .ZN(new_n997));
  INV_X1    g572(.A(new_n959), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n905), .A2(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n896), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n997), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n894), .A2(new_n898), .A3(new_n992), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n990), .A3(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(new_n595), .ZN(new_n1004));
  INV_X1    g579(.A(G2067), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n907), .A2(new_n748), .B1(new_n1005), .B2(new_n927), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n996), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT61), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n995), .A2(KEYINPUT117), .A3(new_n1009), .A4(new_n1003), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1003), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1013), .A2(new_n1009), .B1(new_n995), .B2(new_n1003), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(G1341), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n903), .B2(new_n905), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT114), .B(new_n1016), .C1(new_n903), .C2(new_n905), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1996), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n894), .A2(new_n898), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT112), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n894), .A2(new_n898), .A3(new_n1025), .A4(new_n1022), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1021), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n541), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1027), .A2(KEYINPUT116), .A3(new_n1028), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1011), .A2(new_n1014), .B1(new_n1029), .B2(KEYINPUT59), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1021), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n896), .A2(new_n897), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n893), .B2(new_n892), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1025), .B1(new_n1033), .B2(new_n1022), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1026), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n541), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1028), .B1(new_n1040), .B2(new_n1031), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(KEYINPUT59), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1038), .A2(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT118), .B1(new_n1030), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1029), .B2(KEYINPUT115), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1013), .A2(new_n1009), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n995), .A2(new_n1003), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1010), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1038), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1046), .A2(new_n1050), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1006), .B1(KEYINPUT60), .B2(new_n595), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1044), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n985), .B1(new_n1008), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n686), .A2(new_n922), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT108), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n937), .B1(new_n942), .B2(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1062), .A2(KEYINPUT109), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(KEYINPUT109), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1063), .A2(new_n929), .A3(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n956), .A2(KEYINPUT110), .A3(new_n980), .A4(new_n962), .ZN(new_n1066));
  INV_X1    g641(.A(new_n943), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n948), .A2(new_n954), .A3(new_n953), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n962), .A3(new_n980), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT110), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1066), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n948), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(new_n1074), .B2(new_n952), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n956), .A2(new_n980), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1065), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1068), .A2(new_n943), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n889), .B1(new_n1059), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1058), .A2(new_n1008), .ZN(new_n1082));
  INV_X1    g657(.A(new_n985), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1078), .B(new_n1065), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(KEYINPUT123), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n975), .A2(new_n977), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT120), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n1089));
  INV_X1    g664(.A(new_n982), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n984), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(KEYINPUT62), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n956), .A2(new_n962), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(KEYINPUT62), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1096), .A2(G171), .A3(new_n919), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1081), .A2(new_n1086), .A3(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n769), .B(G2067), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n912), .A2(new_n903), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT105), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n732), .B(G1996), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n676), .A2(new_n678), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n676), .A2(new_n678), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1101), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(G290), .B(G1986), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1101), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1099), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1101), .A2(new_n1022), .ZN(new_n1113));
  NAND2_X1  g688(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1113), .B(new_n1114), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1101), .B1(new_n1100), .B2(new_n732), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1115), .B(new_n1116), .C1(KEYINPUT124), .C2(KEYINPUT46), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT125), .Z(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT47), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n769), .A2(G2067), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1101), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1122), .A2(G1986), .A3(G290), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1124));
  XNOR2_X1  g699(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1121), .A2(new_n1122), .B1(new_n1109), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1112), .A2(new_n1127), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g703(.A1(new_n827), .A2(new_n455), .A3(new_n630), .A4(new_n648), .ZN(new_n1130));
  NOR3_X1   g704(.A1(new_n1130), .A2(new_n887), .A3(G229), .ZN(G308));
  INV_X1    g705(.A(G308), .ZN(G225));
endmodule


