//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G141gat), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT77), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n214), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT78), .A2(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n206), .B1(new_n223), .B2(new_n205), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n214), .B1(new_n218), .B2(KEYINPUT2), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n216), .A2(new_n220), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227));
  INV_X1    g026(.A(G197gat), .ZN(new_n228));
  INV_X1    g027(.A(G204gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G197gat), .A2(G204gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232));
  NAND2_X1  g031(.A1(G211gat), .A2(G218gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n230), .A2(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n227), .B1(new_n234), .B2(KEYINPUT73), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n231), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n232), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT73), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n242), .B1(new_n234), .B2(new_n227), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n234), .A2(new_n242), .A3(new_n227), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n241), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT29), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n226), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n226), .B2(new_n249), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(new_n246), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n204), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n251), .B2(new_n246), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n215), .B1(new_n211), .B2(new_n212), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n209), .A2(KEYINPUT77), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n220), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n224), .A2(new_n225), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n249), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n247), .ZN(new_n262));
  XOR2_X1   g061(.A(G211gat), .B(G218gat), .Z(new_n263));
  OAI21_X1  g062(.A(KEYINPUT74), .B1(new_n238), .B2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n264), .A2(new_n244), .B1(new_n235), .B2(new_n240), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(KEYINPUT83), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n256), .A2(new_n203), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n238), .A2(new_n263), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n245), .B2(new_n243), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n247), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT3), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(KEYINPUT82), .A3(new_n247), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n226), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n253), .B(new_n254), .C1(new_n267), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n264), .A2(new_n244), .B1(new_n263), .B2(new_n238), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n277), .B2(KEYINPUT29), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(new_n273), .A3(new_n249), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n260), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n262), .A2(new_n265), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n204), .B1(new_n282), .B2(new_n255), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n283), .A3(new_n266), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n254), .B1(new_n284), .B2(new_n253), .ZN(new_n285));
  XOR2_X1   g084(.A(G78gat), .B(G106gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(G50gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n287), .B(G22gat), .Z(new_n288));
  XOR2_X1   g087(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n276), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n253), .B1(new_n267), .B2(new_n274), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT84), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n294), .B2(new_n275), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n202), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n291), .B1(new_n276), .B2(new_n285), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n275), .A3(new_n290), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT85), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT24), .ZN(new_n302));
  NOR2_X1   g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n311), .B1(KEYINPUT23), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n310), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(KEYINPUT24), .A3(new_n301), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n313), .A2(new_n320), .A3(new_n306), .A4(new_n308), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n320), .A2(new_n314), .A3(new_n306), .A4(new_n308), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(KEYINPUT25), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(G169gat), .B2(G176gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(new_n311), .ZN(new_n326));
  INV_X1    g125(.A(G169gat), .ZN(new_n327));
  INV_X1    g126(.A(G176gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT26), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n301), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n318), .B1(KEYINPUT65), .B2(KEYINPUT28), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT27), .B(G183gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n317), .A2(KEYINPUT27), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n334), .B1(new_n343), .B2(new_n336), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n331), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n316), .A2(new_n323), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n331), .A2(new_n344), .A3(new_n339), .A4(KEYINPUT66), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n352), .A2(new_n316), .A3(new_n323), .A4(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n350), .B1(new_n354), .B2(new_n347), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n246), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n349), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n316), .A2(new_n323), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(new_n348), .A3(new_n345), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n265), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(KEYINPUT75), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n357), .A2(new_n359), .A3(new_n362), .A4(new_n265), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G8gat), .B(G36gat), .Z(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT76), .ZN(new_n366));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n358), .A2(new_n348), .A3(new_n352), .A4(new_n353), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n265), .B1(new_n372), .B2(new_n350), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n368), .B(new_n363), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(KEYINPUT30), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n364), .A2(new_n376), .A3(new_n369), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379));
  XNOR2_X1  g178(.A(G57gat), .B(G85gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n387));
  INV_X1    g186(.A(G127gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(G134gat), .ZN(new_n389));
  INV_X1    g188(.A(G134gat), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT67), .B1(new_n390), .B2(G127gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n388), .A2(G134gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT68), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT68), .B(new_n389), .C1(new_n391), .C2(new_n392), .ZN(new_n396));
  INV_X1    g195(.A(G113gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G120gat), .ZN(new_n398));
  INV_X1    g197(.A(G120gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G113gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n396), .A3(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n390), .A2(G127gat), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n392), .A2(new_n405), .A3(KEYINPUT1), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT69), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n397), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n400), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(new_n280), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n411), .A2(new_n404), .B1(new_n259), .B2(new_n260), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n386), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n393), .A2(new_n394), .B1(new_n402), .B2(new_n401), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n417), .A2(new_n396), .B1(new_n410), .B2(new_n406), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(KEYINPUT3), .B2(new_n280), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n386), .B1(new_n419), .B2(new_n261), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n226), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n418), .A2(new_n226), .A3(KEYINPUT79), .A4(new_n421), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT4), .B1(new_n412), .B2(new_n280), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n416), .B1(new_n420), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n422), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n420), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n384), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n427), .A2(new_n420), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(new_n383), .A3(new_n431), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT6), .B(new_n384), .C1(new_n428), .C2(new_n432), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n378), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n354), .A2(new_n418), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n358), .A2(new_n412), .A3(new_n352), .A4(new_n353), .ZN(new_n445));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT32), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT70), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT70), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n451), .A3(KEYINPUT32), .ZN(new_n452));
  XNOR2_X1  g251(.A(G15gat), .B(G43gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(G71gat), .B(G99gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n448), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n448), .A2(KEYINPUT32), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n448), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n447), .B1(new_n444), .B2(new_n445), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n458), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n458), .B2(new_n464), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n443), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n464), .ZN(new_n474));
  INV_X1    g273(.A(new_n469), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(KEYINPUT36), .A3(new_n470), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n300), .A2(new_n442), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n374), .A2(KEYINPUT30), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n368), .B1(new_n361), .B2(new_n363), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n377), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n209), .A2(KEYINPUT77), .B1(KEYINPUT2), .B2(new_n214), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n219), .B1(new_n485), .B2(new_n213), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n224), .A2(new_n225), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT3), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(new_n261), .A3(new_n412), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT86), .B(new_n385), .C1(new_n430), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n412), .A2(new_n280), .A3(KEYINPUT4), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n421), .B1(new_n418), .B2(new_n226), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n494), .B2(new_n386), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n484), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n261), .A2(new_n419), .B1(new_n426), .B2(new_n422), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT86), .B1(new_n497), .B2(new_n385), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n494), .A2(new_n491), .A3(new_n386), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n413), .A2(new_n414), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(new_n385), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n503), .A3(new_n383), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n496), .A2(new_n503), .A3(KEYINPUT40), .A4(new_n383), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n483), .A2(new_n433), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n439), .A2(new_n440), .A3(new_n370), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n364), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n361), .A2(KEYINPUT37), .A3(new_n363), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n511), .A2(KEYINPUT38), .A3(new_n368), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT37), .B1(new_n361), .B2(new_n363), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n355), .A2(new_n265), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n357), .A2(new_n246), .A3(new_n359), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n515), .A2(KEYINPUT37), .A3(new_n516), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n514), .A2(new_n369), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n513), .B1(new_n518), .B2(KEYINPUT38), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n292), .A2(new_n295), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n508), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n476), .A2(new_n298), .A3(new_n297), .A4(new_n470), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT35), .B1(new_n523), .B2(new_n442), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n471), .A2(new_n472), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n377), .A2(new_n375), .B1(new_n439), .B2(new_n440), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT35), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n521), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n478), .A2(new_n522), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n530), .A2(KEYINPUT91), .ZN(new_n531));
  XOR2_X1   g330(.A(G57gat), .B(G64gat), .Z(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(KEYINPUT91), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n530), .B(KEYINPUT91), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n534), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n530), .B(new_n540), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n541), .B(new_n532), .C1(KEYINPUT92), .C2(new_n535), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n543), .A2(KEYINPUT21), .ZN(new_n544));
  XOR2_X1   g343(.A(G127gat), .B(G155gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(G1gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT16), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(G1gat), .B2(new_n547), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G8gat), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(KEYINPUT21), .B2(new_n543), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n546), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT94), .ZN(new_n556));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT93), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n554), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G99gat), .B(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT98), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(G92gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G99gat), .ZN(new_n571));
  INV_X1    g370(.A(G106gat), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT8), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT99), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n570), .A2(new_n576), .A3(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(KEYINPUT96), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n581), .B2(new_n583), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n564), .B1(new_n578), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n570), .A2(new_n576), .A3(new_n573), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n576), .B1(new_n570), .B2(new_n573), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n585), .B(new_n564), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592));
  NAND2_X1  g391(.A1(G29gat), .A2(G36gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n594));
  NOR3_X1   g393(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT88), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT14), .ZN(new_n598));
  INV_X1    g397(.A(G29gat), .ZN(new_n599));
  INV_X1    g398(.A(G36gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(KEYINPUT88), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n593), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G43gat), .B(G50gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT15), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n604), .A2(KEYINPUT15), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n601), .A2(new_n594), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n608), .A2(new_n605), .A3(new_n593), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n591), .B1(new_n592), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT89), .B1(new_n611), .B2(new_n592), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT89), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n607), .A2(new_n610), .A3(new_n614), .A4(KEYINPUT17), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G190gat), .B(G218gat), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n620), .B(KEYINPUT95), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n591), .A2(new_n611), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n617), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n619), .B1(new_n617), .B2(new_n623), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OR3_X1    g428(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n629), .B1(new_n624), .B2(new_n625), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n539), .A2(new_n542), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(new_n586), .B2(new_n590), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n637));
  INV_X1    g436(.A(new_n564), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n543), .A3(new_n589), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n543), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n635), .A2(new_n640), .ZN(new_n646));
  INV_X1    g445(.A(new_n644), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT100), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n645), .A2(new_n654), .A3(new_n648), .A4(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n647), .B1(new_n641), .B2(new_n642), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n646), .B2(new_n647), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n658), .A2(new_n651), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G113gat), .B(G141gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G197gat), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT11), .B(G169gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT12), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n552), .B(new_n611), .ZN(new_n668));
  NAND2_X1  g467(.A1(G229gat), .A2(G233gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT13), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n552), .A2(new_n611), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n552), .B1(new_n592), .B2(new_n611), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n616), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT90), .B1(new_n674), .B2(new_n669), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT18), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n669), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n678), .B(new_n672), .C1(new_n616), .C2(new_n673), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(KEYINPUT90), .A3(KEYINPUT18), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n667), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT18), .B1(new_n679), .B2(KEYINPUT90), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n675), .A2(new_n676), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n666), .A4(new_n671), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n661), .A2(new_n685), .ZN(new_n686));
  OR4_X1    g485(.A1(new_n529), .A2(new_n563), .A3(new_n633), .A4(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n441), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(new_n548), .ZN(G1324gat));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n378), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n691), .A2(G8gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT16), .B(G8gat), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT42), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(KEYINPUT42), .B2(new_n694), .ZN(G1325gat));
  NAND2_X1  g495(.A1(new_n473), .A2(new_n477), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n687), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n525), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n699), .A2(G15gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n687), .B2(new_n700), .ZN(G1326gat));
  INV_X1    g500(.A(new_n300), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT43), .B(G22gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n529), .B2(new_n632), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n292), .A2(new_n295), .A3(new_n202), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT85), .B1(new_n297), .B2(new_n298), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n442), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n509), .A2(new_n519), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n506), .A2(new_n507), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n375), .A2(new_n433), .A3(new_n377), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n521), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n710), .B(new_n697), .C1(new_n711), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n524), .A2(new_n528), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(KEYINPUT44), .A3(new_n633), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n707), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n562), .B(KEYINPUT101), .Z(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n686), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n441), .ZN(new_n724));
  INV_X1    g523(.A(new_n685), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n725), .A2(new_n660), .A3(new_n632), .A4(new_n562), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n441), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n599), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT102), .Z(G1328gat));
  NAND3_X1  g531(.A1(new_n727), .A2(new_n600), .A3(new_n483), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT46), .Z(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n723), .B2(new_n378), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n697), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n727), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n699), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n723), .A2(new_n738), .B1(new_n740), .B2(G43gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g541(.A1(new_n719), .A2(new_n300), .A3(new_n722), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G50gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n702), .A2(G50gat), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n727), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(KEYINPUT48), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n521), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n707), .A2(new_n718), .A3(new_n749), .A4(new_n722), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n746), .B1(G50gat), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT103), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n747), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n755), .B(new_n756), .C1(new_n751), .C2(new_n752), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n754), .A2(new_n757), .ZN(G1331gat));
  NAND3_X1  g557(.A1(new_n725), .A2(new_n632), .A3(new_n562), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n661), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT104), .Z(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n717), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n728), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g564(.A1(new_n762), .A2(new_n378), .ZN(new_n766));
  NOR2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  AND2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n766), .B2(new_n767), .ZN(G1333gat));
  NOR3_X1   g569(.A1(new_n762), .A2(G71gat), .A3(new_n699), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n763), .A2(new_n737), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(G71gat), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n763), .A2(new_n300), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g575(.A1(new_n685), .A2(new_n562), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n661), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n707), .A2(new_n718), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT105), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n707), .A2(new_n718), .A3(new_n782), .A4(new_n779), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n781), .A2(new_n728), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n717), .A2(new_n633), .A3(new_n777), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n660), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n728), .A2(new_n569), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n784), .A2(new_n569), .B1(new_n789), .B2(new_n790), .ZN(G1336gat));
  NAND2_X1  g590(.A1(new_n566), .A2(new_n568), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n780), .B2(new_n378), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n378), .A2(G92gat), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n793), .B(new_n794), .C1(new_n789), .C2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n483), .A3(new_n783), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n798), .A2(KEYINPUT106), .A3(new_n792), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT106), .B1(new_n798), .B2(new_n792), .ZN(new_n800));
  INV_X1    g599(.A(new_n785), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n786), .B1(new_n801), .B2(KEYINPUT107), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT107), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n803), .A3(KEYINPUT51), .ZN(new_n804));
  AND4_X1   g603(.A1(new_n660), .A2(new_n802), .A3(new_n804), .A4(new_n795), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n799), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n797), .B1(new_n806), .B2(new_n794), .ZN(G1337gat));
  AND3_X1   g606(.A1(new_n781), .A2(new_n737), .A3(new_n783), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n525), .A2(new_n571), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n808), .A2(new_n571), .B1(new_n789), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT108), .ZN(G1338gat));
  AND2_X1   g610(.A1(new_n802), .A2(new_n804), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n749), .A2(new_n572), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n661), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n781), .A2(new_n300), .A3(new_n783), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n812), .A2(new_n814), .B1(new_n815), .B2(G106gat), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  INV_X1    g616(.A(new_n780), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n572), .B1(new_n818), .B2(new_n749), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n789), .B2(new_n813), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n816), .A2(new_n817), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  NAND3_X1  g620(.A1(new_n641), .A2(new_n642), .A3(new_n647), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT109), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT109), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n641), .A2(new_n642), .A3(new_n824), .A4(new_n647), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n823), .A2(new_n645), .A3(KEYINPUT54), .A4(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n651), .B1(new_n657), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n826), .A2(KEYINPUT110), .A3(KEYINPUT55), .A4(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n656), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n828), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n830), .A2(new_n685), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n674), .A2(new_n669), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n668), .A2(new_n670), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n665), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n660), .A2(new_n684), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n633), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n836), .A2(new_n833), .A3(new_n656), .A4(new_n829), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n630), .A2(new_n631), .A3(new_n684), .A4(new_n840), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n720), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n759), .A2(new_n660), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n300), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n849), .A2(new_n728), .A3(new_n378), .A4(new_n525), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n725), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n441), .B1(new_n846), .B2(new_n848), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n523), .A2(new_n483), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT111), .Z(new_n855));
  NAND2_X1  g654(.A1(new_n685), .A2(new_n397), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(G1340gat));
  OAI21_X1  g656(.A(G120gat), .B1(new_n850), .B2(new_n661), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n660), .A2(new_n399), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n860), .A2(new_n861), .B1(new_n855), .B2(new_n862), .ZN(G1341gat));
  NOR3_X1   g662(.A1(new_n850), .A2(new_n388), .A3(new_n720), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n854), .A2(KEYINPUT113), .A3(new_n563), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(G127gat), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT113), .B1(new_n854), .B2(new_n563), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(G1342gat));
  NAND2_X1  g667(.A1(new_n633), .A2(new_n390), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n854), .A2(KEYINPUT56), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n850), .B2(new_n632), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT56), .B1(new_n854), .B2(new_n869), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT114), .Z(G1343gat));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n728), .A2(new_n378), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n737), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT115), .ZN(new_n879));
  XNOR2_X1  g678(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n831), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n830), .A2(new_n685), .A3(new_n836), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n633), .B1(new_n882), .B2(new_n841), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n563), .B1(new_n883), .B2(new_n845), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n702), .B1(new_n884), .B2(new_n848), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n879), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n841), .B1(new_n843), .B2(new_n725), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n845), .B1(new_n888), .B2(new_n632), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n848), .B1(new_n889), .B2(new_n721), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n749), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n876), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n836), .A2(new_n656), .A3(new_n829), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n685), .A2(new_n881), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n841), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n632), .ZN(new_n897));
  INV_X1    g696(.A(new_n845), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n562), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n300), .B1(new_n899), .B2(new_n847), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT57), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n521), .B1(new_n846), .B2(new_n848), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n886), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT117), .A4(new_n879), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n893), .A2(new_n685), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n697), .A2(new_n749), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n378), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n852), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n725), .A2(G141gat), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n905), .A2(new_n223), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n901), .A2(new_n903), .A3(new_n685), .A4(new_n879), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT58), .B1(new_n913), .B2(new_n223), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n852), .A2(new_n909), .A3(new_n911), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n914), .B2(new_n917), .ZN(new_n920));
  OAI22_X1  g719(.A1(new_n875), .A2(new_n912), .B1(new_n919), .B2(new_n920), .ZN(G1344gat));
  XOR2_X1   g720(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n922));
  AOI211_X1 g721(.A(G148gat), .B(new_n922), .C1(new_n910), .C2(new_n660), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n886), .B(new_n300), .C1(new_n899), .C2(new_n847), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n661), .A2(new_n922), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n924), .A2(new_n879), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n893), .A2(new_n660), .A3(new_n904), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(KEYINPUT59), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n923), .B1(new_n929), .B2(G148gat), .ZN(G1345gat));
  INV_X1    g729(.A(G155gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n931), .A3(new_n562), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n893), .A2(new_n721), .A3(new_n904), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n931), .ZN(G1346gat));
  INV_X1    g733(.A(G162gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n910), .A2(new_n935), .A3(new_n633), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n893), .A2(new_n633), .A3(new_n904), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G162gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(KEYINPUT122), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(G1347gat));
  NAND2_X1  g740(.A1(new_n483), .A2(new_n441), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n699), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n849), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n849), .A2(new_n948), .A3(new_n944), .A4(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n950), .A2(new_n327), .A3(new_n725), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n728), .B1(new_n846), .B2(new_n848), .ZN(new_n952));
  AND4_X1   g751(.A1(new_n521), .A2(new_n952), .A3(new_n483), .A4(new_n525), .ZN(new_n953));
  AOI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n685), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n951), .A2(new_n954), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n950), .B2(new_n661), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n328), .A3(new_n660), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1349gat));
  OAI21_X1  g757(.A(G183gat), .B1(new_n950), .B2(new_n720), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n953), .A2(new_n338), .A3(new_n562), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT60), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n959), .A2(new_n963), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n953), .A2(new_n318), .A3(new_n633), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT125), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n318), .B1(new_n968), .B2(KEYINPUT61), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n969), .B1(new_n950), .B2(new_n632), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n970), .A2(KEYINPUT126), .A3(new_n971), .ZN(new_n972));
  OAI221_X1 g771(.A(new_n969), .B1(new_n968), .B2(KEYINPUT61), .C1(new_n950), .C2(new_n632), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n967), .A2(new_n972), .A3(new_n973), .ZN(G1351gat));
  AND4_X1   g773(.A1(new_n749), .A2(new_n952), .A3(new_n483), .A4(new_n697), .ZN(new_n975));
  AOI21_X1  g774(.A(G197gat), .B1(new_n975), .B2(new_n685), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n737), .A2(new_n942), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n925), .B(new_n977), .C1(new_n902), .C2(new_n886), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n978), .A2(new_n228), .A3(new_n725), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n976), .A2(new_n979), .ZN(G1352gat));
  NAND3_X1  g779(.A1(new_n975), .A2(new_n229), .A3(new_n660), .ZN(new_n981));
  XOR2_X1   g780(.A(new_n981), .B(KEYINPUT62), .Z(new_n982));
  OAI21_X1  g781(.A(G204gat), .B1(new_n978), .B2(new_n661), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1353gat));
  INV_X1    g783(.A(G211gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n975), .A2(new_n985), .A3(new_n562), .ZN(new_n986));
  OAI211_X1 g785(.A(KEYINPUT63), .B(G211gat), .C1(new_n978), .C2(new_n563), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n924), .A2(new_n562), .A3(new_n925), .A4(new_n977), .ZN(new_n989));
  AOI21_X1  g788(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n986), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g792(.A(KEYINPUT127), .B(new_n986), .C1(new_n988), .C2(new_n990), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1354gat));
  INV_X1    g794(.A(G218gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n975), .A2(new_n996), .A3(new_n633), .ZN(new_n997));
  OAI21_X1  g796(.A(G218gat), .B1(new_n978), .B2(new_n632), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(G1355gat));
endmodule


