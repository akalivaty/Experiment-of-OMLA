

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593;

  XNOR2_X1 U322 ( .A(KEYINPUT25), .B(KEYINPUT104), .ZN(n464) );
  XOR2_X1 U323 ( .A(G120GAT), .B(G71GAT), .Z(n438) );
  XNOR2_X1 U324 ( .A(n422), .B(n292), .ZN(n352) );
  XNOR2_X1 U325 ( .A(n482), .B(KEYINPUT110), .ZN(n483) );
  XOR2_X1 U326 ( .A(n318), .B(n317), .Z(n290) );
  AND2_X1 U327 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U329 ( .A(KEYINPUT45), .B(KEYINPUT66), .ZN(n362) );
  XNOR2_X1 U330 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U331 ( .A(n438), .B(n291), .ZN(n311) );
  XNOR2_X1 U332 ( .A(n465), .B(n464), .ZN(n470) );
  XNOR2_X1 U333 ( .A(n311), .B(n343), .ZN(n313) );
  XNOR2_X1 U334 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U335 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n310) );
  XNOR2_X1 U336 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U337 ( .A(n319), .B(n290), .ZN(n320) );
  INV_X1 U338 ( .A(KEYINPUT37), .ZN(n482) );
  XNOR2_X1 U339 ( .A(n321), .B(n320), .ZN(n327) );
  XNOR2_X1 U340 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U341 ( .A(KEYINPUT36), .B(n553), .Z(n590) );
  XNOR2_X1 U342 ( .A(n367), .B(KEYINPUT41), .ZN(n368) );
  XNOR2_X1 U343 ( .A(n484), .B(n483), .ZN(n524) );
  XNOR2_X1 U344 ( .A(n583), .B(n368), .ZN(n561) );
  XNOR2_X1 U345 ( .A(n361), .B(n360), .ZN(n553) );
  XNOR2_X1 U346 ( .A(n458), .B(KEYINPUT58), .ZN(n459) );
  XNOR2_X1 U347 ( .A(n488), .B(G43GAT), .ZN(n489) );
  XNOR2_X1 U348 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n490), .B(n489), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT8), .B(G43GAT), .Z(n294) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G29GAT), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U353 ( .A(KEYINPUT7), .B(n295), .Z(n359) );
  XOR2_X1 U354 ( .A(G169GAT), .B(G8GAT), .Z(n391) );
  XOR2_X1 U355 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n297) );
  XNOR2_X1 U356 ( .A(G197GAT), .B(G113GAT), .ZN(n296) );
  XNOR2_X1 U357 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U358 ( .A(n391), .B(n298), .Z(n300) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U361 ( .A(KEYINPUT30), .B(KEYINPUT74), .Z(n302) );
  XNOR2_X1 U362 ( .A(KEYINPUT71), .B(KEYINPUT73), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U364 ( .A(n304), .B(n303), .Z(n308) );
  XNOR2_X1 U365 ( .A(G50GAT), .B(G22GAT), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n305), .B(G141GAT), .ZN(n423) );
  XNOR2_X1 U367 ( .A(G15GAT), .B(G1GAT), .ZN(n306) );
  XNOR2_X1 U368 ( .A(n306), .B(KEYINPUT72), .ZN(n344) );
  XNOR2_X1 U369 ( .A(n423), .B(n344), .ZN(n307) );
  XNOR2_X1 U370 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n359), .B(n309), .ZN(n579) );
  XNOR2_X1 U372 ( .A(KEYINPUT75), .B(n579), .ZN(n485) );
  INV_X1 U373 ( .A(n485), .ZN(n544) );
  XNOR2_X1 U374 ( .A(n310), .B(KEYINPUT76), .ZN(n343) );
  INV_X1 U375 ( .A(KEYINPUT79), .ZN(n312) );
  NAND2_X1 U376 ( .A1(n313), .A2(n312), .ZN(n316) );
  INV_X1 U377 ( .A(n313), .ZN(n314) );
  NAND2_X1 U378 ( .A1(n314), .A2(KEYINPUT79), .ZN(n315) );
  NAND2_X1 U379 ( .A1(n316), .A2(n315), .ZN(n321) );
  XOR2_X1 U380 ( .A(G176GAT), .B(G64GAT), .Z(n390) );
  XNOR2_X1 U381 ( .A(n390), .B(KEYINPUT32), .ZN(n319) );
  XOR2_X1 U382 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n318) );
  XNOR2_X1 U383 ( .A(KEYINPUT77), .B(KEYINPUT80), .ZN(n317) );
  XOR2_X1 U384 ( .A(G78GAT), .B(G148GAT), .Z(n323) );
  XNOR2_X1 U385 ( .A(G106GAT), .B(G204GAT), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n434) );
  XOR2_X1 U387 ( .A(KEYINPUT78), .B(G92GAT), .Z(n325) );
  XNOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n353) );
  XNOR2_X1 U390 ( .A(n434), .B(n353), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n583) );
  XOR2_X1 U392 ( .A(G155GAT), .B(G78GAT), .Z(n329) );
  XNOR2_X1 U393 ( .A(G22GAT), .B(G211GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U395 ( .A(G71GAT), .B(G183GAT), .Z(n331) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(G127GAT), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U398 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U399 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n335) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U402 ( .A(KEYINPUT85), .B(n336), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U404 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n340) );
  XNOR2_X1 U405 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U407 ( .A(n342), .B(n341), .Z(n346) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n587) );
  XOR2_X1 U410 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n348) );
  XNOR2_X1 U411 ( .A(G218GAT), .B(G106GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U413 ( .A(n349), .B(KEYINPUT67), .Z(n351) );
  XOR2_X1 U414 ( .A(G190GAT), .B(G134GAT), .Z(n439) );
  XNOR2_X1 U415 ( .A(G50GAT), .B(n439), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U417 ( .A(KEYINPUT81), .B(G162GAT), .Z(n422) );
  XOR2_X1 U418 ( .A(n355), .B(n354), .Z(n361) );
  XOR2_X1 U419 ( .A(KEYINPUT11), .B(KEYINPUT68), .Z(n357) );
  XNOR2_X1 U420 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  NAND2_X1 U423 ( .A1(n587), .A2(n590), .ZN(n363) );
  NOR2_X1 U424 ( .A1(n583), .A2(n364), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n365), .B(KEYINPUT117), .ZN(n366) );
  OR2_X1 U426 ( .A1(n544), .A2(n366), .ZN(n375) );
  INV_X1 U427 ( .A(KEYINPUT64), .ZN(n367) );
  NAND2_X1 U428 ( .A1(n579), .A2(n561), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT46), .ZN(n371) );
  INV_X1 U430 ( .A(n553), .ZN(n565) );
  NOR2_X1 U431 ( .A1(n565), .A2(n587), .ZN(n370) );
  NAND2_X1 U432 ( .A1(n371), .A2(n370), .ZN(n373) );
  INV_X1 U433 ( .A(KEYINPUT47), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n374) );
  AND2_X1 U435 ( .A1(n375), .A2(n374), .ZN(n376) );
  XOR2_X1 U436 ( .A(KEYINPUT48), .B(n376), .Z(n539) );
  XOR2_X1 U437 ( .A(KEYINPUT94), .B(KEYINPUT21), .Z(n378) );
  XNOR2_X1 U438 ( .A(G218GAT), .B(KEYINPUT92), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U440 ( .A(n379), .B(KEYINPUT93), .Z(n381) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n430) );
  XOR2_X1 U443 ( .A(G183GAT), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U444 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n449) );
  XOR2_X1 U446 ( .A(KEYINPUT100), .B(n449), .Z(n385) );
  NAND2_X1 U447 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U449 ( .A(G92GAT), .B(G204GAT), .Z(n387) );
  XNOR2_X1 U450 ( .A(G36GAT), .B(G190GAT), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U452 ( .A(n389), .B(n388), .Z(n393) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U455 ( .A(n430), .B(n394), .Z(n501) );
  NAND2_X1 U456 ( .A1(n539), .A2(n501), .ZN(n396) );
  XOR2_X1 U457 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n420) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XOR2_X1 U460 ( .A(G85GAT), .B(G148GAT), .Z(n398) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(G134GAT), .ZN(n397) );
  XNOR2_X1 U462 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U463 ( .A(G29GAT), .B(G162GAT), .Z(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n419) );
  XOR2_X1 U466 ( .A(G155GAT), .B(KEYINPUT2), .Z(n404) );
  XNOR2_X1 U467 ( .A(KEYINPUT3), .B(KEYINPUT95), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n433) );
  XOR2_X1 U469 ( .A(KEYINPUT99), .B(n433), .Z(n409) );
  XOR2_X1 U470 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n406) );
  XNOR2_X1 U471 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U473 ( .A(G113GAT), .B(n407), .Z(n453) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(n453), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n417) );
  XOR2_X1 U476 ( .A(KEYINPUT98), .B(G57GAT), .Z(n411) );
  XNOR2_X1 U477 ( .A(KEYINPUT97), .B(KEYINPUT1), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U479 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n413) );
  XNOR2_X1 U480 ( .A(G120GAT), .B(KEYINPUT5), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U482 ( .A(n415), .B(n414), .Z(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n526) );
  NAND2_X1 U485 ( .A1(n420), .A2(n526), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n421), .B(KEYINPUT65), .ZN(n576) );
  XOR2_X1 U487 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n425) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT96), .Z(n427) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U493 ( .A(n429), .B(n428), .Z(n432) );
  XNOR2_X1 U494 ( .A(n430), .B(KEYINPUT23), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U496 ( .A(n434), .B(n433), .Z(n435) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n475) );
  NAND2_X1 U498 ( .A1(n576), .A2(n475), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n437), .B(KEYINPUT55), .ZN(n454) );
  XOR2_X1 U500 ( .A(G99GAT), .B(n438), .Z(n441) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U503 ( .A(G176GAT), .B(KEYINPUT89), .Z(n443) );
  XNOR2_X1 U504 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n445) );
  AND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XOR2_X1 U507 ( .A(n449), .B(n448), .Z(n451) );
  XNOR2_X1 U508 ( .A(G169GAT), .B(G15GAT), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n477) );
  NAND2_X1 U511 ( .A1(n454), .A2(n477), .ZN(n573) );
  NOR2_X1 U512 ( .A1(n573), .A2(n485), .ZN(n457) );
  XNOR2_X1 U513 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(KEYINPUT124), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(G1348GAT) );
  NOR2_X1 U516 ( .A1(n573), .A2(n553), .ZN(n460) );
  INV_X1 U517 ( .A(G190GAT), .ZN(n458) );
  INV_X1 U518 ( .A(n477), .ZN(n540) );
  NAND2_X1 U519 ( .A1(n501), .A2(n477), .ZN(n462) );
  INV_X1 U520 ( .A(KEYINPUT103), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n463), .A2(n475), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n477), .A2(n475), .ZN(n467) );
  XNOR2_X1 U524 ( .A(KEYINPUT26), .B(KEYINPUT101), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n467), .B(n466), .ZN(n578) );
  XOR2_X1 U526 ( .A(n501), .B(KEYINPUT27), .Z(n474) );
  NOR2_X1 U527 ( .A1(n578), .A2(n474), .ZN(n468) );
  XNOR2_X1 U528 ( .A(KEYINPUT102), .B(n468), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT105), .ZN(n491) );
  INV_X1 U531 ( .A(n587), .ZN(n574) );
  AND2_X1 U532 ( .A1(n574), .A2(n590), .ZN(n473) );
  AND2_X1 U533 ( .A1(n526), .A2(n473), .ZN(n472) );
  NAND2_X1 U534 ( .A1(n491), .A2(n472), .ZN(n481) );
  INV_X1 U535 ( .A(n473), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n474), .A2(n526), .ZN(n538) );
  XNOR2_X1 U537 ( .A(KEYINPUT28), .B(KEYINPUT69), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n476), .B(n475), .ZN(n543) );
  NOR2_X1 U539 ( .A1(n543), .A2(n477), .ZN(n478) );
  NAND2_X1 U540 ( .A1(n538), .A2(n478), .ZN(n492) );
  OR2_X1 U541 ( .A1(n479), .A2(n492), .ZN(n480) );
  NAND2_X1 U542 ( .A1(n481), .A2(n480), .ZN(n484) );
  NOR2_X1 U543 ( .A1(n485), .A2(n583), .ZN(n497) );
  NAND2_X1 U544 ( .A1(n524), .A2(n497), .ZN(n486) );
  XOR2_X1 U545 ( .A(n486), .B(KEYINPUT111), .Z(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT38), .B(n487), .ZN(n513) );
  NOR2_X1 U547 ( .A1(n540), .A2(n513), .ZN(n490) );
  INV_X1 U548 ( .A(KEYINPUT40), .ZN(n488) );
  NAND2_X1 U549 ( .A1(n491), .A2(n526), .ZN(n493) );
  NAND2_X1 U550 ( .A1(n493), .A2(n492), .ZN(n496) );
  NAND2_X1 U551 ( .A1(n553), .A2(n587), .ZN(n494) );
  XOR2_X1 U552 ( .A(KEYINPUT16), .B(n494), .Z(n495) );
  AND2_X1 U553 ( .A1(n496), .A2(n495), .ZN(n515) );
  NAND2_X1 U554 ( .A1(n497), .A2(n515), .ZN(n507) );
  NOR2_X1 U555 ( .A1(n526), .A2(n507), .ZN(n499) );
  XNOR2_X1 U556 ( .A(KEYINPUT34), .B(KEYINPUT106), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U558 ( .A(G1GAT), .B(n500), .Z(G1324GAT) );
  INV_X1 U559 ( .A(n501), .ZN(n528) );
  NOR2_X1 U560 ( .A1(n528), .A2(n507), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G8GAT), .B(KEYINPUT107), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(G1325GAT) );
  NOR2_X1 U563 ( .A1(n540), .A2(n507), .ZN(n505) );
  XNOR2_X1 U564 ( .A(KEYINPUT108), .B(KEYINPUT35), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G15GAT), .B(n506), .ZN(G1326GAT) );
  INV_X1 U567 ( .A(n543), .ZN(n534) );
  NOR2_X1 U568 ( .A1(n534), .A2(n507), .ZN(n509) );
  XNOR2_X1 U569 ( .A(G22GAT), .B(KEYINPUT109), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(G1327GAT) );
  NOR2_X1 U571 ( .A1(n513), .A2(n526), .ZN(n511) );
  XNOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(G1328GAT) );
  NOR2_X1 U574 ( .A1(n513), .A2(n528), .ZN(n512) );
  XOR2_X1 U575 ( .A(G36GAT), .B(n512), .Z(G1329GAT) );
  NOR2_X1 U576 ( .A1(n534), .A2(n513), .ZN(n514) );
  XOR2_X1 U577 ( .A(G50GAT), .B(n514), .Z(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT112), .B(n561), .Z(n568) );
  NOR2_X1 U579 ( .A1(n579), .A2(n568), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n525), .A2(n515), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n526), .A2(n520), .ZN(n516) );
  XOR2_X1 U582 ( .A(G57GAT), .B(n516), .Z(n517) );
  XNOR2_X1 U583 ( .A(KEYINPUT42), .B(n517), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n528), .A2(n520), .ZN(n518) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n518), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n540), .A2(n520), .ZN(n519) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n519), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n534), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U591 ( .A(G78GAT), .B(n523), .Z(G1335GAT) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n533) );
  NOR2_X1 U593 ( .A1(n526), .A2(n533), .ZN(n527) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U595 ( .A1(n528), .A2(n533), .ZN(n529) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(n529), .Z(n530) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  NOR2_X1 U598 ( .A1(n540), .A2(n533), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(G1338GAT) );
  NOR2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT44), .B(KEYINPUT116), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U604 ( .A(G106GAT), .B(n537), .Z(G1339GAT) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n556) );
  NOR2_X1 U606 ( .A1(n540), .A2(n556), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT118), .B(n541), .Z(n542) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n548), .A2(n544), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n545), .ZN(G1340GAT) );
  INV_X1 U611 ( .A(n548), .ZN(n552) );
  NOR2_X1 U612 ( .A1(n568), .A2(n552), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U616 ( .A1(n548), .A2(n587), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NOR2_X1 U622 ( .A1(n578), .A2(n556), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n579), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n557), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n559) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT120), .B(n560), .Z(n563) );
  NAND2_X1 U629 ( .A1(n566), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n587), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n573), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT56), .Z(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(G183GAT), .B(n575), .Z(G1350GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  INV_X1 U643 ( .A(n576), .ZN(n577) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n591) );
  NAND2_X1 U645 ( .A1(n591), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n591), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U653 ( .A1(n591), .A2(n587), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

