//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT0), .B(G128), .Z(new_n193));
  INV_X1    g007(.A(KEYINPUT0), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  MUX2_X1   g011(.A(new_n193), .B(new_n196), .S(new_n197), .Z(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .A4(G104), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT80), .A3(G107), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT4), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G101), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT83), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT83), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n211), .A3(new_n208), .A4(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n214), .B(new_n203), .C1(new_n205), .C2(new_n206), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT82), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n201), .B1(new_n202), .B2(G104), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(new_n202), .A3(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n220), .A2(KEYINPUT82), .A3(new_n214), .A4(new_n203), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n224));
  AOI211_X1 g038(.A(new_n224), .B(new_n214), .C1(new_n220), .C2(new_n203), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT81), .B1(new_n207), .B2(G101), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n199), .B(new_n213), .C1(new_n223), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G137), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G134), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT11), .B1(new_n231), .B2(G137), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n229), .A3(G134), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n230), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G131), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(G137), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(KEYINPUT64), .A3(new_n236), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G143), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(G128), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n246), .B(new_n248), .C1(KEYINPUT1), .C2(new_n195), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n202), .A2(G104), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n204), .A2(G107), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n214), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n222), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT10), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n257), .B1(new_n217), .B2(new_n221), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT10), .A3(new_n254), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n228), .A2(new_n244), .A3(new_n261), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n262), .A2(KEYINPUT10), .A3(new_n254), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT10), .B1(new_n262), .B2(new_n254), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n269), .A2(KEYINPUT84), .A3(new_n244), .A4(new_n228), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  AND4_X1   g085(.A1(KEYINPUT64), .A2(new_n238), .A3(new_n236), .A4(new_n239), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT64), .B1(new_n235), .B2(new_n236), .ZN(new_n273));
  OAI22_X1  g087(.A1(new_n272), .A2(new_n273), .B1(new_n236), .B2(new_n235), .ZN(new_n274));
  INV_X1    g088(.A(new_n259), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n262), .A2(new_n254), .ZN(new_n276));
  OAI211_X1 g090(.A(KEYINPUT12), .B(new_n274), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n222), .A2(new_n258), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n253), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n259), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n282), .A2(KEYINPUT85), .A3(KEYINPUT12), .A4(new_n274), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT12), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(G110), .B(G140), .ZN(new_n288));
  INV_X1    g102(.A(G953), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G227), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n288), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n271), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT87), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT87), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n271), .A2(new_n287), .A3(new_n294), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n269), .A2(new_n228), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n274), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n291), .B1(new_n271), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n192), .B1(new_n301), .B2(new_n190), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n271), .A2(new_n298), .A3(new_n291), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n271), .A2(new_n287), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(new_n291), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT86), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT86), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n307), .B(new_n303), .C1(new_n304), .C2(new_n291), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(G469), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n189), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G128), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n313), .B(new_n314), .C1(G119), .C2(new_n195), .ZN(new_n315));
  OR3_X1    g129(.A1(new_n315), .A2(KEYINPUT76), .A3(G110), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT76), .B1(new_n315), .B2(G110), .ZN(new_n317));
  XOR2_X1   g131(.A(G119), .B(G128), .Z(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT24), .B(G110), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n316), .B(new_n317), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(G140), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT71), .A3(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g142(.A1(KEYINPUT72), .A2(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT72), .A2(G125), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G140), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT16), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT73), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n331), .A3(new_n334), .A4(KEYINPUT16), .ZN(new_n335));
  NOR2_X1   g149(.A1(KEYINPUT16), .A2(G140), .ZN(new_n336));
  AND2_X1   g150(.A1(KEYINPUT72), .A2(G125), .ZN(new_n337));
  NOR2_X1   g151(.A1(KEYINPUT72), .A2(G125), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT74), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n341), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n333), .A2(G146), .A3(new_n335), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n326), .A2(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n324), .A2(G140), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n322), .B(new_n344), .C1(G146), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n343), .A2(new_n335), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n337), .A2(new_n338), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n354), .A2(G140), .B1(new_n325), .B2(new_n327), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n334), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n245), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n344), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n319), .A2(new_n321), .B1(new_n315), .B2(G110), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n352), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n359), .ZN(new_n361));
  AOI211_X1 g175(.A(KEYINPUT75), .B(new_n361), .C1(new_n357), .C2(new_n344), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n351), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n289), .A2(G221), .A3(G234), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT79), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT22), .B(G137), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(KEYINPUT78), .B(new_n351), .C1(new_n360), .C2(new_n362), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n363), .A2(new_n370), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G234), .ZN(new_n375));
  OAI21_X1  g189(.A(G217), .B1(new_n375), .B2(G902), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n191), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n372), .A2(new_n191), .A3(new_n373), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n380), .A2(KEYINPUT25), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT25), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n372), .A2(new_n382), .A3(new_n191), .A4(new_n373), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n376), .B(KEYINPUT70), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n379), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(G237), .A2(G953), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G210), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n388), .B(KEYINPUT27), .Z(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT26), .B(G101), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT28), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n272), .A2(new_n273), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n231), .A3(G137), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT65), .B1(new_n231), .B2(G137), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n229), .A3(G134), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n394), .A2(new_n396), .A3(new_n397), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G131), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n252), .A3(new_n251), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n244), .A2(new_n198), .B1(new_n393), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n312), .A2(G116), .ZN(new_n404));
  INV_X1    g218(.A(G116), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G119), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT67), .ZN(new_n408));
  XNOR2_X1  g222(.A(G116), .B(G119), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT67), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT2), .B(G113), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n408), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n407), .A2(new_n412), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT68), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(KEYINPUT68), .A3(new_n415), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n403), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n413), .A2(KEYINPUT68), .A3(new_n415), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n274), .A2(new_n199), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n253), .B1(G131), .B2(new_n400), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n242), .A2(new_n243), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n392), .B1(new_n420), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n403), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT28), .B1(new_n429), .B2(new_n422), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n391), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT69), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n433), .B(new_n391), .C1(new_n428), .C2(new_n430), .ZN(new_n434));
  INV_X1    g248(.A(new_n427), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n403), .A2(KEYINPUT30), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n423), .A2(new_n426), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n435), .B1(new_n439), .B2(new_n419), .ZN(new_n440));
  INV_X1    g254(.A(new_n391), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT31), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n422), .B1(new_n436), .B2(new_n438), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT31), .ZN(new_n444));
  NOR4_X1   g258(.A1(new_n443), .A2(new_n435), .A3(new_n444), .A4(new_n391), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n432), .B(new_n434), .C1(new_n442), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G472), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n191), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT32), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT32), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n446), .A2(new_n450), .A3(new_n447), .A4(new_n191), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n440), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT29), .B1(new_n453), .B2(new_n391), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n428), .A2(new_n430), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n391), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n391), .ZN(new_n457));
  AOI21_X1  g271(.A(G902), .B1(new_n457), .B2(KEYINPUT29), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G472), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n386), .B1(new_n452), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G214), .B1(G237), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n354), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n198), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n198), .A2(KEYINPUT89), .A3(new_n463), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n253), .A2(new_n354), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT90), .B(G224), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G953), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n470), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT5), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n408), .B2(new_n411), .ZN(new_n475));
  OAI21_X1  g289(.A(G113), .B1(new_n404), .B2(KEYINPUT5), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n415), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n262), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n213), .B1(new_n223), .B2(new_n227), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n422), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G122), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n479), .B(new_n484), .C1(new_n480), .C2(new_n422), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(KEYINPUT6), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n481), .A2(new_n489), .A3(new_n485), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n473), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G210), .B1(G237), .B2(G902), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n492), .B(KEYINPUT94), .Z(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT92), .B1(new_n253), .B2(new_n354), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n496), .B(new_n463), .C1(new_n251), .C2(new_n252), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n464), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT7), .B1(new_n471), .B2(G953), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n498), .B2(new_n500), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n484), .B(KEYINPUT8), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n262), .B2(new_n477), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n407), .A2(new_n474), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n415), .B1(new_n507), .B2(new_n476), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n262), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n504), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n478), .A2(new_n280), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n512), .A2(KEYINPUT91), .A3(new_n509), .A4(new_n505), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n500), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n468), .A2(new_n469), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n503), .A2(new_n514), .A3(new_n487), .A4(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n491), .A2(new_n191), .A3(new_n494), .A4(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n516), .B1(new_n501), .B2(new_n502), .ZN(new_n520));
  INV_X1    g334(.A(new_n487), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(G902), .B1(new_n522), .B2(new_n514), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n494), .B1(new_n523), .B2(new_n491), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n462), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n289), .A2(G952), .ZN(new_n526));
  INV_X1    g340(.A(G237), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n526), .B1(new_n375), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n191), .B(new_n289), .C1(G234), .C2(G237), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT21), .B(G898), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(G143), .B1(new_n387), .B2(G214), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n387), .A2(G143), .A3(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT17), .A3(G131), .ZN(new_n537));
  INV_X1    g351(.A(new_n535), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n533), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n236), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(G131), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n357), .A2(new_n344), .A3(new_n537), .A4(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(G113), .B(G122), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n204), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n539), .B1(new_n547), .B2(new_n236), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n350), .A2(G146), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n355), .A2(new_n245), .ZN(new_n550));
  OAI221_X1 g364(.A(new_n548), .B1(new_n541), .B2(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n544), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n546), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT19), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n245), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n344), .A2(new_n556), .A3(KEYINPUT95), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n540), .A2(new_n541), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT95), .B1(new_n344), .B2(new_n556), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n551), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n552), .B1(new_n553), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G475), .A2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT20), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n553), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n544), .A2(new_n546), .A3(new_n551), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT20), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n563), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n546), .B1(new_n544), .B2(new_n551), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n191), .B1(new_n552), .B2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT96), .B(G475), .Z(new_n573));
  AOI22_X1  g387(.A1(new_n565), .A2(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G217), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n187), .A2(new_n575), .A3(G953), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n195), .A2(G143), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n195), .A3(G143), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT97), .B1(new_n247), .B2(G128), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n578), .B(new_n579), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n581), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n247), .A2(G128), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT99), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n231), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(G116), .B(G122), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G107), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT13), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n582), .A2(new_n581), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n593), .A2(KEYINPUT98), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n593), .A2(KEYINPUT98), .B1(KEYINPUT13), .B2(new_n579), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n231), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n577), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n580), .B1(new_n195), .B2(G143), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n247), .A2(KEYINPUT97), .A3(G128), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n585), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n578), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n584), .A2(KEYINPUT99), .A3(new_n585), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n589), .B1(new_n603), .B2(new_n231), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n593), .A2(KEYINPUT98), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n579), .A2(KEYINPUT13), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n593), .A2(KEYINPUT98), .ZN(new_n608));
  OAI21_X1  g422(.A(G134), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n604), .A2(new_n609), .A3(KEYINPUT100), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n597), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G122), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G116), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n202), .B1(new_n613), .B2(KEYINPUT14), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n588), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n601), .A2(G134), .A3(new_n602), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n587), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n576), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n576), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n618), .B(new_n621), .C1(new_n597), .C2(new_n610), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n191), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G478), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(KEYINPUT15), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n623), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n574), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n525), .A2(new_n532), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n310), .A2(new_n461), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G101), .ZN(G3));
  NAND2_X1  g445(.A1(new_n448), .A2(KEYINPUT101), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n447), .B1(new_n446), .B2(new_n191), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n386), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n310), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n518), .A2(KEYINPUT102), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n517), .A2(new_n191), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n473), .A2(new_n488), .A3(new_n490), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n493), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n523), .A2(new_n642), .A3(new_n494), .A4(new_n491), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n638), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n462), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n624), .B(new_n191), .C1(new_n620), .C2(new_n622), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n620), .A2(new_n622), .A3(KEYINPUT33), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n591), .A2(new_n596), .A3(new_n577), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT100), .B1(new_n604), .B2(new_n609), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n619), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n621), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n611), .A2(new_n619), .A3(new_n576), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n191), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n647), .B1(new_n656), .B2(G478), .ZN(new_n657));
  INV_X1    g471(.A(new_n532), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n572), .A2(new_n573), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n569), .B1(new_n568), .B2(new_n563), .ZN(new_n660));
  AOI211_X1 g474(.A(KEYINPUT20), .B(new_n564), .C1(new_n566), .C2(new_n567), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n645), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n637), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT103), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT34), .B(G104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NOR2_X1   g482(.A1(new_n662), .A2(new_n627), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n658), .A2(new_n644), .A3(new_n462), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n637), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  OR2_X1    g487(.A1(new_n370), .A2(KEYINPUT36), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n365), .A2(new_n371), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n674), .B1(new_n365), .B2(new_n371), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n378), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n381), .B2(new_n385), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n634), .A2(new_n310), .A3(new_n629), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT37), .B(G110), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT104), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(G12));
  INV_X1    g497(.A(new_n385), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n380), .A2(KEYINPUT25), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n452), .A2(new_n460), .B1(new_n686), .B2(new_n678), .ZN(new_n687));
  INV_X1    g501(.A(new_n645), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n623), .B(new_n625), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n574), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n529), .B1(new_n530), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n687), .A2(new_n310), .A3(new_n688), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  XOR2_X1   g509(.A(new_n692), .B(KEYINPUT39), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n310), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT40), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n440), .A2(new_n441), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n420), .A2(new_n427), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n700), .B1(new_n441), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n447), .B1(new_n702), .B2(new_n191), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n449), .B2(new_n451), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n641), .A2(new_n518), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n662), .A2(new_n689), .A3(new_n462), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n679), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n699), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND2_X1  g526(.A1(new_n656), .A2(G478), .ZN(new_n713));
  INV_X1    g527(.A(new_n692), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n662), .A3(new_n646), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT106), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n657), .A2(new_n717), .A3(new_n662), .A4(new_n714), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n687), .A2(new_n310), .A3(new_n719), .A4(new_n688), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  INV_X1    g535(.A(new_n461), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n296), .A2(new_n300), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n190), .A3(new_n191), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n299), .B1(new_n293), .B2(new_n295), .ZN(new_n725));
  OAI21_X1  g539(.A(G469), .B1(new_n725), .B2(G902), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n188), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n664), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT107), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND2_X1  g546(.A1(new_n728), .A2(new_n670), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  NOR2_X1   g548(.A1(new_n727), .A2(new_n645), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n628), .A2(new_n532), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n687), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  AND4_X1   g552(.A1(new_n188), .A2(new_n724), .A3(new_n658), .A4(new_n726), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n662), .A2(new_n689), .A3(KEYINPUT108), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT108), .B1(new_n662), .B2(new_n689), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n645), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n447), .A2(new_n191), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n700), .A2(new_n444), .ZN(new_n745));
  INV_X1    g559(.A(new_n445), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n744), .B1(new_n747), .B2(new_n431), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n386), .A2(new_n633), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n739), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NOR2_X1   g565(.A1(new_n633), .A2(new_n748), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n679), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n735), .A2(new_n719), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NAND4_X1  g569(.A1(new_n641), .A2(new_n188), .A3(new_n462), .A4(new_n518), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n305), .A2(new_n190), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n756), .B1(new_n302), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n719), .A2(new_n758), .A3(new_n461), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT42), .Z(new_n760));
  XOR2_X1   g574(.A(KEYINPUT109), .B(G131), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G33));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n693), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n693), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n758), .B(new_n461), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  INV_X1    g582(.A(new_n679), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n634), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n657), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n662), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT43), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT44), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(KEYINPUT44), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n641), .A2(new_n462), .A3(new_n518), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n306), .B2(new_n308), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  OAI21_X1  g594(.A(G469), .B1(new_n305), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n192), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT46), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n724), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(KEYINPUT46), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n188), .B(new_n696), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n778), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  INV_X1    g605(.A(new_n719), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n449), .A2(new_n451), .B1(G472), .B2(new_n459), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n792), .A2(new_n794), .A3(new_n635), .A4(new_n777), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n188), .B1(new_n786), .B2(new_n787), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT47), .B(new_n188), .C1(new_n786), .C2(new_n787), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n795), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  NAND2_X1  g617(.A1(new_n724), .A2(new_n726), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT49), .Z(new_n805));
  INV_X1    g619(.A(new_n462), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n189), .A2(new_n806), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n635), .A2(new_n708), .A3(new_n772), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n805), .A2(new_n808), .A3(new_n704), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n758), .A2(new_n719), .A3(new_n811), .A4(new_n753), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n724), .A2(new_n783), .A3(new_n757), .ZN(new_n813));
  INV_X1    g627(.A(new_n756), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n716), .A2(new_n679), .A3(new_n718), .A4(new_n752), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT114), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n777), .A2(new_n628), .A3(new_n692), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n687), .A2(new_n310), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n767), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n810), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n812), .A2(new_n817), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n823), .A2(KEYINPUT115), .A3(new_n767), .A4(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n663), .A2(new_n525), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n690), .A2(KEYINPUT112), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT112), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n574), .A2(new_n689), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n706), .A2(new_n658), .A3(new_n462), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT113), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n525), .A2(new_n532), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n827), .A4(new_n829), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n826), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n630), .B(new_n680), .C1(new_n836), .C2(new_n636), .ZN(new_n837));
  INV_X1    g651(.A(new_n727), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(new_n461), .C1(new_n664), .C2(new_n670), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n737), .A3(new_n750), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT111), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n839), .A2(new_n737), .A3(new_n750), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n837), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n692), .B(KEYINPUT116), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n188), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n679), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n743), .A2(new_n705), .A3(new_n813), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n720), .A2(new_n694), .A3(new_n754), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n724), .A2(new_n309), .A3(new_n783), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n688), .A2(new_n852), .A3(new_n188), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n793), .A2(new_n769), .A3(new_n765), .ZN(new_n854));
  INV_X1    g668(.A(new_n816), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n853), .A2(new_n854), .B1(new_n855), .B2(new_n735), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n720), .A4(new_n848), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n825), .A2(new_n760), .A3(new_n844), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n837), .A2(new_n860), .A3(new_n840), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n825), .A2(new_n760), .A3(new_n858), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n773), .A2(new_n529), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n749), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n838), .A2(new_n806), .A3(new_n708), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT50), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n804), .A2(new_n756), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n869), .A2(new_n753), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n386), .A2(new_n528), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n704), .A3(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n878), .A2(new_n662), .A3(new_n657), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n874), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n798), .B(new_n800), .C1(new_n188), .C2(new_n804), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n706), .A2(new_n806), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n871), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n883), .A3(KEYINPUT51), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n869), .A2(new_n461), .A3(new_n875), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT48), .Z(new_n886));
  NOR3_X1   g700(.A1(new_n878), .A2(new_n574), .A3(new_n771), .ZN(new_n887));
  INV_X1    g701(.A(new_n735), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n526), .B1(new_n870), .B2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT51), .B1(new_n880), .B2(new_n883), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n868), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(G952), .A2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n809), .B1(new_n893), .B2(new_n894), .ZN(G75));
  XNOR2_X1  g709(.A(new_n473), .B(KEYINPUT55), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n488), .A2(new_n490), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT117), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n191), .B1(new_n863), .B2(new_n866), .ZN(new_n901));
  AOI211_X1 g715(.A(KEYINPUT56), .B(new_n900), .C1(new_n901), .C2(new_n493), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n863), .A2(new_n866), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(G902), .A3(new_n493), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n897), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n191), .B(new_n494), .C1(new_n863), .C2(new_n866), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n900), .B1(new_n908), .B2(KEYINPUT56), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n904), .A2(new_n905), .A3(new_n899), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n896), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n289), .A2(G952), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT118), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n907), .A2(new_n911), .A3(new_n913), .ZN(G51));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n867), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n863), .A2(KEYINPUT120), .A3(new_n864), .A4(new_n866), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n783), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n723), .ZN(new_n923));
  INV_X1    g737(.A(new_n901), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n924), .A2(new_n782), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n912), .B1(new_n923), .B2(new_n925), .ZN(G54));
  INV_X1    g740(.A(new_n912), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n568), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n568), .B2(new_n928), .ZN(G60));
  XNOR2_X1  g744(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n624), .A2(new_n191), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n931), .B(new_n932), .Z(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n862), .B2(new_n867), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n648), .A2(new_n655), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n913), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n933), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n919), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n936), .A2(new_n938), .ZN(G63));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT60), .B1(new_n575), .B2(new_n191), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n575), .A2(new_n191), .A3(KEYINPUT60), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n903), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n677), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n913), .B1(new_n943), .B2(new_n374), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n943), .A2(new_n374), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n913), .A4(new_n944), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(G953), .B1(new_n531), .B2(new_n471), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n844), .B2(G953), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n900), .B1(G898), .B2(new_n289), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  AOI21_X1  g769(.A(new_n289), .B1(G227), .B2(G900), .ZN(new_n956));
  INV_X1    g770(.A(new_n796), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n743), .A2(new_n461), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n957), .A2(new_n958), .A3(new_n696), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT126), .B1(new_n788), .B2(new_n959), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n760), .A2(new_n767), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n856), .A2(new_n720), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n778), .B2(new_n789), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n802), .A2(new_n963), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(G953), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n554), .A2(new_n555), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n439), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n970), .ZN(new_n973));
  INV_X1    g787(.A(new_n965), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n711), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n697), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n830), .B1(new_n574), .B2(new_n771), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n980), .A2(new_n461), .A3(new_n882), .A4(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n979), .A2(new_n802), .A3(new_n790), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n973), .B1(new_n983), .B2(new_n289), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n956), .B1(new_n972), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n956), .B(KEYINPUT125), .Z(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n968), .B2(new_n971), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n984), .A2(new_n986), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n985), .A2(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(new_n453), .A2(new_n441), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n440), .A2(new_n391), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT63), .Z(new_n997));
  OAI21_X1  g811(.A(new_n927), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI22_X1  g812(.A1(new_n983), .A2(new_n993), .B1(new_n967), .B2(new_n994), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(new_n844), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n861), .A2(new_n997), .A3(new_n995), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n1002), .A2(new_n1001), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(G57));
endmodule


